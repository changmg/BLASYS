module max_12_0(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , po0 , po1 , po2 , po3 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 ;
  output po0 , po1 , po2 , po3 ;
  wire new_n8, new_n9, new_n10, new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22;
  assign new_n8 = pi0 & ~pi5 ;
  assign new_n9 = ~pi4 & ~new_n8 ;
  assign new_n10 = ~pi0 & pi5 ;
  assign new_n11 = ~pi1 & pi6 ;
  assign new_n12 = ~new_n10 & ~new_n11 ;
  assign new_n13 = ~new_n9 & new_n12 ;
  assign new_n14 = pi1 & ~pi6 ;
  assign new_n15 = ~pi2 & ~new_n14 ;
  assign new_n16 = ~new_n13 & new_n15 ;
  assign new_n17 = pi3 & ~pi5 ;
  assign new_n18 = ~pi0 & ~pi3 ;
  assign new_n19 = ~new_n17 & ~new_n18 ;
  assign new_n20 = pi3 & ~pi6 ;
  assign new_n21 = ~pi1 & ~pi3 ;
  assign new_n22 = ~new_n20 & ~new_n21 ;
  assign po0 = pi3 ;
  assign po1 = new_n16 ;
  assign po2 = new_n19 ;
  assign po3 = new_n22 ;
endmodule
