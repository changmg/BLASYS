// Benchmark "ex" written by ABC on Thu Jul 14 00:31:25 2022

module ex ( 
    a, b, c, d, e, f, g,
    F  );
  input  a, b, c, d, e, f, g;
  output F;
  assign F = e;
endmodule


