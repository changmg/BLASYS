module adder(\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] 
, \a[21] , \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] 
, \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] 
, \a[63] , \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] 
, \a[84] , \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] 
, \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] , \a[125] 
, \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] 
, \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] 
, \b[40] , \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] 
, \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] 
, \b[82] , \b[83] , \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] , \b[100] , \b[101] , \b[102] 
, \b[103] , \b[104] , \b[105] , \b[106] , \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] , \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] , \b[121] , \b[122] , \b[123] 
, \b[124] , \b[125] , \b[126] , \b[127] , \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] 
, \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] 
, \f[38] , \f[39] , \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] , \f[57] , \f[58] 
, \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] 
, \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] , \f[97] , \f[98] , \f[99] , \f[100] 
, \f[101] , \f[102] , \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] , \f[118] , \f[119] , \f[120] , \f[121] 
, \f[122] , \f[123] , \f[124] , \f[125] , \f[126] , \f[127] , cOut);
  input \a[0] ;
  input \a[100] ;
  input \a[101] ;
  input \a[102] ;
  input \a[103] ;
  input \a[104] ;
  input \a[105] ;
  input \a[106] ;
  input \a[107] ;
  input \a[108] ;
  input \a[109] ;
  input \a[10] ;
  input \a[110] ;
  input \a[111] ;
  input \a[112] ;
  input \a[113] ;
  input \a[114] ;
  input \a[115] ;
  input \a[116] ;
  input \a[117] ;
  input \a[118] ;
  input \a[119] ;
  input \a[11] ;
  input \a[120] ;
  input \a[121] ;
  input \a[122] ;
  input \a[123] ;
  input \a[124] ;
  input \a[125] ;
  input \a[126] ;
  input \a[127] ;
  input \a[12] ;
  input \a[13] ;
  input \a[14] ;
  input \a[15] ;
  input \a[16] ;
  input \a[17] ;
  input \a[18] ;
  input \a[19] ;
  input \a[1] ;
  input \a[20] ;
  input \a[21] ;
  input \a[22] ;
  input \a[23] ;
  input \a[24] ;
  input \a[25] ;
  input \a[26] ;
  input \a[27] ;
  input \a[28] ;
  input \a[29] ;
  input \a[2] ;
  input \a[30] ;
  input \a[31] ;
  input \a[32] ;
  input \a[33] ;
  input \a[34] ;
  input \a[35] ;
  input \a[36] ;
  input \a[37] ;
  input \a[38] ;
  input \a[39] ;
  input \a[3] ;
  input \a[40] ;
  input \a[41] ;
  input \a[42] ;
  input \a[43] ;
  input \a[44] ;
  input \a[45] ;
  input \a[46] ;
  input \a[47] ;
  input \a[48] ;
  input \a[49] ;
  input \a[4] ;
  input \a[50] ;
  input \a[51] ;
  input \a[52] ;
  input \a[53] ;
  input \a[54] ;
  input \a[55] ;
  input \a[56] ;
  input \a[57] ;
  input \a[58] ;
  input \a[59] ;
  input \a[5] ;
  input \a[60] ;
  input \a[61] ;
  input \a[62] ;
  input \a[63] ;
  input \a[64] ;
  input \a[65] ;
  input \a[66] ;
  input \a[67] ;
  input \a[68] ;
  input \a[69] ;
  input \a[6] ;
  input \a[70] ;
  input \a[71] ;
  input \a[72] ;
  input \a[73] ;
  input \a[74] ;
  input \a[75] ;
  input \a[76] ;
  input \a[77] ;
  input \a[78] ;
  input \a[79] ;
  input \a[7] ;
  input \a[80] ;
  input \a[81] ;
  input \a[82] ;
  input \a[83] ;
  input \a[84] ;
  input \a[85] ;
  input \a[86] ;
  input \a[87] ;
  input \a[88] ;
  input \a[89] ;
  input \a[8] ;
  input \a[90] ;
  input \a[91] ;
  input \a[92] ;
  input \a[93] ;
  input \a[94] ;
  input \a[95] ;
  input \a[96] ;
  input \a[97] ;
  input \a[98] ;
  input \a[99] ;
  input \a[9] ;
  input \b[0] ;
  input \b[100] ;
  input \b[101] ;
  input \b[102] ;
  input \b[103] ;
  input \b[104] ;
  input \b[105] ;
  input \b[106] ;
  input \b[107] ;
  input \b[108] ;
  input \b[109] ;
  input \b[10] ;
  input \b[110] ;
  input \b[111] ;
  input \b[112] ;
  input \b[113] ;
  input \b[114] ;
  input \b[115] ;
  input \b[116] ;
  input \b[117] ;
  input \b[118] ;
  input \b[119] ;
  input \b[11] ;
  input \b[120] ;
  input \b[121] ;
  input \b[122] ;
  input \b[123] ;
  input \b[124] ;
  input \b[125] ;
  input \b[126] ;
  input \b[127] ;
  input \b[12] ;
  input \b[13] ;
  input \b[14] ;
  input \b[15] ;
  input \b[16] ;
  input \b[17] ;
  input \b[18] ;
  input \b[19] ;
  input \b[1] ;
  input \b[20] ;
  input \b[21] ;
  input \b[22] ;
  input \b[23] ;
  input \b[24] ;
  input \b[25] ;
  input \b[26] ;
  input \b[27] ;
  input \b[28] ;
  input \b[29] ;
  input \b[2] ;
  input \b[30] ;
  input \b[31] ;
  input \b[32] ;
  input \b[33] ;
  input \b[34] ;
  input \b[35] ;
  input \b[36] ;
  input \b[37] ;
  input \b[38] ;
  input \b[39] ;
  input \b[3] ;
  input \b[40] ;
  input \b[41] ;
  input \b[42] ;
  input \b[43] ;
  input \b[44] ;
  input \b[45] ;
  input \b[46] ;
  input \b[47] ;
  input \b[48] ;
  input \b[49] ;
  input \b[4] ;
  input \b[50] ;
  input \b[51] ;
  input \b[52] ;
  input \b[53] ;
  input \b[54] ;
  input \b[55] ;
  input \b[56] ;
  input \b[57] ;
  input \b[58] ;
  input \b[59] ;
  input \b[5] ;
  input \b[60] ;
  input \b[61] ;
  input \b[62] ;
  input \b[63] ;
  input \b[64] ;
  input \b[65] ;
  input \b[66] ;
  input \b[67] ;
  input \b[68] ;
  input \b[69] ;
  input \b[6] ;
  input \b[70] ;
  input \b[71] ;
  input \b[72] ;
  input \b[73] ;
  input \b[74] ;
  input \b[75] ;
  input \b[76] ;
  input \b[77] ;
  input \b[78] ;
  input \b[79] ;
  input \b[7] ;
  input \b[80] ;
  input \b[81] ;
  input \b[82] ;
  input \b[83] ;
  input \b[84] ;
  input \b[85] ;
  input \b[86] ;
  input \b[87] ;
  input \b[88] ;
  input \b[89] ;
  input \b[8] ;
  input \b[90] ;
  input \b[91] ;
  input \b[92] ;
  input \b[93] ;
  input \b[94] ;
  input \b[95] ;
  input \b[96] ;
  input \b[97] ;
  input \b[98] ;
  input \b[99] ;
  input \b[9] ;
  output cOut;
  output \f[0] ;
  output \f[100] ;
  output \f[101] ;
  output \f[102] ;
  output \f[103] ;
  output \f[104] ;
  output \f[105] ;
  output \f[106] ;
  output \f[107] ;
  output \f[108] ;
  output \f[109] ;
  output \f[10] ;
  output \f[110] ;
  output \f[111] ;
  output \f[112] ;
  output \f[113] ;
  output \f[114] ;
  output \f[115] ;
  output \f[116] ;
  output \f[117] ;
  output \f[118] ;
  output \f[119] ;
  output \f[11] ;
  output \f[120] ;
  output \f[121] ;
  output \f[122] ;
  output \f[123] ;
  output \f[124] ;
  output \f[125] ;
  output \f[126] ;
  output \f[127] ;
  output \f[12] ;
  output \f[13] ;
  output \f[14] ;
  output \f[15] ;
  output \f[16] ;
  output \f[17] ;
  output \f[18] ;
  output \f[19] ;
  output \f[1] ;
  output \f[20] ;
  output \f[21] ;
  output \f[22] ;
  output \f[23] ;
  output \f[24] ;
  output \f[25] ;
  output \f[26] ;
  output \f[27] ;
  output \f[28] ;
  output \f[29] ;
  output \f[2] ;
  output \f[30] ;
  output \f[31] ;
  output \f[32] ;
  output \f[33] ;
  output \f[34] ;
  output \f[35] ;
  output \f[36] ;
  output \f[37] ;
  output \f[38] ;
  output \f[39] ;
  output \f[3] ;
  output \f[40] ;
  output \f[41] ;
  output \f[42] ;
  output \f[43] ;
  output \f[44] ;
  output \f[45] ;
  output \f[46] ;
  output \f[47] ;
  output \f[48] ;
  output \f[49] ;
  output \f[4] ;
  output \f[50] ;
  output \f[51] ;
  output \f[52] ;
  output \f[53] ;
  output \f[54] ;
  output \f[55] ;
  output \f[56] ;
  output \f[57] ;
  output \f[58] ;
  output \f[59] ;
  output \f[5] ;
  output \f[60] ;
  output \f[61] ;
  output \f[62] ;
  output \f[63] ;
  output \f[64] ;
  output \f[65] ;
  output \f[66] ;
  output \f[67] ;
  output \f[68] ;
  output \f[69] ;
  output \f[6] ;
  output \f[70] ;
  output \f[71] ;
  output \f[72] ;
  output \f[73] ;
  output \f[74] ;
  output \f[75] ;
  output \f[76] ;
  output \f[77] ;
  output \f[78] ;
  output \f[79] ;
  output \f[7] ;
  output \f[80] ;
  output \f[81] ;
  output \f[82] ;
  output \f[83] ;
  output \f[84] ;
  output \f[85] ;
  output \f[86] ;
  output \f[87] ;
  output \f[88] ;
  output \f[89] ;
  output \f[8] ;
  output \f[90] ;
  output \f[91] ;
  output \f[92] ;
  output \f[93] ;
  output \f[94] ;
  output \f[95] ;
  output \f[96] ;
  output \f[97] ;
  output \f[98] ;
  output \f[99] ;
  output \f[9] ;
  top U0 ( .pi000( \a[0] ) , .pi001( \a[1] ) , .pi002( \a[2] ) , .pi003( \a[3] ) , .pi004( \a[4] ) , .pi005( \a[5] ) , .pi006( \a[6] ) , .pi007( \a[7] ) , .pi008( \a[8] ) , .pi009( \a[9] ) , .pi010( \a[10] ) , .pi011( \a[11] ) , .pi012( \a[12] ) , .pi013( \a[13] ) , .pi014( \a[14] ) , .pi015( \a[15] ) , .pi016( \a[16] ) , .pi017( \a[17] ) , .pi018( \a[18] ) , .pi019( \a[19] ) , .pi020( \a[20] ) , .pi021( \a[21] ) , .pi022( \a[22] ) , .pi023( \a[23] ) , .pi024( \a[24] ) , .pi025( \a[25] ) , .pi026( \a[26] ) , .pi027( \a[27] ) , .pi028( \a[28] ) , .pi029( \a[29] ) , .pi030( \a[30] ) , .pi031( \a[31] ) , .pi032( \a[32] ) , .pi033( \a[33] ) , .pi034( \a[34] ) , .pi035( \a[35] ) , .pi036( \a[36] ) , .pi037( \a[37] ) , .pi038( \a[38] ) , .pi039( \a[39] ) , .pi040( \a[40] ) , .pi041( \a[41] ) , .pi042( \a[42] ) , .pi043( \a[43] ) , .pi044( \a[44] ) , .pi045( \a[45] ) , .pi046( \a[46] ) , .pi047( \a[47] ) , .pi048( \a[48] ) , .pi049( \a[49] ) , .pi050( \a[50] ) , .pi051( \a[51] ) , .pi052( \a[52] ) , .pi053( \a[53] ) , .pi054( \a[54] ) , .pi055( \a[55] ) , .pi056( \a[56] ) , .pi057( \a[57] ) , .pi058( \a[58] ) , .pi059( \a[59] ) , .pi060( \a[60] ) , .pi061( \a[61] ) , .pi062( \a[62] ) , .pi063( \a[63] ) , .pi064( \a[64] ) , .pi065( \a[65] ) , .pi066( \a[66] ) , .pi067( \a[67] ) , .pi068( \a[68] ) , .pi069( \a[69] ) , .pi070( \a[70] ) , .pi071( \a[71] ) , .pi072( \a[72] ) , .pi073( \a[73] ) , .pi074( \a[74] ) , .pi075( \a[75] ) , .pi076( \a[76] ) , .pi077( \a[77] ) , .pi078( \a[78] ) , .pi079( \a[79] ) , .pi080( \a[80] ) , .pi081( \a[81] ) , .pi082( \a[82] ) , .pi083( \a[83] ) , .pi084( \a[84] ) , .pi085( \a[85] ) , .pi086( \a[86] ) , .pi087( \a[87] ) , .pi088( \a[88] ) , .pi089( \a[89] ) , .pi090( \a[90] ) , .pi091( \a[91] ) , .pi092( \a[92] ) , .pi093( \a[93] ) , .pi094( \a[94] ) , .pi095( \a[95] ) , .pi096( \a[96] ) , .pi097( \a[97] ) , .pi098( \a[98] ) , .pi099( \a[99] ) , .pi100( \a[100] ) , .pi101( \a[101] ) , .pi102( \a[102] ) , .pi103( \a[103] ) , .pi104( \a[104] ) , .pi105( \a[105] ) , .pi106( \a[106] ) , .pi107( \a[107] ) , .pi108( \a[108] ) , .pi109( \a[109] ) , .pi110( \a[110] ) , .pi111( \a[111] ) , .pi112( \a[112] ) , .pi113( \a[113] ) , .pi114( \a[114] ) , .pi115( \a[115] ) , .pi116( \a[116] ) , .pi117( \a[117] ) , .pi118( \a[118] ) , .pi119( \a[119] ) , .pi120( \a[120] ) , .pi121( \a[121] ) , .pi122( \a[122] ) , .pi123( \a[123] ) , .pi124( \a[124] ) , .pi125( \a[125] ) , .pi126( \a[126] ) , .pi127( \a[127] ) , .pi128( \b[0] ) , .pi129( \b[1] ) , .pi130( \b[2] ) , .pi131( \b[3] ) , .pi132( \b[4] ) , .pi133( \b[5] ) , .pi134( \b[6] ) , .pi135( \b[7] ) , .pi136( \b[8] ) , .pi137( \b[9] ) , .pi138( \b[10] ) , .pi139( \b[11] ) , .pi140( \b[12] ) , .pi141( \b[13] ) , .pi142( \b[14] ) , .pi143( \b[15] ) , .pi144( \b[16] ) , .pi145( \b[17] ) , .pi146( \b[18] ) , .pi147( \b[19] ) , .pi148( \b[20] ) , .pi149( \b[21] ) , .pi150( \b[22] ) , .pi151( \b[23] ) , .pi152( \b[24] ) , .pi153( \b[25] ) , .pi154( \b[26] ) , .pi155( \b[27] ) , .pi156( \b[28] ) , .pi157( \b[29] ) , .pi158( \b[30] ) , .pi159( \b[31] ) , .pi160( \b[32] ) , .pi161( \b[33] ) , .pi162( \b[34] ) , .pi163( \b[35] ) , .pi164( \b[36] ) , .pi165( \b[37] ) , .pi166( \b[38] ) , .pi167( \b[39] ) , .pi168( \b[40] ) , .pi169( \b[41] ) , .pi170( \b[42] ) , .pi171( \b[43] ) , .pi172( \b[44] ) , .pi173( \b[45] ) , .pi174( \b[46] ) , .pi175( \b[47] ) , .pi176( \b[48] ) , .pi177( \b[49] ) , .pi178( \b[50] ) , .pi179( \b[51] ) , .pi180( \b[52] ) , .pi181( \b[53] ) , .pi182( \b[54] ) , .pi183( \b[55] ) , .pi184( \b[56] ) , .pi185( \b[57] ) , .pi186( \b[58] ) , .pi187( \b[59] ) , .pi188( \b[60] ) , .pi189( \b[61] ) , .pi190( \b[62] ) , .pi191( \b[63] ) , .pi192( \b[64] ) , .pi193( \b[65] ) , .pi194( \b[66] ) , .pi195( \b[67] ) , .pi196( \b[68] ) , .pi197( \b[69] ) , .pi198( \b[70] ) , .pi199( \b[71] ) , .pi200( \b[72] ) , .pi201( \b[73] ) , .pi202( \b[74] ) , .pi203( \b[75] ) , .pi204( \b[76] ) , .pi205( \b[77] ) , .pi206( \b[78] ) , .pi207( \b[79] ) , .pi208( \b[80] ) , .pi209( \b[81] ) , .pi210( \b[82] ) , .pi211( \b[83] ) , .pi212( \b[84] ) , .pi213( \b[85] ) , .pi214( \b[86] ) , .pi215( \b[87] ) , .pi216( \b[88] ) , .pi217( \b[89] ) , .pi218( \b[90] ) , .pi219( \b[91] ) , .pi220( \b[92] ) , .pi221( \b[93] ) , .pi222( \b[94] ) , .pi223( \b[95] ) , .pi224( \b[96] ) , .pi225( \b[97] ) , .pi226( \b[98] ) , .pi227( \b[99] ) , .pi228( \b[100] ) , .pi229( \b[101] ) , .pi230( \b[102] ) , .pi231( \b[103] ) , .pi232( \b[104] ) , .pi233( \b[105] ) , .pi234( \b[106] ) , .pi235( \b[107] ) , .pi236( \b[108] ) , .pi237( \b[109] ) , .pi238( \b[110] ) , .pi239( \b[111] ) , .pi240( \b[112] ) , .pi241( \b[113] ) , .pi242( \b[114] ) , .pi243( \b[115] ) , .pi244( \b[116] ) , .pi245( \b[117] ) , .pi246( \b[118] ) , .pi247( \b[119] ) , .pi248( \b[120] ) , .pi249( \b[121] ) , .pi250( \b[122] ) , .pi251( \b[123] ) , .pi252( \b[124] ) , .pi253( \b[125] ) , .pi254( \b[126] ) , .pi255( \b[127] ) , .po000( \f[0] ) , .po001( \f[1] ) , .po002( \f[2] ) , .po003( \f[3] ) , .po004( \f[4] ) , .po005( \f[5] ) , .po006( \f[6] ) , .po007( \f[7] ) , .po008( \f[8] ) , .po009( \f[9] ) , .po010( \f[10] ) , .po011( \f[11] ) , .po012( \f[12] ) , .po013( \f[13] ) , .po014( \f[14] ) , .po015( \f[15] ) , .po016( \f[16] ) , .po017( \f[17] ) , .po018( \f[18] ) , .po019( \f[19] ) , .po020( \f[20] ) , .po021( \f[21] ) , .po022( \f[22] ) , .po023( \f[23] ) , .po024( \f[24] ) , .po025( \f[25] ) , .po026( \f[26] ) , .po027( \f[27] ) , .po028( \f[28] ) , .po029( \f[29] ) , .po030( \f[30] ) , .po031( \f[31] ) , .po032( \f[32] ) , .po033( \f[33] ) , .po034( \f[34] ) , .po035( \f[35] ) , .po036( \f[36] ) , .po037( \f[37] ) , .po038( \f[38] ) , .po039( \f[39] ) , .po040( \f[40] ) , .po041( \f[41] ) , .po042( \f[42] ) , .po043( \f[43] ) , .po044( \f[44] ) , .po045( \f[45] ) , .po046( \f[46] ) , .po047( \f[47] ) , .po048( \f[48] ) , .po049( \f[49] ) , .po050( \f[50] ) , .po051( \f[51] ) , .po052( \f[52] ) , .po053( \f[53] ) , .po054( \f[54] ) , .po055( \f[55] ) , .po056( \f[56] ) , .po057( \f[57] ) , .po058( \f[58] ) , .po059( \f[59] ) , .po060( \f[60] ) , .po061( \f[61] ) , .po062( \f[62] ) , .po063( \f[63] ) , .po064( \f[64] ) , .po065( \f[65] ) , .po066( \f[66] ) , .po067( \f[67] ) , .po068( \f[68] ) , .po069( \f[69] ) , .po070( \f[70] ) , .po071( \f[71] ) , .po072( \f[72] ) , .po073( \f[73] ) , .po074( \f[74] ) , .po075( \f[75] ) , .po076( \f[76] ) , .po077( \f[77] ) , .po078( \f[78] ) , .po079( \f[79] ) , .po080( \f[80] ) , .po081( \f[81] ) , .po082( \f[82] ) , .po083( \f[83] ) , .po084( \f[84] ) , .po085( \f[85] ) , .po086( \f[86] ) , .po087( \f[87] ) , .po088( \f[88] ) , .po089( \f[89] ) , .po090( \f[90] ) , .po091( \f[91] ) , .po092( \f[92] ) , .po093( \f[93] ) , .po094( \f[94] ) , .po095( \f[95] ) , .po096( \f[96] ) , .po097( \f[97] ) , .po098( \f[98] ) , .po099( \f[99] ) , .po100( \f[100] ) , .po101( \f[101] ) , .po102( \f[102] ) , .po103( \f[103] ) , .po104( \f[104] ) , .po105( \f[105] ) , .po106( \f[106] ) , .po107( \f[107] ) , .po108( \f[108] ) , .po109( \f[109] ) , .po110( \f[110] ) , .po111( \f[111] ) , .po112( \f[112] ) , .po113( \f[113] ) , .po114( \f[114] ) , .po115( \f[115] ) , .po116( \f[116] ) , .po117( \f[117] ) , .po118( \f[118] ) , .po119( \f[119] ) , .po120( \f[120] ) , .po121( \f[121] ) , .po122( \f[122] ) , .po123( \f[123] ) , .po124( \f[124] ) , .po125( \f[125] ) , .po126( \f[126] ) , .po127( \f[127] ) , .po128( cOut ) );
endmodule

module top(pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128);
  input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128;
  wire n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, tpo000, tpo001, tpo002, tpo003, tpo004, tpo005, tpo006, tpo007, tpo008, tpo009, tpo010, tpo011, tpo012, tpo013, tpo014, tpo015, tpo016, tpo017, tpo018, tpo019, tpo020, tpo021, tpo022, tpo023, tpo024, tpo025, tpo026, tpo027, tpo028, tpo029, tpo030, tpo031, tpo032, tpo033, tpo034, tpo035, tpo036, tpo037, tpo038, tpo039, tpo040, tpo041, tpo042, tpo043, tpo044, tpo045, tpo046, tpo047, tpo048, tpo049, tpo050, tpo051, tpo052, tpo053, tpo054, tpo055, tpo056, tpo057, tpo058, tpo059, tpo060, tpo061, tpo062, tpo063, tpo064, tpo065, tpo066, tpo067, tpo068, tpo069, tpo070, tpo071, tpo072, tpo073, tpo074, tpo075, tpo076, tpo077, tpo078, tpo079, tpo080, tpo081, tpo082, tpo083, tpo084, tpo085, tpo086, tpo087, tpo088, tpo089, tpo090, tpo091, tpo092, tpo093, tpo094, tpo095, tpo096, tpo097, tpo098, tpo099, tpo100, tpo101, tpo102, tpo103, tpo104, tpo105, tpo106, tpo107, tpo108, tpo109, tpo110, tpo111, tpo112, tpo113, tpo114, tpo115, tpo116, tpo117, tpo118, tpo119, tpo120, tpo121, tpo122, tpo123, tpo124, tpo125, tpo126, tpo127, tpo128;
  assign po000 = tpo000;
  assign po001 = ~tpo001;
  assign po002 = ~tpo002;
  assign po003 = ~tpo003;
  assign po004 = ~tpo004;
  assign po005 = ~tpo005;
  assign po006 = ~tpo006;
  assign po007 = ~tpo007;
  assign po008 = ~tpo008;
  assign po009 = ~tpo009;
  assign po010 = ~tpo010;
  assign po011 = ~tpo011;
  assign po012 = ~tpo012;
  assign po013 = ~tpo013;
  assign po014 = ~tpo014;
  assign po015 = ~tpo015;
  assign po016 = ~tpo016;
  assign po017 = ~tpo017;
  assign po018 = ~tpo018;
  assign po019 = ~tpo019;
  assign po020 = ~tpo020;
  assign po021 = ~tpo021;
  assign po022 = ~tpo022;
  assign po023 = ~tpo023;
  assign po024 = ~tpo024;
  assign po025 = ~tpo025;
  assign po026 = ~tpo026;
  assign po027 = ~tpo027;
  assign po028 = ~tpo028;
  assign po029 = ~tpo029;
  assign po030 = ~tpo030;
  assign po031 = ~tpo031;
  assign po032 = ~tpo032;
  assign po033 = ~tpo033;
  assign po034 = ~tpo034;
  assign po035 = ~tpo035;
  assign po036 = ~tpo036;
  assign po037 = ~tpo037;
  assign po038 = ~tpo038;
  assign po039 = ~tpo039;
  assign po040 = ~tpo040;
  assign po041 = ~tpo041;
  assign po042 = ~tpo042;
  assign po043 = ~tpo043;
  assign po044 = ~tpo044;
  assign po045 = ~tpo045;
  assign po046 = ~tpo046;
  assign po047 = ~tpo047;
  assign po048 = ~tpo048;
  assign po049 = ~tpo049;
  assign po050 = ~tpo050;
  assign po051 = ~tpo051;
  assign po052 = ~tpo052;
  assign po053 = ~tpo053;
  assign po054 = ~tpo054;
  assign po055 = ~tpo055;
  assign po056 = ~tpo056;
  assign po057 = ~tpo057;
  assign po058 = ~tpo058;
  assign po059 = ~tpo059;
  assign po060 = ~tpo060;
  assign po061 = ~tpo061;
  assign po062 = ~tpo062;
  assign po063 = ~tpo063;
  assign po064 = ~tpo064;
  assign po065 = ~tpo065;
  assign po066 = ~tpo066;
  assign po067 = ~tpo067;
  assign po068 = ~tpo068;
  assign po069 = ~tpo069;
  assign po070 = ~tpo070;
  assign po071 = ~tpo071;
  assign po072 = ~tpo072;
  assign po073 = ~tpo073;
  assign po074 = ~tpo074;
  assign po075 = ~tpo075;
  assign po076 = ~tpo076;
  assign po077 = ~tpo077;
  assign po078 = ~tpo078;
  assign po079 = ~tpo079;
  assign po080 = ~tpo080;
  assign po081 = ~tpo081;
  assign po082 = ~tpo082;
  assign po083 = ~tpo083;
  assign po084 = ~tpo084;
  assign po085 = ~tpo085;
  assign po086 = ~tpo086;
  assign po087 = ~tpo087;
  assign po088 = ~tpo088;
  assign po089 = ~tpo089;
  assign po090 = ~tpo090;
  assign po091 = ~tpo091;
  assign po092 = ~tpo092;
  assign po093 = ~tpo093;
  assign po094 = ~tpo094;
  assign po095 = ~tpo095;
  assign po096 = ~tpo096;
  assign po097 = ~tpo097;
  assign po098 = ~tpo098;
  assign po099 = ~tpo099;
  assign po100 = ~tpo100;
  assign po101 = ~tpo101;
  assign po102 = ~tpo102;
  assign po103 = ~tpo103;
  assign po104 = ~tpo104;
  assign po105 = ~tpo105;
  assign po106 = ~tpo106;
  assign po107 = ~tpo107;
  assign po108 = ~tpo108;
  assign po109 = ~tpo109;
  assign po110 = ~tpo110;
  assign po111 = ~tpo111;
  assign po112 = ~tpo112;
  assign po113 = ~tpo113;
  assign po114 = ~tpo114;
  assign po115 = ~tpo115;
  assign po116 = ~tpo116;
  assign po117 = ~tpo117;
  assign po118 = ~tpo118;
  assign po119 = ~tpo119;
  assign po120 = ~tpo120;
  assign po121 = ~tpo121;
  assign po122 = ~tpo122;
  assign po123 = ~tpo123;
  assign po124 = ~tpo124;
  assign po125 = ~tpo125;
  assign po126 = ~tpo126;
  assign po127 = ~tpo127;
  assign po128 = ~tpo128;
  adder_0 U0 ( .pi00( pi089 ), .pi01( pi090 ), .pi02( pi091 ), .pi03( pi092 ), .pi04( pi093 ), .pi05( pi218 ), .pi06( pi219 ), .pi07( pi220 ), .pi08( pi221 ), .pi09( n36 ), .pi10( n37 ), .po0( tpo089 ), .po1( tpo090 ), .po2( tpo091 ), .po3( tpo092 ), .po4( tpo093 ), .po5( n38 ), .po6( n39 ) );
  adder_1 U1 ( .pi00( pi080 ), .pi01( pi081 ), .pi02( pi082 ), .pi03( pi083 ), .pi04( pi084 ), .pi05( pi208 ), .pi06( pi209 ), .pi07( pi210 ), .pi08( pi211 ), .pi09( pi212 ), .pi10( n32 ), .pi11( n33 ), .po0( tpo080 ), .po1( tpo081 ), .po2( tpo082 ), .po3( tpo083 ), .po4( tpo084 ), .po5( n34 ), .po6( n35 ) );
  adder_2 U2 ( .pi00( pi085 ), .pi01( pi086 ), .pi02( pi087 ), .pi03( pi088 ), .pi04( pi213 ), .pi05( pi214 ), .pi06( pi215 ), .pi07( pi216 ), .pi08( pi217 ), .pi09( n34 ), .pi10( n35 ), .po0( tpo085 ), .po1( tpo086 ), .po2( tpo087 ), .po3( tpo088 ), .po4( n36 ), .po5( n37 ) );
  adder_3 U3 ( .pi00( pi075 ), .pi01( pi076 ), .pi02( pi077 ), .pi03( pi078 ), .pi04( pi079 ), .pi05( pi203 ), .pi06( pi204 ), .pi07( pi205 ), .pi08( pi206 ), .pi09( pi207 ), .pi10( n30 ), .pi11( n31 ), .po0( tpo075 ), .po1( tpo076 ), .po2( tpo077 ), .po3( tpo078 ), .po4( tpo079 ), .po5( n32 ), .po6( n33 ) );
  adder_4 U4 ( .pi00( pi070 ), .pi01( pi071 ), .pi02( pi072 ), .pi03( pi073 ), .pi04( pi074 ), .pi05( pi198 ), .pi06( pi199 ), .pi07( pi200 ), .pi08( pi201 ), .pi09( pi202 ), .pi10( n28 ), .pi11( n29 ), .po0( tpo070 ), .po1( tpo071 ), .po2( tpo072 ), .po3( tpo073 ), .po4( tpo074 ), .po5( n30 ), .po6( n31 ) );
  adder_5 U5 ( .pi00( pi065 ), .pi01( pi066 ), .pi02( pi067 ), .pi03( pi068 ), .pi04( pi069 ), .pi05( pi194 ), .pi06( pi195 ), .pi07( pi196 ), .pi08( pi197 ), .pi09( n26 ), .pi10( n27 ), .po0( tpo065 ), .po1( tpo066 ), .po2( tpo067 ), .po3( tpo068 ), .po4( tpo069 ), .po5( n28 ), .po6( n29 ) );
  adder_6 U6 ( .pi00( pi061 ), .pi01( pi062 ), .pi02( pi063 ), .pi03( pi064 ), .pi04( pi189 ), .pi05( pi190 ), .pi06( pi191 ), .pi07( pi192 ), .pi08( pi193 ), .pi09( n25 ), .po0( tpo061 ), .po1( tpo062 ), .po2( tpo063 ), .po3( tpo064 ), .po4( n26 ), .po5( n27 ) );
  adder_7 U7 ( .pi00( pi094 ), .pi01( pi095 ), .pi02( pi096 ), .pi03( pi097 ), .pi04( pi098 ), .pi05( pi222 ), .pi06( pi223 ), .pi07( pi224 ), .pi08( pi225 ), .pi09( pi226 ), .pi10( pi227 ), .pi11( n38 ), .pi12( n39 ), .po0( tpo094 ), .po1( tpo095 ), .po2( tpo096 ), .po3( tpo097 ), .po4( tpo098 ), .po5( n40 ), .po6( n41 ) );
  adder_8 U8 ( .pi00( pi105 ), .pi01( pi106 ), .pi02( pi107 ), .pi03( pi108 ), .pi04( pi109 ), .pi05( pi233 ), .pi06( pi234 ), .pi07( pi235 ), .pi08( pi236 ), .pi09( pi237 ), .pi10( n42 ), .pi11( n43 ), .po0( tpo105 ), .po1( tpo106 ), .po2( tpo107 ), .po3( tpo108 ), .po4( tpo109 ), .po5( n44 ) );
  adder_9 U9 ( .pi00( pi099 ), .pi01( pi100 ), .pi02( pi101 ), .pi03( pi102 ), .pi04( pi103 ), .pi05( pi104 ), .pi06( pi228 ), .pi07( pi229 ), .pi08( pi230 ), .pi09( pi231 ), .pi10( pi232 ), .pi11( n40 ), .pi12( n41 ), .po0( tpo099 ), .po1( tpo100 ), .po2( tpo101 ), .po3( tpo102 ), .po4( tpo103 ), .po5( tpo104 ), .po6( n42 ), .po7( n43 ) );
  adder_10 U10 ( .pi0( pi126 ), .pi1( pi127 ), .pi2( pi254 ), .pi3( pi255 ), .pi4( n49 ), .po0( tpo126 ), .po1( tpo127 ), .po2( tpo128 ) );
  adder_11 U11 ( .pi00( pi119 ), .pi01( pi120 ), .pi02( pi121 ), .pi03( pi122 ), .pi04( pi123 ), .pi05( pi124 ), .pi06( pi125 ), .pi07( pi247 ), .pi08( pi248 ), .pi09( pi249 ), .pi10( pi250 ), .pi11( pi251 ), .pi12( pi252 ), .pi13( pi253 ), .pi14( n47 ), .pi15( n48 ), .po0( tpo119 ), .po1( tpo120 ), .po2( tpo121 ), .po3( tpo122 ), .po4( tpo123 ), .po5( tpo124 ), .po6( tpo125 ), .po7( n49 ) );
  adder_12 U12 ( .pi00( pi110 ), .pi01( pi111 ), .pi02( pi112 ), .pi03( pi113 ), .pi04( pi114 ), .pi05( pi238 ), .pi06( pi239 ), .pi07( pi240 ), .pi08( pi241 ), .pi09( pi242 ), .pi10( n44 ), .po0( tpo110 ), .po1( tpo111 ), .po2( tpo112 ), .po3( tpo113 ), .po4( tpo114 ), .po5( n45 ), .po6( n46 ) );
  adder_13 U13 ( .pi00( pi115 ), .pi01( pi116 ), .pi02( pi117 ), .pi03( pi118 ), .pi04( pi243 ), .pi05( pi244 ), .pi06( pi245 ), .pi07( pi246 ), .pi08( n45 ), .pi09( n46 ), .po0( tpo115 ), .po1( tpo116 ), .po2( tpo117 ), .po3( tpo118 ), .po4( n47 ), .po5( n48 ) );
  adder_14 U14 ( .pi00( pi018 ), .pi01( pi019 ), .pi02( pi020 ), .pi03( pi021 ), .pi04( pi146 ), .pi05( pi147 ), .pi06( pi148 ), .pi07( pi149 ), .pi08( n5 ), .pi09( n6 ), .po0( tpo018 ), .po1( tpo019 ), .po2( tpo020 ), .po3( tpo021 ), .po4( n7 ), .po5( n8 ) );
  adder_15 U15 ( .pi00( pi027 ), .pi01( pi028 ), .pi02( pi029 ), .pi03( pi030 ), .pi04( pi155 ), .pi05( pi156 ), .pi06( pi157 ), .pi07( pi158 ), .pi08( n9 ), .pi09( n10 ), .po0( tpo027 ), .po1( tpo028 ), .po2( tpo029 ), .po3( tpo030 ), .po4( n11 ), .po5( n12 ) );
  adder_16 U16 ( .pi00( pi022 ), .pi01( pi023 ), .pi02( pi024 ), .pi03( pi025 ), .pi04( pi026 ), .pi05( pi150 ), .pi06( pi151 ), .pi07( pi152 ), .pi08( pi153 ), .pi09( pi154 ), .pi10( n7 ), .pi11( n8 ), .po0( tpo022 ), .po1( tpo023 ), .po2( tpo024 ), .po3( tpo025 ), .po4( tpo026 ), .po5( n9 ), .po6( n10 ) );
  adder_17 U17 ( .pi00( pi013 ), .pi01( pi014 ), .pi02( pi015 ), .pi03( pi016 ), .pi04( pi017 ), .pi05( pi142 ), .pi06( pi143 ), .pi07( pi144 ), .pi08( pi145 ), .pi09( n3 ), .pi10( n4 ), .po0( tpo013 ), .po1( tpo014 ), .po2( tpo015 ), .po3( tpo016 ), .po4( tpo017 ), .po5( n5 ), .po6( n6 ) );
  adder_18 U18 ( .pi00( pi009 ), .pi01( pi010 ), .pi02( pi011 ), .pi03( pi012 ), .pi04( pi137 ), .pi05( pi138 ), .pi06( pi139 ), .pi07( pi140 ), .pi08( pi141 ), .pi09( n1 ), .pi10( n2 ), .po0( tpo009 ), .po1( tpo010 ), .po2( tpo011 ), .po3( tpo012 ), .po4( n3 ), .po5( n4 ) );
  adder_19 U19 ( .pi0( pi000 ), .pi1( pi001 ), .pi2( pi002 ), .pi3( pi128 ), .pi4( pi129 ), .pi5( pi130 ), .po0( tpo000 ), .po1( tpo001 ), .po2( tpo002 ), .po3( n0 ) );
  adder_20 U20 ( .pi00( pi003 ), .pi01( pi004 ), .pi02( pi005 ), .pi03( pi006 ), .pi04( pi007 ), .pi05( pi008 ), .pi06( pi131 ), .pi07( pi132 ), .pi08( pi133 ), .pi09( pi134 ), .pi10( pi135 ), .pi11( pi136 ), .pi12( n0 ), .po0( tpo003 ), .po1( tpo004 ), .po2( tpo005 ), .po3( tpo006 ), .po4( tpo007 ), .po5( tpo008 ), .po6( n1 ), .po7( n2 ) );
  adder_21 U21 ( .pi00( pi048 ), .pi01( pi049 ), .pi02( pi050 ), .pi03( pi051 ), .pi04( pi176 ), .pi05( pi177 ), .pi06( pi178 ), .pi07( pi179 ), .pi08( n19 ), .pi09( n20 ), .po0( tpo048 ), .po1( tpo049 ), .po2( tpo050 ), .po3( tpo051 ), .po4( n21 ), .po5( n22 ) );
  adder_22 U22 ( .pi00( pi056 ), .pi01( pi057 ), .pi02( pi058 ), .pi03( pi059 ), .pi04( pi060 ), .pi05( pi184 ), .pi06( pi185 ), .pi07( pi186 ), .pi08( pi187 ), .pi09( pi188 ), .pi10( n23 ), .pi11( n24 ), .po0( tpo056 ), .po1( tpo057 ), .po2( tpo058 ), .po3( tpo059 ), .po4( n25 ), .po5( tpo060 ) );
  adder_23 U23 ( .pi00( pi052 ), .pi01( pi053 ), .pi02( pi054 ), .pi03( pi055 ), .pi04( pi180 ), .pi05( pi181 ), .pi06( pi182 ), .pi07( pi183 ), .pi08( n21 ), .pi09( n22 ), .po0( tpo052 ), .po1( tpo053 ), .po2( tpo054 ), .po3( tpo055 ), .po4( n23 ), .po5( n24 ) );
  adder_24 U24 ( .pi00( pi039 ), .pi01( pi040 ), .pi02( pi041 ), .pi03( pi042 ), .pi04( pi168 ), .pi05( pi169 ), .pi06( pi170 ), .pi07( pi171 ), .pi08( n15 ), .pi09( n16 ), .po0( tpo039 ), .po1( tpo040 ), .po2( tpo041 ), .po3( tpo042 ), .po4( n17 ), .po5( n18 ) );
  adder_25 U25 ( .pi00( pi043 ), .pi01( pi044 ), .pi02( pi045 ), .pi03( pi046 ), .pi04( pi047 ), .pi05( pi172 ), .pi06( pi173 ), .pi07( pi174 ), .pi08( pi175 ), .pi09( n17 ), .pi10( n18 ), .po0( tpo043 ), .po1( tpo044 ), .po2( tpo045 ), .po3( tpo046 ), .po4( tpo047 ), .po5( n19 ), .po6( n20 ) );
  adder_26 U26 ( .pi00( pi035 ), .pi01( pi036 ), .pi02( pi037 ), .pi03( pi038 ), .pi04( pi163 ), .pi05( pi164 ), .pi06( pi165 ), .pi07( pi166 ), .pi08( pi167 ), .pi09( n13 ), .pi10( n14 ), .po0( tpo035 ), .po1( tpo036 ), .po2( tpo037 ), .po3( tpo038 ), .po4( n15 ), .po5( n16 ) );
  adder_27 U27 ( .pi00( pi031 ), .pi01( pi032 ), .pi02( pi033 ), .pi03( pi034 ), .pi04( pi159 ), .pi05( pi160 ), .pi06( pi161 ), .pi07( pi162 ), .pi08( n11 ), .pi09( n12 ), .po0( tpo031 ), .po1( tpo032 ), .po2( tpo033 ), .po3( tpo034 ), .po4( n13 ), .po5( n14 ) );
endmodule
