module mult16_15(pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 , po0 , po1 , po2 , po3 , po4 );
  input pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 ;
  output po0 , po1 , po2 , po3 , po4 ;
  wire new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36, new_n37, new_n38, new_n39, new_n40, new_n41, new_n42, new_n43, new_n44, new_n45, new_n46, new_n47, new_n48, new_n49, new_n50, new_n51, new_n52, new_n53, new_n54, new_n55, new_n56, new_n57, new_n58, new_n59, new_n60, new_n61, new_n62, new_n63, new_n64, new_n65, new_n66;
  assign new_n12 = ~pi03 & pi04 ;
  assign new_n13 = pi03 & ~pi04 ;
  assign new_n14 = ~new_n12 & ~new_n13 ;
  assign new_n15 = ~pi05 & pi06 ;
  assign new_n16 = pi05 & ~pi06 ;
  assign new_n17 = ~new_n15 & ~new_n16 ;
  assign new_n18 = new_n14 & new_n17 ;
  assign new_n19 = ~new_n14 & ~new_n17 ;
  assign new_n20 = ~new_n18 & ~new_n19 ;
  assign new_n21 = ~pi02 & new_n20 ;
  assign new_n22 = pi02 & ~new_n20 ;
  assign new_n23 = ~new_n21 & ~new_n22 ;
  assign new_n24 = pi00 & new_n23 ;
  assign new_n25 = ~pi00 & ~new_n23 ;
  assign new_n26 = ~new_n24 & ~new_n25 ;
  assign new_n27 = ~pi01 & new_n26 ;
  assign new_n28 = pi01 & ~new_n26 ;
  assign new_n29 = ~new_n27 & ~new_n28 ;
  assign new_n30 = ~new_n12 & ~new_n18 ;
  assign new_n31 = pi07 & ~new_n30 ;
  assign new_n32 = ~pi07 & new_n30 ;
  assign new_n33 = ~new_n31 & ~new_n32 ;
  assign new_n34 = new_n15 & new_n33 ;
  assign new_n35 = ~new_n15 & ~new_n33 ;
  assign new_n36 = ~new_n34 & ~new_n35 ;
  assign new_n37 = ~new_n21 & ~new_n24 ;
  assign new_n38 = new_n36 & ~new_n37 ;
  assign new_n39 = ~new_n36 & new_n37 ;
  assign new_n40 = ~new_n38 & ~new_n39 ;
  assign new_n41 = new_n27 & new_n40 ;
  assign new_n42 = ~new_n27 & ~new_n40 ;
  assign new_n43 = ~new_n41 & ~new_n42 ;
  assign new_n44 = ~pi08 & new_n43 ;
  assign new_n45 = pi08 & ~new_n43 ;
  assign new_n46 = ~new_n44 & ~new_n45 ;
  assign new_n47 = ~new_n31 & ~new_n34 ;
  assign new_n48 = pi09 & ~new_n47 ;
  assign new_n49 = ~pi09 & new_n47 ;
  assign new_n50 = ~new_n48 & ~new_n49 ;
  assign new_n51 = ~new_n44 & ~new_n50 ;
  assign new_n52 = new_n38 & ~new_n51 ;
  assign new_n53 = ~new_n41 & ~new_n44 ;
  assign new_n54 = new_n50 & ~new_n53 ;
  assign new_n55 = ~new_n50 & new_n53 ;
  assign new_n56 = ~new_n54 & ~new_n55 ;
  assign new_n57 = ~new_n38 & ~new_n56 ;
  assign new_n58 = ~new_n52 & ~new_n57 ;
  assign new_n59 = pi10 & new_n48 ;
  assign new_n60 = ~pi10 & ~new_n48 ;
  assign new_n61 = ~new_n59 & ~new_n60 ;
  assign new_n62 = ~new_n52 & ~new_n54 ;
  assign new_n63 = new_n61 & ~new_n62 ;
  assign new_n64 = ~new_n61 & new_n62 ;
  assign new_n65 = ~new_n63 & ~new_n64 ;
  assign new_n66 = ~new_n59 & ~new_n63 ;
  assign po0 = new_n29 ;
  assign po1 = new_n46 ;
  assign po2 = new_n58 ;
  assign po3 = new_n65 ;
  assign po4 = new_n66 ;
endmodule
