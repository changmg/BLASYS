module max_44_2(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 ;
  wire new_n9, new_n10, new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26;
  assign new_n9 = ~pi0 & pi2 ;
  assign new_n10 = ~pi7 & ~new_n9 ;
  assign new_n11 = pi1 & ~pi3 ;
  assign new_n12 = pi0 & ~pi2 ;
  assign new_n13 = ~new_n11 & ~new_n12 ;
  assign new_n14 = ~new_n10 & new_n13 ;
  assign new_n15 = ~pi1 & pi3 ;
  assign new_n16 = pi0 & pi4 ;
  assign new_n17 = pi2 & ~pi4 ;
  assign new_n18 = ~new_n16 & ~new_n17 ;
  assign new_n19 = pi1 & pi4 ;
  assign new_n20 = pi3 & ~pi4 ;
  assign new_n21 = ~new_n19 & ~new_n20 ;
  assign new_n22 = ~pi5 & new_n21 ;
  assign new_n23 = pi5 & ~new_n21 ;
  assign new_n24 = pi6 & ~new_n21 ;
  assign new_n25 = ~pi5 & ~pi6 ;
  assign new_n26 = ~new_n24 & ~new_n25 ;
  assign po0 = pi4 ;
  assign po1 = pi6 ;
  assign po2 = new_n14 ;
  assign po3 = new_n15 ;
  assign po4 = new_n18 ;
  assign po5 = new_n22 ;
  assign po6 = new_n23 ;
  assign po7 = new_n26 ;
endmodule
