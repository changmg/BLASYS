module mult16_10(pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , po00 , po01 , po02 , po03 , po04 , po05 , po06 , po07 , po08 , po09 , po10 , po11 , po12 , po13 , po14 , po15 );
  input pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 ;
  output po00 , po01 , po02 , po03 , po04 , po05 , po06 , po07 , po08 , po09 , po10 , po11 , po12 , po13 , po14 , po15 ;
  wire new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36, new_n37, new_n38, new_n39, new_n40, new_n41, new_n42, new_n43, new_n44, new_n45, new_n46, new_n47, new_n48, new_n49, new_n50, new_n51, new_n52, new_n53;
  assign new_n11 = pi00 & pi04 ;
  assign new_n12 = pi01 & pi05 ;
  assign new_n13 = new_n11 & new_n12 ;
  assign new_n14 = pi01 & pi04 ;
  assign new_n15 = pi00 & pi05 ;
  assign new_n16 = ~new_n14 & ~new_n15 ;
  assign new_n17 = ~new_n13 & ~new_n16 ;
  assign new_n18 = pi00 & pi06 ;
  assign new_n19 = pi02 & pi04 ;
  assign new_n20 = new_n12 & new_n19 ;
  assign new_n21 = ~new_n12 & ~new_n19 ;
  assign new_n22 = ~new_n20 & ~new_n21 ;
  assign new_n23 = new_n18 & new_n22 ;
  assign new_n24 = ~new_n18 & ~new_n22 ;
  assign new_n25 = ~new_n23 & ~new_n24 ;
  assign new_n26 = pi03 & pi05 ;
  assign new_n27 = pi01 & pi06 ;
  assign new_n28 = new_n19 & new_n26 ;
  assign new_n29 = pi03 & pi04 ;
  assign new_n30 = pi02 & pi05 ;
  assign new_n31 = ~new_n29 & ~new_n30 ;
  assign new_n32 = ~new_n28 & ~new_n31 ;
  assign new_n33 = new_n27 & new_n32 ;
  assign new_n34 = ~new_n27 & ~new_n32 ;
  assign new_n35 = ~new_n33 & ~new_n34 ;
  assign new_n36 = pi00 & pi07 ;
  assign new_n37 = ~new_n20 & ~new_n23 ;
  assign new_n38 = ~pi08 & ~new_n37 ;
  assign new_n39 = pi08 & new_n37 ;
  assign new_n40 = ~new_n38 & ~new_n39 ;
  assign new_n41 = new_n36 & new_n40 ;
  assign new_n42 = ~new_n36 & ~new_n40 ;
  assign new_n43 = ~new_n41 & ~new_n42 ;
  assign new_n44 = ~new_n38 & ~new_n41 ;
  assign new_n45 = pi01 & pi07 ;
  assign new_n46 = ~new_n28 & ~new_n33 ;
  assign new_n47 = ~pi09 & ~new_n46 ;
  assign new_n48 = pi09 & new_n46 ;
  assign new_n49 = ~new_n47 & ~new_n48 ;
  assign new_n50 = new_n45 & new_n49 ;
  assign new_n51 = ~new_n45 & ~new_n49 ;
  assign new_n52 = ~new_n50 & ~new_n51 ;
  assign new_n53 = ~new_n47 & ~new_n50 ;
  assign po00 = pi01 ;
  assign po01 = pi03 ;
  assign po02 = pi04 ;
  assign po03 = pi05 ;
  assign po04 = pi06 ;
  assign po05 = pi07 ;
  assign po06 = new_n11 ;
  assign po07 = new_n13 ;
  assign po08 = new_n17 ;
  assign po09 = new_n25 ;
  assign po10 = new_n26 ;
  assign po11 = new_n35 ;
  assign po12 = new_n43 ;
  assign po13 = new_n44 ;
  assign po14 = new_n52 ;
  assign po15 = new_n53 ;
endmodule
