module mult8_12(pi0 , pi1 , pi2 , pi3 , pi4 , po0 , po1 , po2 );
  input pi0 , pi1 , pi2 , pi3 , pi4 ;
  output po0 , po1 , po2 ;
  wire new_n6, new_n7, new_n8, new_n9, new_n10, new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24;
  assign new_n6 = pi1 & ~pi2 ;
  assign new_n7 = ~pi1 & pi2 ;
  assign new_n8 = ~new_n6 & ~new_n7 ;
  assign new_n9 = ~pi3 & ~new_n8 ;
  assign new_n10 = ~pi1 & ~pi2 ;
  assign new_n11 = pi1 & pi2 ;
  assign new_n12 = ~new_n10 & ~new_n11 ;
  assign new_n13 = pi3 & ~new_n12 ;
  assign new_n14 = ~new_n9 & ~new_n13 ;
  assign new_n15 = ~pi4 & new_n14 ;
  assign new_n16 = pi4 & ~new_n14 ;
  assign new_n17 = ~new_n15 & ~new_n16 ;
  assign new_n18 = ~pi0 & ~new_n17 ;
  assign new_n19 = ~pi4 & ~new_n14 ;
  assign new_n20 = pi4 & new_n14 ;
  assign new_n21 = ~new_n19 & ~new_n20 ;
  assign new_n22 = pi0 & ~new_n21 ;
  assign new_n23 = pi4 & ~new_n13 ;
  assign new_n24 = ~new_n9 & ~new_n23 ;
  assign po0 = new_n18 ;
  assign po1 = new_n22 ;
  assign po2 = new_n24 ;
endmodule
