module mac_0_tb;
reg [4:0] pi;
wire [2:0] po;
mac_0 dut(pi[4], pi[3], pi[2], pi[1], pi[0], po[2], po[1], po[0]);
initial
begin
# 1  pi=5'b00000;
#1 $display("%b", po);
# 1  pi=5'b00001;
#1 $display("%b", po);
# 1  pi=5'b00010;
#1 $display("%b", po);
# 1  pi=5'b00011;
#1 $display("%b", po);
# 1  pi=5'b00100;
#1 $display("%b", po);
# 1  pi=5'b00101;
#1 $display("%b", po);
# 1  pi=5'b00110;
#1 $display("%b", po);
# 1  pi=5'b00111;
#1 $display("%b", po);
# 1  pi=5'b01000;
#1 $display("%b", po);
# 1  pi=5'b01001;
#1 $display("%b", po);
# 1  pi=5'b01010;
#1 $display("%b", po);
# 1  pi=5'b01011;
#1 $display("%b", po);
# 1  pi=5'b01100;
#1 $display("%b", po);
# 1  pi=5'b01101;
#1 $display("%b", po);
# 1  pi=5'b01110;
#1 $display("%b", po);
# 1  pi=5'b01111;
#1 $display("%b", po);
# 1  pi=5'b10000;
#1 $display("%b", po);
# 1  pi=5'b10001;
#1 $display("%b", po);
# 1  pi=5'b10010;
#1 $display("%b", po);
# 1  pi=5'b10011;
#1 $display("%b", po);
# 1  pi=5'b10100;
#1 $display("%b", po);
# 1  pi=5'b10101;
#1 $display("%b", po);
# 1  pi=5'b10110;
#1 $display("%b", po);
# 1  pi=5'b10111;
#1 $display("%b", po);
# 1  pi=5'b11000;
#1 $display("%b", po);
# 1  pi=5'b11001;
#1 $display("%b", po);
# 1  pi=5'b11010;
#1 $display("%b", po);
# 1  pi=5'b11011;
#1 $display("%b", po);
# 1  pi=5'b11100;
#1 $display("%b", po);
# 1  pi=5'b11101;
#1 $display("%b", po);
# 1  pi=5'b11110;
#1 $display("%b", po);
# 1  pi=5'b11111;
#1 $display("%b", po);
end
endmodule
