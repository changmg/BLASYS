module max_28_1(pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , po0 , po1 , po2 , po3 , po4 , po5 );
  input pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 ;
  output po0 , po1 , po2 , po3 , po4 , po5 ;
  wire new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31;
  assign new_n11 = ~pi01 & pi03 ;
  assign new_n12 = ~pi06 & ~new_n11 ;
  assign new_n13 = ~pi00 & pi02 ;
  assign new_n14 = ~pi07 & ~new_n13 ;
  assign new_n15 = new_n12 & new_n14 ;
  assign new_n16 = ~pi04 & new_n15 ;
  assign new_n17 = pi00 & ~pi02 ;
  assign new_n18 = pi01 & ~pi03 ;
  assign new_n19 = ~new_n17 & ~new_n18 ;
  assign new_n20 = new_n12 & ~new_n19 ;
  assign new_n21 = pi00 & pi08 ;
  assign new_n22 = pi02 & ~pi08 ;
  assign new_n23 = ~new_n21 & ~new_n22 ;
  assign new_n24 = pi01 & pi08 ;
  assign new_n25 = pi03 & ~pi08 ;
  assign new_n26 = ~new_n24 & ~new_n25 ;
  assign new_n27 = ~pi05 & new_n26 ;
  assign new_n28 = pi05 & ~new_n26 ;
  assign new_n29 = ~pi05 & pi09 ;
  assign new_n30 = ~pi09 & ~new_n26 ;
  assign new_n31 = ~new_n29 & ~new_n30 ;
  assign po0 = new_n16 ;
  assign po1 = new_n20 ;
  assign po2 = new_n23 ;
  assign po3 = new_n27 ;
  assign po4 = new_n28 ;
  assign po5 = new_n31 ;
endmodule
