module max_63_0(pi0 , pi1 , pi2 , pi3 , pi4 , po0 , po1 , po2 , po3 , po4 , po5 , po6 );
  input pi0 , pi1 , pi2 , pi3 , pi4 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 ;
  wire new_n6, new_n7, new_n8, new_n9, new_n10, new_n11, new_n12, new_n13, new_n14, new_n15;
  assign new_n6 = pi0 & ~pi1 ;
  assign new_n7 = ~pi0 & pi1 ;
  assign new_n8 = pi0 & pi2 ;
  assign new_n9 = pi1 & ~pi2 ;
  assign new_n10 = ~new_n8 & ~new_n9 ;
  assign new_n11 = ~pi3 & new_n10 ;
  assign new_n12 = pi3 & ~new_n10 ;
  assign new_n13 = ~pi3 & pi4 ;
  assign new_n14 = ~pi4 & ~new_n10 ;
  assign new_n15 = ~new_n13 & ~new_n14 ;
  assign po0 = pi2 ;
  assign po1 = pi4 ;
  assign po2 = new_n6 ;
  assign po3 = new_n7 ;
  assign po4 = new_n11 ;
  assign po5 = new_n12 ;
  assign po6 = new_n15 ;
endmodule
