module mult16_12(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , po00 , po01 , po02 , po03 , po04 , po05 , po06 , po07 , po08 , po09 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ;
  output po00 , po01 , po02 , po03 , po04 , po05 , po06 , po07 , po08 , po09 ;
  wire new_n9, new_n10, new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33;
  assign new_n9 = pi1 & pi4 ;
  assign new_n10 = pi0 & pi6 ;
  assign new_n11 = pi2 & pi5 ;
  assign new_n12 = new_n9 & new_n11 ;
  assign new_n13 = pi2 & pi4 ;
  assign new_n14 = pi1 & pi5 ;
  assign new_n15 = ~new_n13 & ~new_n14 ;
  assign new_n16 = ~new_n12 & ~new_n15 ;
  assign new_n17 = new_n10 & new_n16 ;
  assign new_n18 = ~new_n10 & ~new_n16 ;
  assign new_n19 = ~new_n17 & ~new_n18 ;
  assign new_n20 = pi3 & pi4 ;
  assign new_n21 = ~new_n12 & ~new_n17 ;
  assign new_n22 = pi1 & pi6 ;
  assign new_n23 = new_n11 & new_n20 ;
  assign new_n24 = ~new_n11 & ~new_n20 ;
  assign new_n25 = ~new_n23 & ~new_n24 ;
  assign new_n26 = new_n22 & new_n25 ;
  assign new_n27 = ~new_n22 & ~new_n25 ;
  assign new_n28 = ~new_n26 & ~new_n27 ;
  assign new_n29 = ~new_n21 & new_n28 ;
  assign new_n30 = new_n21 & ~new_n28 ;
  assign new_n31 = ~new_n29 & ~new_n30 ;
  assign new_n32 = ~pi7 & ~new_n29 ;
  assign new_n33 = ~new_n23 & ~new_n26 ;
  assign po00 = pi1 ;
  assign po01 = pi4 ;
  assign po02 = pi5 ;
  assign po03 = pi6 ;
  assign po04 = new_n9 ;
  assign po05 = new_n19 ;
  assign po06 = new_n20 ;
  assign po07 = new_n31 ;
  assign po08 = new_n32 ;
  assign po09 = new_n33 ;
endmodule
