module max_1_2(pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , po0 , po1 , po2 , po3 );
  input pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 ;
  output po0 , po1 , po2 , po3 ;
  wire new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29;
  assign new_n11 = ~pi01 & pi03 ;
  assign new_n12 = ~pi00 & pi02 ;
  assign new_n13 = ~pi07 & ~new_n12 ;
  assign new_n14 = ~pi05 & ~pi08 ;
  assign new_n15 = new_n13 & new_n14 ;
  assign new_n16 = ~pi04 & new_n15 ;
  assign new_n17 = ~pi09 & new_n13 ;
  assign new_n18 = pi00 & ~pi02 ;
  assign new_n19 = pi01 & ~pi03 ;
  assign new_n20 = ~new_n18 & ~new_n19 ;
  assign new_n21 = ~new_n17 & new_n20 ;
  assign new_n22 = ~new_n16 & new_n21 ;
  assign new_n23 = ~new_n11 & ~new_n22 ;
  assign new_n24 = pi00 & pi06 ;
  assign new_n25 = pi02 & ~pi06 ;
  assign new_n26 = ~new_n24 & ~new_n25 ;
  assign new_n27 = pi01 & pi06 ;
  assign new_n28 = pi03 & ~pi06 ;
  assign new_n29 = ~new_n27 & ~new_n28 ;
  assign po0 = pi06 ;
  assign po1 = new_n23 ;
  assign po2 = new_n26 ;
  assign po3 = new_n29 ;
endmodule
