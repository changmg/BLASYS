// Benchmark "c1908" written by ABC on Thu Jul 14 21:13:58 2022

module c1908 ( 
    G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
    G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237,
    G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_new_n59__, new_new_n60__, new_new_n61__, new_new_n62__,
    new_new_n63__, new_new_n64__, new_new_n65__, new_new_n66__,
    new_new_n67__, new_new_n68__, new_new_n69__, new_new_n70__,
    new_new_n71__, new_new_n72__, new_new_n73__, new_new_n74__,
    new_new_n75__, new_new_n76__, new_new_n77__, new_new_n78__,
    new_new_n79__, new_new_n80__, new_new_n81__, new_new_n82__,
    new_new_n83__, new_new_n84__, new_new_n85__, new_new_n86__,
    new_new_n87__, new_new_n88__, new_new_n89__, new_new_n90__,
    new_new_n91__, new_new_n92__, new_new_n93__, new_new_n94__,
    new_new_n95__, new_new_n96__, new_new_n97__, new_new_n98__,
    new_new_n99__, new_new_n100__, new_new_n101__, new_new_n102__,
    new_new_n103__, new_new_n104__, new_new_n105__, new_new_n106__,
    new_new_n107__, new_new_n108__, new_new_n109__, new_new_n110__,
    new_new_n111__, new_new_n112__, new_new_n113__, new_new_n114__,
    new_new_n115__, new_new_n116__, new_new_n117__, new_new_n118__,
    new_new_n119__, new_new_n120__, new_new_n121__, new_new_n122__,
    new_new_n123__, new_new_n124__, new_new_n125__, new_new_n126__,
    new_new_n127__, new_new_n128__, new_new_n129__, new_new_n130__,
    new_new_n131__, new_new_n132__, new_new_n133__, new_new_n134__,
    new_new_n135__, new_new_n136__, new_new_n137__, new_new_n138__,
    new_new_n139__, new_new_n140__, new_new_n141__, new_new_n142__,
    new_new_n143__, new_new_n144__, new_new_n145__, new_new_n146__,
    new_new_n147__, new_new_n148__, new_new_n149__, new_new_n150__,
    new_new_n151__, new_new_n152__, new_new_n153__, new_new_n154__,
    new_new_n155__, new_new_n156__, new_new_n157__, new_new_n158__,
    new_new_n159__, new_new_n160__, new_new_n161__, new_new_n162__,
    new_new_n163__, new_new_n164__, new_new_n165__, new_new_n166__,
    new_new_n167__, new_new_n168__, new_new_n169__, new_new_n170__,
    new_new_n171__, new_new_n172__, new_new_n173__, new_new_n174__,
    new_new_n175__, new_new_n176__, new_new_n177__, new_new_n178__,
    new_new_n179__, new_new_n180__, new_new_n181__, new_new_n182__,
    new_new_n183__, new_new_n184__, new_new_n185__, new_new_n186__,
    new_new_n187__, new_new_n188__, new_new_n189__, new_new_n190__,
    new_new_n191__, new_new_n192__, new_new_n193__, new_new_n194__,
    new_new_n195__, new_new_n196__, new_new_n197__, new_new_n198__,
    new_new_n199__, new_new_n200__, new_new_n201__, new_new_n202__,
    new_new_n203__, new_new_n204__, new_new_n205__, new_new_n206__,
    new_new_n207__, new_new_n208__, new_new_n209__, new_new_n210__,
    new_new_n211__, new_new_n212__, new_new_n213__, new_new_n214__,
    new_new_n215__, new_new_n216__, new_new_n217__, new_new_n218__,
    new_new_n219__, new_new_n220__, new_new_n221__, new_new_n222__,
    new_new_n223__, new_new_n224__, new_new_n225__, new_new_n226__,
    new_new_n227__, new_new_n228__, new_new_n229__, new_new_n230__,
    new_new_n231__, new_new_n232__, new_new_n233__, new_new_n234__,
    new_new_n235__, new_new_n236__, new_new_n237__, new_new_n238__,
    new_new_n240__, new_new_n241__, new_new_n242__, new_new_n243__,
    new_new_n244__, new_new_n245__, new_new_n246__, new_new_n248__,
    new_new_n249__, new_new_n250__, new_new_n251__, new_new_n252__,
    new_new_n254__, new_new_n255__, new_new_n256__, new_new_n257__,
    new_new_n258__, new_new_n259__, new_new_n261__, new_new_n262__,
    new_new_n263__, new_new_n264__, new_new_n265__, new_new_n266__,
    new_new_n267__, new_new_n268__, new_new_n269__, new_new_n271__,
    new_new_n272__, new_new_n273__, new_new_n274__, new_new_n275__,
    new_new_n277__, new_new_n278__, new_new_n279__, new_new_n280__,
    new_new_n282__, new_new_n283__, new_new_n284__, new_new_n285__,
    new_new_n286__, new_new_n287__, new_new_n289__, new_new_n290__,
    new_new_n291__, new_new_n293__, new_new_n294__, new_new_n295__,
    new_new_n296__, new_new_n298__, new_new_n299__, new_new_n300__,
    new_new_n301__, new_new_n302__, new_new_n304__, new_new_n305__,
    new_new_n306__, new_new_n307__, new_new_n309__, new_new_n310__,
    new_new_n311__, new_new_n312__, new_new_n313__, new_new_n314__,
    new_new_n316__, new_new_n317__, new_new_n318__, new_new_n320__,
    new_new_n321__, new_new_n322__, new_new_n323__, new_new_n324__,
    new_new_n326__, new_new_n327__, new_new_n328__, new_new_n330__,
    new_new_n331__, new_new_n332__, new_new_n333__, new_new_n334__,
    new_new_n335__, new_new_n336__, new_new_n337__, new_new_n338__,
    new_new_n339__, new_new_n340__, new_new_n341__, new_new_n342__,
    new_new_n343__, new_new_n344__, new_new_n345__, new_new_n346__,
    new_new_n347__, new_new_n348__, new_new_n349__, new_new_n350__,
    new_new_n351__, new_new_n352__, new_new_n353__, new_new_n354__,
    new_new_n355__, new_new_n356__, new_new_n357__, new_new_n358__,
    new_new_n359__, new_new_n360__, new_new_n361__, new_new_n362__,
    new_new_n363__, new_new_n364__, new_new_n365__, new_new_n366__,
    new_new_n367__, new_new_n368__, new_new_n369__, new_new_n371__,
    new_new_n372__, new_new_n373__, new_new_n374__, new_new_n375__,
    new_new_n376__, new_new_n378__, new_new_n379__, new_new_n380__,
    new_new_n381__, new_new_n382__, new_new_n384__, new_new_n385__,
    new_new_n386__, new_new_n387__, new_new_n388__, new_new_n390__,
    new_new_n391__, new_new_n392__, new_new_n393__, new_new_n394__,
    new_new_n396__, new_new_n397__, new_new_n398__, new_new_n399__,
    new_new_n400__, new_new_n402__, new_new_n403__, new_new_n404__,
    new_new_n405__, new_new_n406__, new_new_n407__, new_new_n409__,
    new_new_n410__, new_new_n411__, new_new_n412__, new_new_n413__,
    new_new_n414__, new_new_n415__, new_new_n416__, new_new_n417__,
    new_new_n418__, new_new_n420__, new_new_n421__, new_new_n422__,
    new_new_n423__, new_new_n424__;
  assign new_new_n59__ = ~G125 & ~G140;
  assign new_new_n60__ = G125 & G140;
  assign new_new_n61__ = ~new_new_n59__ & ~new_new_n60__;
  assign new_new_n62__ = G146 & ~new_new_n61__;
  assign new_new_n63__ = ~G146 & new_new_n61__;
  assign new_new_n64__ = ~new_new_n62__ & ~new_new_n63__;
  assign new_new_n65__ = G221 & G234;
  assign new_new_n66__ = ~G953 & new_new_n65__;
  assign new_new_n67__ = G137 & new_new_n66__;
  assign new_new_n68__ = ~G137 & ~new_new_n66__;
  assign new_new_n69__ = ~new_new_n67__ & ~new_new_n68__;
  assign new_new_n70__ = G119 & ~G128;
  assign new_new_n71__ = ~G119 & G128;
  assign new_new_n72__ = ~new_new_n70__ & ~new_new_n71__;
  assign new_new_n73__ = new_new_n69__ & new_new_n72__;
  assign new_new_n74__ = ~new_new_n69__ & ~new_new_n72__;
  assign new_new_n75__ = ~new_new_n73__ & ~new_new_n74__;
  assign new_new_n76__ = G110 & ~new_new_n75__;
  assign new_new_n77__ = ~G110 & new_new_n75__;
  assign new_new_n78__ = ~new_new_n76__ & ~new_new_n77__;
  assign new_new_n79__ = new_new_n64__ & new_new_n78__;
  assign new_new_n80__ = ~new_new_n64__ & ~new_new_n78__;
  assign new_new_n81__ = ~new_new_n79__ & ~new_new_n80__;
  assign new_new_n82__ = ~G902 & ~new_new_n81__;
  assign new_new_n83__ = G234 & ~G902;
  assign new_new_n84__ = G217 & ~new_new_n83__;
  assign new_new_n85__ = ~new_new_n82__ & new_new_n84__;
  assign new_new_n86__ = new_new_n82__ & ~new_new_n84__;
  assign new_new_n87__ = ~new_new_n85__ & ~new_new_n86__;
  assign new_new_n88__ = ~G134 & ~G137;
  assign new_new_n89__ = G134 & G137;
  assign new_new_n90__ = ~new_new_n88__ & ~new_new_n89__;
  assign new_new_n91__ = ~G143 & ~G146;
  assign new_new_n92__ = G143 & G146;
  assign new_new_n93__ = ~new_new_n91__ & ~new_new_n92__;
  assign new_new_n94__ = G128 & new_new_n93__;
  assign new_new_n95__ = ~G128 & ~new_new_n93__;
  assign new_new_n96__ = ~new_new_n94__ & ~new_new_n95__;
  assign new_new_n97__ = G131 & ~new_new_n96__;
  assign new_new_n98__ = ~G131 & new_new_n96__;
  assign new_new_n99__ = ~new_new_n97__ & ~new_new_n98__;
  assign new_new_n100__ = new_new_n90__ & new_new_n99__;
  assign new_new_n101__ = ~new_new_n90__ & ~new_new_n99__;
  assign new_new_n102__ = ~new_new_n100__ & ~new_new_n101__;
  assign new_new_n103__ = ~G116 & ~G119;
  assign new_new_n104__ = G116 & G119;
  assign new_new_n105__ = ~new_new_n103__ & ~new_new_n104__;
  assign new_new_n106__ = G113 & new_new_n105__;
  assign new_new_n107__ = ~G113 & ~new_new_n105__;
  assign new_new_n108__ = ~new_new_n106__ & ~new_new_n107__;
  assign new_new_n109__ = G210 & ~G237;
  assign new_new_n110__ = ~G953 & new_new_n109__;
  assign new_new_n111__ = G101 & ~new_new_n110__;
  assign new_new_n112__ = ~G101 & new_new_n110__;
  assign new_new_n113__ = ~new_new_n111__ & ~new_new_n112__;
  assign new_new_n114__ = new_new_n108__ & ~new_new_n113__;
  assign new_new_n115__ = ~new_new_n108__ & new_new_n113__;
  assign new_new_n116__ = ~new_new_n114__ & ~new_new_n115__;
  assign new_new_n117__ = new_new_n102__ & new_new_n116__;
  assign new_new_n118__ = ~new_new_n102__ & ~new_new_n116__;
  assign new_new_n119__ = ~new_new_n117__ & ~new_new_n118__;
  assign new_new_n120__ = ~G902 & ~new_new_n119__;
  assign new_new_n121__ = G472 & ~new_new_n120__;
  assign new_new_n122__ = ~G472 & new_new_n120__;
  assign new_new_n123__ = ~new_new_n121__ & ~new_new_n122__;
  assign new_new_n124__ = new_new_n87__ & ~new_new_n123__;
  assign new_new_n125__ = ~G237 & ~G902;
  assign new_new_n126__ = G214 & ~new_new_n125__;
  assign new_new_n127__ = G210 & ~new_new_n125__;
  assign new_new_n128__ = G110 & ~G122;
  assign new_new_n129__ = ~G110 & G122;
  assign new_new_n130__ = ~new_new_n128__ & ~new_new_n129__;
  assign new_new_n131__ = ~G104 & ~G107;
  assign new_new_n132__ = G104 & G107;
  assign new_new_n133__ = ~new_new_n131__ & ~new_new_n132__;
  assign new_new_n134__ = G101 & new_new_n133__;
  assign new_new_n135__ = ~G101 & ~new_new_n133__;
  assign new_new_n136__ = ~new_new_n134__ & ~new_new_n135__;
  assign new_new_n137__ = new_new_n108__ & ~new_new_n136__;
  assign new_new_n138__ = ~new_new_n108__ & new_new_n136__;
  assign new_new_n139__ = ~new_new_n137__ & ~new_new_n138__;
  assign new_new_n140__ = new_new_n130__ & new_new_n139__;
  assign new_new_n141__ = ~new_new_n130__ & ~new_new_n139__;
  assign new_new_n142__ = ~new_new_n140__ & ~new_new_n141__;
  assign new_new_n143__ = G224 & ~G953;
  assign new_new_n144__ = G125 & ~new_new_n96__;
  assign new_new_n145__ = ~G125 & new_new_n96__;
  assign new_new_n146__ = ~new_new_n144__ & ~new_new_n145__;
  assign new_new_n147__ = new_new_n143__ & ~new_new_n146__;
  assign new_new_n148__ = ~new_new_n143__ & new_new_n146__;
  assign new_new_n149__ = ~new_new_n147__ & ~new_new_n148__;
  assign new_new_n150__ = new_new_n142__ & new_new_n149__;
  assign new_new_n151__ = ~new_new_n142__ & ~new_new_n149__;
  assign new_new_n152__ = ~new_new_n150__ & ~new_new_n151__;
  assign new_new_n153__ = ~G902 & new_new_n152__;
  assign new_new_n154__ = ~new_new_n127__ & new_new_n153__;
  assign new_new_n155__ = new_new_n127__ & ~new_new_n153__;
  assign new_new_n156__ = ~new_new_n154__ & ~new_new_n155__;
  assign new_new_n157__ = ~new_new_n126__ & ~new_new_n156__;
  assign new_new_n158__ = G221 & ~new_new_n83__;
  assign new_new_n159__ = ~G110 & ~G140;
  assign new_new_n160__ = G110 & G140;
  assign new_new_n161__ = ~new_new_n159__ & ~new_new_n160__;
  assign new_new_n162__ = G227 & ~G953;
  assign new_new_n163__ = new_new_n136__ & ~new_new_n162__;
  assign new_new_n164__ = ~new_new_n136__ & new_new_n162__;
  assign new_new_n165__ = ~new_new_n163__ & ~new_new_n164__;
  assign new_new_n166__ = new_new_n161__ & ~new_new_n165__;
  assign new_new_n167__ = ~new_new_n161__ & new_new_n165__;
  assign new_new_n168__ = ~new_new_n166__ & ~new_new_n167__;
  assign new_new_n169__ = new_new_n102__ & new_new_n168__;
  assign new_new_n170__ = ~new_new_n102__ & ~new_new_n168__;
  assign new_new_n171__ = ~new_new_n169__ & ~new_new_n170__;
  assign new_new_n172__ = ~G902 & ~new_new_n171__;
  assign new_new_n173__ = G469 & ~new_new_n172__;
  assign new_new_n174__ = ~G469 & new_new_n172__;
  assign new_new_n175__ = ~new_new_n173__ & ~new_new_n174__;
  assign new_new_n176__ = ~new_new_n158__ & ~new_new_n175__;
  assign new_new_n177__ = new_new_n157__ & new_new_n176__;
  assign new_new_n178__ = new_new_n124__ & new_new_n177__;
  assign new_new_n179__ = G128 & ~G143;
  assign new_new_n180__ = ~G128 & G143;
  assign new_new_n181__ = ~new_new_n179__ & ~new_new_n180__;
  assign new_new_n182__ = G217 & G234;
  assign new_new_n183__ = ~G953 & new_new_n182__;
  assign new_new_n184__ = ~G116 & ~G122;
  assign new_new_n185__ = G116 & G122;
  assign new_new_n186__ = ~new_new_n184__ & ~new_new_n185__;
  assign new_new_n187__ = G107 & ~G134;
  assign new_new_n188__ = ~G107 & G134;
  assign new_new_n189__ = ~new_new_n187__ & ~new_new_n188__;
  assign new_new_n190__ = new_new_n186__ & new_new_n189__;
  assign new_new_n191__ = ~new_new_n186__ & ~new_new_n189__;
  assign new_new_n192__ = ~new_new_n190__ & ~new_new_n191__;
  assign new_new_n193__ = new_new_n183__ & ~new_new_n192__;
  assign new_new_n194__ = ~new_new_n183__ & new_new_n192__;
  assign new_new_n195__ = ~new_new_n193__ & ~new_new_n194__;
  assign new_new_n196__ = new_new_n181__ & new_new_n195__;
  assign new_new_n197__ = ~new_new_n181__ & ~new_new_n195__;
  assign new_new_n198__ = ~new_new_n196__ & ~new_new_n197__;
  assign new_new_n199__ = ~G902 & ~new_new_n198__;
  assign new_new_n200__ = G478 & ~new_new_n199__;
  assign new_new_n201__ = ~G478 & new_new_n199__;
  assign new_new_n202__ = ~new_new_n200__ & ~new_new_n201__;
  assign new_new_n203__ = G131 & ~G143;
  assign new_new_n204__ = ~G131 & G143;
  assign new_new_n205__ = ~new_new_n203__ & ~new_new_n204__;
  assign new_new_n206__ = G214 & ~G237;
  assign new_new_n207__ = ~G953 & new_new_n206__;
  assign new_new_n208__ = ~new_new_n64__ & ~new_new_n207__;
  assign new_new_n209__ = new_new_n64__ & new_new_n207__;
  assign new_new_n210__ = ~new_new_n208__ & ~new_new_n209__;
  assign new_new_n211__ = ~G113 & ~G122;
  assign new_new_n212__ = G113 & G122;
  assign new_new_n213__ = ~new_new_n211__ & ~new_new_n212__;
  assign new_new_n214__ = G104 & new_new_n213__;
  assign new_new_n215__ = ~G104 & ~new_new_n213__;
  assign new_new_n216__ = ~new_new_n214__ & ~new_new_n215__;
  assign new_new_n217__ = new_new_n210__ & ~new_new_n216__;
  assign new_new_n218__ = ~new_new_n210__ & new_new_n216__;
  assign new_new_n219__ = ~new_new_n217__ & ~new_new_n218__;
  assign new_new_n220__ = new_new_n205__ & new_new_n219__;
  assign new_new_n221__ = ~new_new_n205__ & ~new_new_n219__;
  assign new_new_n222__ = ~new_new_n220__ & ~new_new_n221__;
  assign new_new_n223__ = ~G902 & ~new_new_n222__;
  assign new_new_n224__ = G475 & ~new_new_n223__;
  assign new_new_n225__ = ~G475 & new_new_n223__;
  assign new_new_n226__ = ~new_new_n224__ & ~new_new_n225__;
  assign new_new_n227__ = new_new_n202__ & new_new_n226__;
  assign new_new_n228__ = ~G898 & G953;
  assign new_new_n229__ = G234 & G237;
  assign new_new_n230__ = G902 & ~new_new_n229__;
  assign new_new_n231__ = new_new_n228__ & new_new_n230__;
  assign new_new_n232__ = G952 & ~G953;
  assign new_new_n233__ = ~new_new_n229__ & new_new_n232__;
  assign new_new_n234__ = ~new_new_n231__ & ~new_new_n233__;
  assign new_new_n235__ = new_new_n227__ & ~new_new_n234__;
  assign new_new_n236__ = new_new_n178__ & new_new_n235__;
  assign new_new_n237__ = ~G101 & ~new_new_n236__;
  assign new_new_n238__ = G101 & new_new_n236__;
  assign G3 = ~new_new_n237__ & ~new_new_n238__;
  assign new_new_n240__ = new_new_n87__ & new_new_n123__;
  assign new_new_n241__ = new_new_n177__ & new_new_n240__;
  assign new_new_n242__ = new_new_n202__ & ~new_new_n226__;
  assign new_new_n243__ = ~new_new_n234__ & new_new_n242__;
  assign new_new_n244__ = new_new_n241__ & new_new_n243__;
  assign new_new_n245__ = ~G104 & ~new_new_n244__;
  assign new_new_n246__ = G104 & new_new_n244__;
  assign G6 = ~new_new_n245__ & ~new_new_n246__;
  assign new_new_n248__ = ~new_new_n202__ & new_new_n226__;
  assign new_new_n249__ = ~new_new_n234__ & new_new_n248__;
  assign new_new_n250__ = new_new_n241__ & new_new_n249__;
  assign new_new_n251__ = ~G107 & ~new_new_n250__;
  assign new_new_n252__ = G107 & new_new_n250__;
  assign G9 = ~new_new_n251__ & ~new_new_n252__;
  assign new_new_n254__ = ~new_new_n87__ & new_new_n123__;
  assign new_new_n255__ = new_new_n227__ & new_new_n254__;
  assign new_new_n256__ = new_new_n177__ & ~new_new_n234__;
  assign new_new_n257__ = new_new_n255__ & new_new_n256__;
  assign new_new_n258__ = ~G110 & ~new_new_n257__;
  assign new_new_n259__ = G110 & new_new_n257__;
  assign G12 = ~new_new_n258__ & ~new_new_n259__;
  assign new_new_n261__ = ~new_new_n87__ & ~new_new_n123__;
  assign new_new_n262__ = new_new_n177__ & new_new_n261__;
  assign new_new_n263__ = ~G900 & G953;
  assign new_new_n264__ = new_new_n230__ & new_new_n263__;
  assign new_new_n265__ = ~new_new_n233__ & ~new_new_n264__;
  assign new_new_n266__ = new_new_n248__ & ~new_new_n265__;
  assign new_new_n267__ = new_new_n262__ & new_new_n266__;
  assign new_new_n268__ = ~G128 & ~new_new_n267__;
  assign new_new_n269__ = G128 & new_new_n267__;
  assign G30 = ~new_new_n268__ & ~new_new_n269__;
  assign new_new_n271__ = ~new_new_n202__ & ~new_new_n226__;
  assign new_new_n272__ = ~new_new_n265__ & new_new_n271__;
  assign new_new_n273__ = new_new_n178__ & new_new_n272__;
  assign new_new_n274__ = ~G143 & ~new_new_n273__;
  assign new_new_n275__ = G143 & new_new_n273__;
  assign G45 = ~new_new_n274__ & ~new_new_n275__;
  assign new_new_n277__ = new_new_n242__ & ~new_new_n265__;
  assign new_new_n278__ = new_new_n262__ & new_new_n277__;
  assign new_new_n279__ = ~G146 & ~new_new_n278__;
  assign new_new_n280__ = G146 & new_new_n278__;
  assign G48 = ~new_new_n279__ & ~new_new_n280__;
  assign new_new_n282__ = ~new_new_n158__ & new_new_n175__;
  assign new_new_n283__ = new_new_n157__ & new_new_n282__;
  assign new_new_n284__ = new_new_n124__ & new_new_n283__;
  assign new_new_n285__ = new_new_n243__ & new_new_n284__;
  assign new_new_n286__ = ~G113 & ~new_new_n285__;
  assign new_new_n287__ = G113 & new_new_n285__;
  assign G15 = ~new_new_n286__ & ~new_new_n287__;
  assign new_new_n289__ = new_new_n249__ & new_new_n284__;
  assign new_new_n290__ = ~G116 & ~new_new_n289__;
  assign new_new_n291__ = G116 & new_new_n289__;
  assign G18 = ~new_new_n290__ & ~new_new_n291__;
  assign new_new_n293__ = new_new_n235__ & new_new_n261__;
  assign new_new_n294__ = new_new_n283__ & new_new_n293__;
  assign new_new_n295__ = ~G119 & ~new_new_n294__;
  assign new_new_n296__ = G119 & new_new_n294__;
  assign G21 = ~new_new_n295__ & ~new_new_n296__;
  assign new_new_n298__ = ~new_new_n234__ & new_new_n240__;
  assign new_new_n299__ = new_new_n271__ & new_new_n298__;
  assign new_new_n300__ = new_new_n283__ & new_new_n299__;
  assign new_new_n301__ = ~G122 & ~new_new_n300__;
  assign new_new_n302__ = G122 & new_new_n300__;
  assign G24 = ~new_new_n301__ & ~new_new_n302__;
  assign new_new_n304__ = new_new_n254__ & new_new_n277__;
  assign new_new_n305__ = new_new_n283__ & new_new_n304__;
  assign new_new_n306__ = ~G125 & ~new_new_n305__;
  assign new_new_n307__ = G125 & new_new_n305__;
  assign G27 = ~new_new_n306__ & ~new_new_n307__;
  assign new_new_n309__ = ~new_new_n126__ & new_new_n156__;
  assign new_new_n310__ = new_new_n176__ & new_new_n309__;
  assign new_new_n311__ = new_new_n124__ & new_new_n310__;
  assign new_new_n312__ = new_new_n277__ & new_new_n311__;
  assign new_new_n313__ = ~G131 & ~new_new_n312__;
  assign new_new_n314__ = G131 & new_new_n312__;
  assign G33 = ~new_new_n313__ & ~new_new_n314__;
  assign new_new_n316__ = new_new_n266__ & new_new_n311__;
  assign new_new_n317__ = ~G134 & ~new_new_n316__;
  assign new_new_n318__ = G134 & new_new_n316__;
  assign G36 = ~new_new_n317__ & ~new_new_n318__;
  assign new_new_n320__ = new_new_n227__ & ~new_new_n265__;
  assign new_new_n321__ = new_new_n261__ & new_new_n320__;
  assign new_new_n322__ = new_new_n310__ & new_new_n321__;
  assign new_new_n323__ = ~G137 & ~new_new_n322__;
  assign new_new_n324__ = G137 & new_new_n322__;
  assign G39 = ~new_new_n323__ & ~new_new_n324__;
  assign new_new_n326__ = new_new_n304__ & new_new_n310__;
  assign new_new_n327__ = ~G140 & ~new_new_n326__;
  assign new_new_n328__ = G140 & new_new_n326__;
  assign G42 = ~new_new_n327__ & ~new_new_n328__;
  assign new_new_n330__ = ~new_new_n236__ & ~new_new_n244__;
  assign new_new_n331__ = ~new_new_n250__ & ~new_new_n257__;
  assign new_new_n332__ = ~new_new_n285__ & ~new_new_n289__;
  assign new_new_n333__ = ~new_new_n294__ & ~new_new_n300__;
  assign new_new_n334__ = new_new_n332__ & new_new_n333__;
  assign new_new_n335__ = new_new_n330__ & new_new_n331__;
  assign new_new_n336__ = new_new_n334__ & new_new_n335__;
  assign new_new_n337__ = ~new_new_n267__ & ~new_new_n273__;
  assign new_new_n338__ = ~new_new_n278__ & ~new_new_n305__;
  assign new_new_n339__ = ~new_new_n312__ & ~new_new_n316__;
  assign new_new_n340__ = ~new_new_n322__ & ~new_new_n326__;
  assign new_new_n341__ = new_new_n339__ & new_new_n340__;
  assign new_new_n342__ = new_new_n337__ & new_new_n338__;
  assign new_new_n343__ = new_new_n341__ & new_new_n342__;
  assign new_new_n344__ = new_new_n336__ & new_new_n343__;
  assign new_new_n345__ = new_new_n282__ & new_new_n309__;
  assign new_new_n346__ = ~new_new_n227__ & new_new_n240__;
  assign new_new_n347__ = ~new_new_n271__ & new_new_n346__;
  assign new_new_n348__ = ~new_new_n255__ & ~new_new_n347__;
  assign new_new_n349__ = new_new_n345__ & ~new_new_n348__;
  assign new_new_n350__ = new_new_n227__ & new_new_n240__;
  assign new_new_n351__ = new_new_n126__ & new_new_n158__;
  assign new_new_n352__ = ~new_new_n126__ & ~new_new_n158__;
  assign new_new_n353__ = ~new_new_n351__ & ~new_new_n352__;
  assign new_new_n354__ = new_new_n156__ & new_new_n353__;
  assign new_new_n355__ = new_new_n175__ & new_new_n354__;
  assign new_new_n356__ = new_new_n350__ & new_new_n355__;
  assign new_new_n357__ = ~new_new_n349__ & ~new_new_n356__;
  assign new_new_n358__ = ~new_new_n229__ & ~new_new_n357__;
  assign new_new_n359__ = new_new_n124__ & new_new_n345__;
  assign new_new_n360__ = ~new_new_n283__ & ~new_new_n310__;
  assign new_new_n361__ = new_new_n240__ & ~new_new_n360__;
  assign new_new_n362__ = ~new_new_n359__ & ~new_new_n361__;
  assign new_new_n363__ = new_new_n227__ & new_new_n233__;
  assign new_new_n364__ = ~new_new_n362__ & new_new_n363__;
  assign new_new_n365__ = ~new_new_n358__ & ~new_new_n364__;
  assign new_new_n366__ = new_new_n344__ & new_new_n365__;
  assign new_new_n367__ = G952 & ~new_new_n366__;
  assign new_new_n368__ = new_new_n345__ & new_new_n350__;
  assign new_new_n369__ = ~G953 & ~new_new_n368__;
  assign G75 = new_new_n367__ | ~new_new_n369__;
  assign new_new_n371__ = ~G952 & G953;
  assign new_new_n372__ = G210 & G902;
  assign new_new_n373__ = ~new_new_n344__ & new_new_n372__;
  assign new_new_n374__ = new_new_n152__ & new_new_n373__;
  assign new_new_n375__ = ~new_new_n152__ & ~new_new_n373__;
  assign new_new_n376__ = ~new_new_n371__ & ~new_new_n374__;
  assign G51 = ~new_new_n375__ & new_new_n376__;
  assign new_new_n378__ = G469 & G902;
  assign new_new_n379__ = ~new_new_n344__ & new_new_n378__;
  assign new_new_n380__ = ~new_new_n171__ & new_new_n379__;
  assign new_new_n381__ = new_new_n171__ & ~new_new_n379__;
  assign new_new_n382__ = ~new_new_n371__ & ~new_new_n380__;
  assign G54 = ~new_new_n381__ & new_new_n382__;
  assign new_new_n384__ = G475 & G902;
  assign new_new_n385__ = ~new_new_n344__ & new_new_n384__;
  assign new_new_n386__ = new_new_n222__ & ~new_new_n385__;
  assign new_new_n387__ = ~new_new_n222__ & new_new_n385__;
  assign new_new_n388__ = ~new_new_n371__ & ~new_new_n386__;
  assign G60 = ~new_new_n387__ & new_new_n388__;
  assign new_new_n390__ = G478 & G902;
  assign new_new_n391__ = ~new_new_n344__ & new_new_n390__;
  assign new_new_n392__ = new_new_n198__ & ~new_new_n391__;
  assign new_new_n393__ = ~new_new_n198__ & new_new_n391__;
  assign new_new_n394__ = ~new_new_n371__ & ~new_new_n392__;
  assign G63 = ~new_new_n393__ & new_new_n394__;
  assign new_new_n396__ = G217 & G902;
  assign new_new_n397__ = ~new_new_n344__ & new_new_n396__;
  assign new_new_n398__ = ~new_new_n81__ & new_new_n397__;
  assign new_new_n399__ = new_new_n81__ & ~new_new_n397__;
  assign new_new_n400__ = ~new_new_n371__ & ~new_new_n398__;
  assign G66 = ~new_new_n399__ & new_new_n400__;
  assign new_new_n402__ = ~G953 & ~new_new_n336__;
  assign new_new_n403__ = ~G224 & G953;
  assign new_new_n404__ = ~new_new_n402__ & ~new_new_n403__;
  assign new_new_n405__ = ~new_new_n142__ & ~new_new_n404__;
  assign new_new_n406__ = new_new_n142__ & new_new_n404__;
  assign new_new_n407__ = ~new_new_n405__ & ~new_new_n406__;
  assign G69 = new_new_n228__ | new_new_n407__;
  assign new_new_n409__ = ~G953 & ~new_new_n343__;
  assign new_new_n410__ = ~G227 & G953;
  assign new_new_n411__ = ~new_new_n263__ & ~new_new_n410__;
  assign new_new_n412__ = ~new_new_n409__ & new_new_n411__;
  assign new_new_n413__ = new_new_n61__ & ~new_new_n102__;
  assign new_new_n414__ = ~new_new_n61__ & new_new_n102__;
  assign new_new_n415__ = ~new_new_n413__ & ~new_new_n414__;
  assign new_new_n416__ = ~new_new_n263__ & ~new_new_n415__;
  assign new_new_n417__ = ~new_new_n412__ & new_new_n416__;
  assign new_new_n418__ = new_new_n412__ & ~new_new_n416__;
  assign G72 = ~new_new_n417__ & ~new_new_n418__;
  assign new_new_n420__ = G472 & G902;
  assign new_new_n421__ = ~new_new_n344__ & new_new_n420__;
  assign new_new_n422__ = ~new_new_n119__ & new_new_n421__;
  assign new_new_n423__ = new_new_n119__ & ~new_new_n421__;
  assign new_new_n424__ = ~new_new_n371__ & ~new_new_n422__;
  assign G57 = ~new_new_n423__ & new_new_n424__;
endmodule


