module max_2(pi0 , po0 );
  input pi0 ;
  output po0 ;
  assign po0 = pi0 ;
endmodule
