module adder32_2(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , po0 , po1 , po2 , po3 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 ;
  output po0 , po1 , po2 , po3 ;
  wire new_n7, new_n8, new_n9, new_n10, new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23;
  assign new_n7 = pi0 & pi3 ;
  assign new_n8 = ~pi0 & ~pi3 ;
  assign new_n9 = ~new_n7 & ~new_n8 ;
  assign new_n10 = pi1 & pi4 ;
  assign new_n11 = ~pi1 & ~pi4 ;
  assign new_n12 = ~new_n10 & ~new_n11 ;
  assign new_n13 = new_n7 & new_n12 ;
  assign new_n14 = ~new_n7 & ~new_n12 ;
  assign new_n15 = ~new_n13 & ~new_n14 ;
  assign new_n16 = ~new_n10 & ~new_n13 ;
  assign new_n17 = pi2 & pi5 ;
  assign new_n18 = ~pi2 & ~pi5 ;
  assign new_n19 = ~new_n17 & ~new_n18 ;
  assign new_n20 = ~new_n16 & new_n19 ;
  assign new_n21 = new_n16 & ~new_n19 ;
  assign new_n22 = ~new_n20 & ~new_n21 ;
  assign new_n23 = ~new_n17 & ~new_n20 ;
  assign po0 = new_n9 ;
  assign po1 = new_n15 ;
  assign po2 = new_n22 ;
  assign po3 = new_n23 ;
endmodule
