// Benchmark "c3540" written by ABC on Thu Jul 14 21:14:18 2022

module c3540 ( 
    G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
    G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200,
    G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274,
    G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698,
    G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107,
    G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
    G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270,
    G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_new_n73__, new_new_n74__, new_new_n76__, new_new_n78__,
    new_new_n79__, new_new_n80__, new_new_n81__, new_new_n82__,
    new_new_n83__, new_new_n84__, new_new_n85__, new_new_n86__,
    new_new_n87__, new_new_n88__, new_new_n89__, new_new_n90__,
    new_new_n91__, new_new_n92__, new_new_n93__, new_new_n94__,
    new_new_n95__, new_new_n96__, new_new_n97__, new_new_n98__,
    new_new_n99__, new_new_n100__, new_new_n101__, new_new_n102__,
    new_new_n103__, new_new_n104__, new_new_n106__, new_new_n107__,
    new_new_n108__, new_new_n109__, new_new_n110__, new_new_n111__,
    new_new_n112__, new_new_n113__, new_new_n114__, new_new_n115__,
    new_new_n116__, new_new_n117__, new_new_n118__, new_new_n119__,
    new_new_n120__, new_new_n121__, new_new_n122__, new_new_n123__,
    new_new_n124__, new_new_n125__, new_new_n127__, new_new_n128__,
    new_new_n129__, new_new_n130__, new_new_n131__, new_new_n132__,
    new_new_n133__, new_new_n134__, new_new_n135__, new_new_n136__,
    new_new_n137__, new_new_n138__, new_new_n139__, new_new_n140__,
    new_new_n141__, new_new_n142__, new_new_n143__, new_new_n144__,
    new_new_n145__, new_new_n147__, new_new_n148__, new_new_n149__,
    new_new_n150__, new_new_n151__, new_new_n152__, new_new_n153__,
    new_new_n154__, new_new_n155__, new_new_n156__, new_new_n157__,
    new_new_n158__, new_new_n159__, new_new_n160__, new_new_n161__,
    new_new_n162__, new_new_n163__, new_new_n164__, new_new_n165__,
    new_new_n166__, new_new_n167__, new_new_n168__, new_new_n169__,
    new_new_n170__, new_new_n171__, new_new_n172__, new_new_n173__,
    new_new_n174__, new_new_n175__, new_new_n176__, new_new_n177__,
    new_new_n178__, new_new_n179__, new_new_n180__, new_new_n181__,
    new_new_n182__, new_new_n183__, new_new_n184__, new_new_n185__,
    new_new_n186__, new_new_n187__, new_new_n188__, new_new_n189__,
    new_new_n190__, new_new_n191__, new_new_n192__, new_new_n193__,
    new_new_n194__, new_new_n195__, new_new_n196__, new_new_n197__,
    new_new_n198__, new_new_n199__, new_new_n200__, new_new_n201__,
    new_new_n202__, new_new_n203__, new_new_n204__, new_new_n205__,
    new_new_n206__, new_new_n207__, new_new_n208__, new_new_n209__,
    new_new_n210__, new_new_n211__, new_new_n212__, new_new_n213__,
    new_new_n214__, new_new_n215__, new_new_n216__, new_new_n217__,
    new_new_n218__, new_new_n219__, new_new_n220__, new_new_n221__,
    new_new_n222__, new_new_n223__, new_new_n224__, new_new_n225__,
    new_new_n226__, new_new_n227__, new_new_n228__, new_new_n229__,
    new_new_n230__, new_new_n231__, new_new_n232__, new_new_n233__,
    new_new_n234__, new_new_n235__, new_new_n236__, new_new_n237__,
    new_new_n238__, new_new_n239__, new_new_n240__, new_new_n241__,
    new_new_n242__, new_new_n243__, new_new_n244__, new_new_n245__,
    new_new_n246__, new_new_n247__, new_new_n248__, new_new_n249__,
    new_new_n250__, new_new_n251__, new_new_n252__, new_new_n253__,
    new_new_n254__, new_new_n255__, new_new_n256__, new_new_n257__,
    new_new_n258__, new_new_n259__, new_new_n260__, new_new_n261__,
    new_new_n262__, new_new_n263__, new_new_n264__, new_new_n265__,
    new_new_n266__, new_new_n267__, new_new_n268__, new_new_n269__,
    new_new_n270__, new_new_n271__, new_new_n272__, new_new_n273__,
    new_new_n274__, new_new_n275__, new_new_n276__, new_new_n277__,
    new_new_n278__, new_new_n279__, new_new_n280__, new_new_n281__,
    new_new_n282__, new_new_n283__, new_new_n284__, new_new_n285__,
    new_new_n286__, new_new_n287__, new_new_n288__, new_new_n289__,
    new_new_n290__, new_new_n291__, new_new_n292__, new_new_n293__,
    new_new_n294__, new_new_n295__, new_new_n296__, new_new_n297__,
    new_new_n298__, new_new_n299__, new_new_n300__, new_new_n301__,
    new_new_n302__, new_new_n303__, new_new_n304__, new_new_n305__,
    new_new_n306__, new_new_n307__, new_new_n308__, new_new_n309__,
    new_new_n310__, new_new_n311__, new_new_n312__, new_new_n313__,
    new_new_n314__, new_new_n315__, new_new_n316__, new_new_n317__,
    new_new_n318__, new_new_n319__, new_new_n320__, new_new_n321__,
    new_new_n322__, new_new_n323__, new_new_n324__, new_new_n325__,
    new_new_n326__, new_new_n327__, new_new_n328__, new_new_n329__,
    new_new_n330__, new_new_n331__, new_new_n332__, new_new_n333__,
    new_new_n334__, new_new_n335__, new_new_n336__, new_new_n337__,
    new_new_n338__, new_new_n339__, new_new_n340__, new_new_n341__,
    new_new_n342__, new_new_n343__, new_new_n344__, new_new_n345__,
    new_new_n346__, new_new_n347__, new_new_n348__, new_new_n349__,
    new_new_n350__, new_new_n351__, new_new_n352__, new_new_n353__,
    new_new_n354__, new_new_n355__, new_new_n356__, new_new_n357__,
    new_new_n358__, new_new_n359__, new_new_n360__, new_new_n361__,
    new_new_n362__, new_new_n363__, new_new_n364__, new_new_n365__,
    new_new_n366__, new_new_n367__, new_new_n368__, new_new_n369__,
    new_new_n370__, new_new_n371__, new_new_n372__, new_new_n373__,
    new_new_n374__, new_new_n375__, new_new_n376__, new_new_n377__,
    new_new_n378__, new_new_n379__, new_new_n380__, new_new_n381__,
    new_new_n382__, new_new_n383__, new_new_n384__, new_new_n385__,
    new_new_n386__, new_new_n387__, new_new_n388__, new_new_n389__,
    new_new_n390__, new_new_n391__, new_new_n392__, new_new_n393__,
    new_new_n394__, new_new_n395__, new_new_n396__, new_new_n397__,
    new_new_n398__, new_new_n399__, new_new_n400__, new_new_n401__,
    new_new_n402__, new_new_n403__, new_new_n404__, new_new_n405__,
    new_new_n406__, new_new_n407__, new_new_n408__, new_new_n409__,
    new_new_n410__, new_new_n412__, new_new_n413__, new_new_n414__,
    new_new_n415__, new_new_n416__, new_new_n417__, new_new_n418__,
    new_new_n419__, new_new_n420__, new_new_n421__, new_new_n422__,
    new_new_n423__, new_new_n424__, new_new_n426__, new_new_n427__,
    new_new_n428__, new_new_n429__, new_new_n430__, new_new_n431__,
    new_new_n432__, new_new_n433__, new_new_n434__, new_new_n435__,
    new_new_n436__, new_new_n437__, new_new_n438__, new_new_n439__,
    new_new_n440__, new_new_n441__, new_new_n442__, new_new_n444__,
    new_new_n445__, new_new_n446__, new_new_n447__, new_new_n448__,
    new_new_n449__, new_new_n450__, new_new_n451__, new_new_n452__,
    new_new_n453__, new_new_n454__, new_new_n455__, new_new_n456__,
    new_new_n457__, new_new_n458__, new_new_n459__, new_new_n460__,
    new_new_n461__, new_new_n462__, new_new_n463__, new_new_n464__,
    new_new_n466__, new_new_n467__, new_new_n468__, new_new_n469__,
    new_new_n470__, new_new_n471__, new_new_n472__, new_new_n473__,
    new_new_n474__, new_new_n475__, new_new_n476__, new_new_n477__,
    new_new_n478__, new_new_n479__, new_new_n480__, new_new_n481__,
    new_new_n482__, new_new_n483__, new_new_n484__, new_new_n485__,
    new_new_n486__, new_new_n487__, new_new_n488__, new_new_n489__,
    new_new_n490__, new_new_n491__, new_new_n492__, new_new_n493__,
    new_new_n494__, new_new_n495__, new_new_n496__, new_new_n497__,
    new_new_n498__, new_new_n499__, new_new_n500__, new_new_n501__,
    new_new_n502__, new_new_n503__, new_new_n504__, new_new_n505__,
    new_new_n506__, new_new_n507__, new_new_n508__, new_new_n509__,
    new_new_n510__, new_new_n511__, new_new_n512__, new_new_n513__,
    new_new_n514__, new_new_n515__, new_new_n516__, new_new_n517__,
    new_new_n518__, new_new_n519__, new_new_n520__, new_new_n521__,
    new_new_n522__, new_new_n523__, new_new_n524__, new_new_n525__,
    new_new_n526__, new_new_n527__, new_new_n528__, new_new_n529__,
    new_new_n530__, new_new_n531__, new_new_n532__, new_new_n533__,
    new_new_n534__, new_new_n535__, new_new_n536__, new_new_n537__,
    new_new_n538__, new_new_n539__, new_new_n540__, new_new_n541__,
    new_new_n543__, new_new_n544__, new_new_n545__, new_new_n546__,
    new_new_n547__, new_new_n548__, new_new_n549__, new_new_n550__,
    new_new_n551__, new_new_n552__, new_new_n553__, new_new_n554__,
    new_new_n555__, new_new_n556__, new_new_n557__, new_new_n558__,
    new_new_n559__, new_new_n560__, new_new_n561__, new_new_n562__,
    new_new_n563__, new_new_n564__, new_new_n565__, new_new_n566__,
    new_new_n567__, new_new_n568__, new_new_n569__, new_new_n570__,
    new_new_n571__, new_new_n572__, new_new_n573__, new_new_n574__,
    new_new_n575__, new_new_n576__, new_new_n577__, new_new_n578__,
    new_new_n579__, new_new_n580__, new_new_n581__, new_new_n582__,
    new_new_n583__, new_new_n584__, new_new_n585__, new_new_n586__,
    new_new_n587__, new_new_n588__, new_new_n589__, new_new_n590__,
    new_new_n591__, new_new_n592__, new_new_n593__, new_new_n595__,
    new_new_n596__, new_new_n597__, new_new_n598__, new_new_n599__,
    new_new_n600__, new_new_n601__, new_new_n602__, new_new_n603__,
    new_new_n604__, new_new_n605__, new_new_n606__, new_new_n607__,
    new_new_n608__, new_new_n609__, new_new_n610__, new_new_n611__,
    new_new_n612__, new_new_n613__, new_new_n614__, new_new_n615__,
    new_new_n616__, new_new_n617__, new_new_n618__, new_new_n619__,
    new_new_n620__, new_new_n621__, new_new_n622__, new_new_n623__,
    new_new_n624__, new_new_n625__, new_new_n626__, new_new_n627__,
    new_new_n628__, new_new_n629__, new_new_n630__, new_new_n631__,
    new_new_n632__, new_new_n633__, new_new_n635__, new_new_n636__,
    new_new_n637__, new_new_n638__, new_new_n639__, new_new_n640__,
    new_new_n641__, new_new_n642__, new_new_n643__, new_new_n644__,
    new_new_n645__, new_new_n646__, new_new_n647__, new_new_n648__,
    new_new_n649__, new_new_n650__, new_new_n651__, new_new_n652__,
    new_new_n653__, new_new_n654__, new_new_n655__, new_new_n656__,
    new_new_n657__, new_new_n658__, new_new_n659__, new_new_n660__,
    new_new_n661__, new_new_n662__, new_new_n663__, new_new_n664__,
    new_new_n665__, new_new_n666__, new_new_n667__, new_new_n668__,
    new_new_n669__, new_new_n670__, new_new_n671__, new_new_n672__,
    new_new_n673__, new_new_n674__, new_new_n675__, new_new_n676__,
    new_new_n677__, new_new_n678__, new_new_n679__, new_new_n680__,
    new_new_n681__, new_new_n682__, new_new_n683__, new_new_n684__,
    new_new_n685__, new_new_n686__, new_new_n687__, new_new_n688__,
    new_new_n689__, new_new_n690__, new_new_n691__, new_new_n692__,
    new_new_n693__, new_new_n694__, new_new_n695__, new_new_n696__,
    new_new_n697__, new_new_n698__, new_new_n699__, new_new_n700__,
    new_new_n701__, new_new_n702__, new_new_n703__, new_new_n704__,
    new_new_n705__, new_new_n706__, new_new_n707__, new_new_n708__,
    new_new_n709__, new_new_n710__, new_new_n712__, new_new_n713__,
    new_new_n714__, new_new_n715__, new_new_n716__, new_new_n717__,
    new_new_n718__, new_new_n719__, new_new_n720__, new_new_n721__,
    new_new_n722__, new_new_n723__, new_new_n724__, new_new_n725__,
    new_new_n726__, new_new_n727__, new_new_n728__, new_new_n729__,
    new_new_n730__, new_new_n731__, new_new_n732__, new_new_n733__,
    new_new_n734__, new_new_n735__, new_new_n736__, new_new_n737__,
    new_new_n738__, new_new_n739__, new_new_n740__, new_new_n741__,
    new_new_n742__, new_new_n743__, new_new_n744__, new_new_n745__,
    new_new_n746__, new_new_n747__, new_new_n748__, new_new_n749__,
    new_new_n750__, new_new_n751__, new_new_n752__, new_new_n753__,
    new_new_n754__, new_new_n755__, new_new_n756__, new_new_n757__,
    new_new_n758__, new_new_n759__, new_new_n760__, new_new_n761__,
    new_new_n762__, new_new_n763__, new_new_n764__, new_new_n765__,
    new_new_n766__, new_new_n768__, new_new_n769__, new_new_n770__,
    new_new_n771__, new_new_n772__, new_new_n773__, new_new_n774__,
    new_new_n775__, new_new_n776__, new_new_n777__, new_new_n778__,
    new_new_n779__, new_new_n780__, new_new_n781__, new_new_n782__,
    new_new_n783__, new_new_n784__, new_new_n785__, new_new_n786__,
    new_new_n787__, new_new_n788__, new_new_n789__, new_new_n790__,
    new_new_n791__, new_new_n792__, new_new_n793__, new_new_n794__,
    new_new_n795__, new_new_n796__, new_new_n797__, new_new_n798__,
    new_new_n799__, new_new_n800__, new_new_n801__, new_new_n802__,
    new_new_n803__, new_new_n804__, new_new_n805__, new_new_n806__,
    new_new_n807__, new_new_n808__, new_new_n809__, new_new_n810__,
    new_new_n811__, new_new_n812__, new_new_n814__, new_new_n815__,
    new_new_n816__, new_new_n817__, new_new_n818__, new_new_n819__,
    new_new_n820__, new_new_n821__, new_new_n822__, new_new_n823__,
    new_new_n824__, new_new_n825__, new_new_n826__, new_new_n827__,
    new_new_n828__, new_new_n829__, new_new_n830__, new_new_n831__,
    new_new_n832__, new_new_n833__, new_new_n834__, new_new_n835__,
    new_new_n836__, new_new_n837__, new_new_n838__, new_new_n839__,
    new_new_n840__, new_new_n841__, new_new_n842__, new_new_n843__,
    new_new_n844__, new_new_n845__, new_new_n846__, new_new_n847__,
    new_new_n848__, new_new_n849__, new_new_n850__, new_new_n851__,
    new_new_n852__, new_new_n853__, new_new_n854__, new_new_n855__,
    new_new_n856__, new_new_n857__, new_new_n858__, new_new_n859__,
    new_new_n860__, new_new_n861__, new_new_n862__, new_new_n863__,
    new_new_n864__, new_new_n865__, new_new_n866__, new_new_n867__,
    new_new_n868__, new_new_n869__, new_new_n870__, new_new_n871__,
    new_new_n872__, new_new_n873__, new_new_n875__, new_new_n876__,
    new_new_n877__, new_new_n878__, new_new_n879__, new_new_n880__,
    new_new_n881__, new_new_n882__, new_new_n883__, new_new_n884__,
    new_new_n885__, new_new_n886__, new_new_n887__, new_new_n888__,
    new_new_n889__, new_new_n890__, new_new_n891__, new_new_n892__,
    new_new_n893__, new_new_n894__, new_new_n895__, new_new_n896__,
    new_new_n897__, new_new_n898__, new_new_n899__, new_new_n900__,
    new_new_n901__, new_new_n902__, new_new_n903__, new_new_n904__,
    new_new_n905__, new_new_n906__, new_new_n907__, new_new_n908__,
    new_new_n909__, new_new_n910__, new_new_n911__, new_new_n912__,
    new_new_n913__, new_new_n914__, new_new_n915__, new_new_n916__,
    new_new_n917__, new_new_n918__, new_new_n919__, new_new_n920__,
    new_new_n921__, new_new_n922__, new_new_n923__, new_new_n924__,
    new_new_n925__, new_new_n926__, new_new_n927__, new_new_n928__,
    new_new_n929__, new_new_n930__, new_new_n931__, new_new_n933__,
    new_new_n934__, new_new_n935__, new_new_n936__, new_new_n937__,
    new_new_n938__, new_new_n939__, new_new_n940__, new_new_n941__,
    new_new_n942__, new_new_n943__, new_new_n944__, new_new_n945__,
    new_new_n946__, new_new_n947__, new_new_n948__, new_new_n949__,
    new_new_n950__, new_new_n951__, new_new_n952__, new_new_n953__,
    new_new_n954__, new_new_n955__, new_new_n956__, new_new_n957__,
    new_new_n958__, new_new_n959__, new_new_n960__, new_new_n961__,
    new_new_n962__, new_new_n963__, new_new_n964__, new_new_n965__,
    new_new_n966__, new_new_n967__, new_new_n968__, new_new_n969__,
    new_new_n970__, new_new_n971__, new_new_n972__, new_new_n973__,
    new_new_n975__, new_new_n976__, new_new_n977__, new_new_n978__,
    new_new_n979__, new_new_n980__, new_new_n982__, new_new_n983__,
    new_new_n984__, new_new_n986__, new_new_n987__, new_new_n988__,
    new_new_n989__, new_new_n990__, new_new_n991__, new_new_n992__,
    new_new_n993__, new_new_n994__, new_new_n995__, new_new_n996__,
    new_new_n997__, new_new_n998__, new_new_n999__, new_new_n1000__,
    new_new_n1001__, new_new_n1002__, new_new_n1003__, new_new_n1004__,
    new_new_n1005__, new_new_n1007__, new_new_n1008__;
  assign new_new_n73__ = ~G58 & ~G68;
  assign new_new_n74__ = ~G50 & new_new_n73__;
  assign G353 = ~G77 & new_new_n74__;
  assign new_new_n76__ = ~G97 & ~G107;
  assign G355 = ~G87 | new_new_n76__;
  assign new_new_n78__ = G1 & G13;
  assign new_new_n79__ = G20 & new_new_n78__;
  assign new_new_n80__ = G50 & ~new_new_n73__;
  assign new_new_n81__ = new_new_n79__ & new_new_n80__;
  assign new_new_n82__ = G1 & G20;
  assign new_new_n83__ = G58 & G232;
  assign new_new_n84__ = G107 & G264;
  assign new_new_n85__ = G77 & G244;
  assign new_new_n86__ = G68 & G238;
  assign new_new_n87__ = G50 & G226;
  assign new_new_n88__ = G116 & G270;
  assign new_new_n89__ = G87 & G250;
  assign new_new_n90__ = G97 & G257;
  assign new_new_n91__ = ~new_new_n83__ & ~new_new_n84__;
  assign new_new_n92__ = ~new_new_n85__ & ~new_new_n86__;
  assign new_new_n93__ = ~new_new_n87__ & ~new_new_n88__;
  assign new_new_n94__ = ~new_new_n89__ & ~new_new_n90__;
  assign new_new_n95__ = new_new_n93__ & new_new_n94__;
  assign new_new_n96__ = new_new_n91__ & new_new_n92__;
  assign new_new_n97__ = new_new_n95__ & new_new_n96__;
  assign new_new_n98__ = ~new_new_n82__ & ~new_new_n97__;
  assign new_new_n99__ = G1 & ~G13;
  assign new_new_n100__ = G20 & new_new_n99__;
  assign new_new_n101__ = ~G257 & ~G264;
  assign new_new_n102__ = G250 & ~new_new_n101__;
  assign new_new_n103__ = new_new_n100__ & new_new_n102__;
  assign new_new_n104__ = ~new_new_n81__ & ~new_new_n103__;
  assign G361 = ~new_new_n98__ & new_new_n104__;
  assign new_new_n106__ = ~G264 & ~G270;
  assign new_new_n107__ = G264 & G270;
  assign new_new_n108__ = ~new_new_n106__ & ~new_new_n107__;
  assign new_new_n109__ = G250 & ~G257;
  assign new_new_n110__ = ~G250 & G257;
  assign new_new_n111__ = ~new_new_n109__ & ~new_new_n110__;
  assign new_new_n112__ = new_new_n108__ & new_new_n111__;
  assign new_new_n113__ = ~new_new_n108__ & ~new_new_n111__;
  assign new_new_n114__ = ~new_new_n112__ & ~new_new_n113__;
  assign new_new_n115__ = ~G238 & ~G244;
  assign new_new_n116__ = G238 & G244;
  assign new_new_n117__ = ~new_new_n115__ & ~new_new_n116__;
  assign new_new_n118__ = G226 & ~G232;
  assign new_new_n119__ = ~G226 & G232;
  assign new_new_n120__ = ~new_new_n118__ & ~new_new_n119__;
  assign new_new_n121__ = new_new_n117__ & new_new_n120__;
  assign new_new_n122__ = ~new_new_n117__ & ~new_new_n120__;
  assign new_new_n123__ = ~new_new_n121__ & ~new_new_n122__;
  assign new_new_n124__ = new_new_n114__ & new_new_n123__;
  assign new_new_n125__ = ~new_new_n114__ & ~new_new_n123__;
  assign G358 = new_new_n124__ | new_new_n125__;
  assign new_new_n127__ = G58 & G68;
  assign new_new_n128__ = ~new_new_n73__ & ~new_new_n127__;
  assign new_new_n129__ = ~G50 & ~G77;
  assign new_new_n130__ = G50 & G77;
  assign new_new_n131__ = ~new_new_n129__ & ~new_new_n130__;
  assign new_new_n132__ = new_new_n128__ & ~new_new_n131__;
  assign new_new_n133__ = ~new_new_n128__ & new_new_n131__;
  assign new_new_n134__ = ~new_new_n132__ & ~new_new_n133__;
  assign new_new_n135__ = ~G87 & ~G97;
  assign new_new_n136__ = G87 & G97;
  assign new_new_n137__ = ~new_new_n135__ & ~new_new_n136__;
  assign new_new_n138__ = G107 & ~G116;
  assign new_new_n139__ = ~G107 & G116;
  assign new_new_n140__ = ~new_new_n138__ & ~new_new_n139__;
  assign new_new_n141__ = new_new_n137__ & new_new_n140__;
  assign new_new_n142__ = ~new_new_n137__ & ~new_new_n140__;
  assign new_new_n143__ = ~new_new_n141__ & ~new_new_n142__;
  assign new_new_n144__ = new_new_n134__ & new_new_n143__;
  assign new_new_n145__ = ~new_new_n134__ & ~new_new_n143__;
  assign G351 = new_new_n144__ | new_new_n145__;
  assign new_new_n147__ = G33 & G41;
  assign new_new_n148__ = new_new_n78__ & ~new_new_n147__;
  assign new_new_n149__ = G33 & G303;
  assign new_new_n150__ = ~G33 & G1698;
  assign new_new_n151__ = G264 & new_new_n150__;
  assign new_new_n152__ = ~G33 & ~G1698;
  assign new_new_n153__ = G257 & new_new_n152__;
  assign new_new_n154__ = ~new_new_n149__ & ~new_new_n151__;
  assign new_new_n155__ = ~new_new_n153__ & new_new_n154__;
  assign new_new_n156__ = new_new_n148__ & ~new_new_n155__;
  assign new_new_n157__ = G274 & ~new_new_n148__;
  assign new_new_n158__ = ~G1 & G45;
  assign new_new_n159__ = ~G41 & new_new_n158__;
  assign new_new_n160__ = new_new_n157__ & new_new_n159__;
  assign new_new_n161__ = ~new_new_n148__ & ~new_new_n159__;
  assign new_new_n162__ = G270 & new_new_n161__;
  assign new_new_n163__ = ~new_new_n160__ & ~new_new_n162__;
  assign new_new_n164__ = ~new_new_n156__ & new_new_n163__;
  assign new_new_n165__ = G169 & ~new_new_n164__;
  assign new_new_n166__ = G179 & new_new_n164__;
  assign new_new_n167__ = ~new_new_n165__ & ~new_new_n166__;
  assign new_new_n168__ = ~G1 & G13;
  assign new_new_n169__ = G20 & ~G116;
  assign new_new_n170__ = new_new_n168__ & new_new_n169__;
  assign new_new_n171__ = ~G1 & G33;
  assign new_new_n172__ = G33 & new_new_n82__;
  assign new_new_n173__ = ~new_new_n78__ & ~new_new_n172__;
  assign new_new_n174__ = G20 & new_new_n168__;
  assign new_new_n175__ = new_new_n173__ & ~new_new_n174__;
  assign new_new_n176__ = G116 & ~new_new_n171__;
  assign new_new_n177__ = new_new_n175__ & new_new_n176__;
  assign new_new_n178__ = G33 & G283;
  assign new_new_n179__ = ~G33 & G97;
  assign new_new_n180__ = ~G20 & ~new_new_n178__;
  assign new_new_n181__ = ~new_new_n179__ & new_new_n180__;
  assign new_new_n182__ = ~new_new_n169__ & ~new_new_n173__;
  assign new_new_n183__ = ~new_new_n181__ & new_new_n182__;
  assign new_new_n184__ = ~new_new_n170__ & ~new_new_n177__;
  assign new_new_n185__ = ~new_new_n183__ & new_new_n184__;
  assign new_new_n186__ = ~new_new_n167__ & ~new_new_n185__;
  assign new_new_n187__ = G200 & ~new_new_n164__;
  assign new_new_n188__ = G190 & new_new_n164__;
  assign new_new_n189__ = new_new_n185__ & ~new_new_n187__;
  assign new_new_n190__ = ~new_new_n188__ & new_new_n189__;
  assign new_new_n191__ = ~new_new_n186__ & ~new_new_n190__;
  assign new_new_n192__ = ~G87 & new_new_n174__;
  assign new_new_n193__ = G33 & G97;
  assign new_new_n194__ = ~G33 & G68;
  assign new_new_n195__ = ~G20 & ~new_new_n193__;
  assign new_new_n196__ = ~new_new_n194__ & new_new_n195__;
  assign new_new_n197__ = ~G107 & new_new_n135__;
  assign new_new_n198__ = G20 & new_new_n197__;
  assign new_new_n199__ = ~new_new_n173__ & ~new_new_n196__;
  assign new_new_n200__ = ~new_new_n198__ & new_new_n199__;
  assign new_new_n201__ = G87 & ~new_new_n171__;
  assign new_new_n202__ = new_new_n175__ & new_new_n201__;
  assign new_new_n203__ = ~new_new_n192__ & ~new_new_n200__;
  assign new_new_n204__ = ~new_new_n202__ & new_new_n203__;
  assign new_new_n205__ = G33 & G116;
  assign new_new_n206__ = G244 & new_new_n150__;
  assign new_new_n207__ = G238 & new_new_n152__;
  assign new_new_n208__ = ~new_new_n205__ & ~new_new_n206__;
  assign new_new_n209__ = ~new_new_n207__ & new_new_n208__;
  assign new_new_n210__ = new_new_n148__ & ~new_new_n209__;
  assign new_new_n211__ = ~G250 & ~new_new_n158__;
  assign new_new_n212__ = ~G274 & new_new_n158__;
  assign new_new_n213__ = ~new_new_n148__ & ~new_new_n211__;
  assign new_new_n214__ = ~new_new_n212__ & new_new_n213__;
  assign new_new_n215__ = ~new_new_n210__ & ~new_new_n214__;
  assign new_new_n216__ = ~G169 & ~new_new_n215__;
  assign new_new_n217__ = ~G179 & new_new_n215__;
  assign new_new_n218__ = ~new_new_n204__ & ~new_new_n216__;
  assign new_new_n219__ = ~new_new_n217__ & new_new_n218__;
  assign new_new_n220__ = G190 & new_new_n215__;
  assign new_new_n221__ = G200 & ~new_new_n215__;
  assign new_new_n222__ = new_new_n204__ & ~new_new_n220__;
  assign new_new_n223__ = ~new_new_n221__ & new_new_n222__;
  assign new_new_n224__ = ~new_new_n219__ & ~new_new_n223__;
  assign new_new_n225__ = ~G97 & new_new_n174__;
  assign new_new_n226__ = G33 & G107;
  assign new_new_n227__ = ~G33 & G77;
  assign new_new_n228__ = ~G20 & ~new_new_n226__;
  assign new_new_n229__ = ~new_new_n227__ & new_new_n228__;
  assign new_new_n230__ = G97 & G107;
  assign new_new_n231__ = G20 & ~new_new_n76__;
  assign new_new_n232__ = ~new_new_n230__ & new_new_n231__;
  assign new_new_n233__ = ~new_new_n173__ & ~new_new_n229__;
  assign new_new_n234__ = ~new_new_n232__ & new_new_n233__;
  assign new_new_n235__ = G97 & ~new_new_n171__;
  assign new_new_n236__ = new_new_n175__ & new_new_n235__;
  assign new_new_n237__ = ~new_new_n225__ & ~new_new_n234__;
  assign new_new_n238__ = ~new_new_n236__ & new_new_n237__;
  assign new_new_n239__ = G257 & new_new_n161__;
  assign new_new_n240__ = G244 & new_new_n152__;
  assign new_new_n241__ = G250 & new_new_n150__;
  assign new_new_n242__ = ~new_new_n178__ & ~new_new_n240__;
  assign new_new_n243__ = ~new_new_n241__ & new_new_n242__;
  assign new_new_n244__ = new_new_n148__ & ~new_new_n243__;
  assign new_new_n245__ = ~new_new_n160__ & ~new_new_n239__;
  assign new_new_n246__ = ~new_new_n244__ & new_new_n245__;
  assign new_new_n247__ = ~G169 & ~new_new_n246__;
  assign new_new_n248__ = ~G179 & new_new_n246__;
  assign new_new_n249__ = ~new_new_n238__ & ~new_new_n247__;
  assign new_new_n250__ = ~new_new_n248__ & new_new_n249__;
  assign new_new_n251__ = G200 & ~new_new_n246__;
  assign new_new_n252__ = G190 & new_new_n246__;
  assign new_new_n253__ = new_new_n238__ & ~new_new_n251__;
  assign new_new_n254__ = ~new_new_n252__ & new_new_n253__;
  assign new_new_n255__ = ~new_new_n250__ & ~new_new_n254__;
  assign new_new_n256__ = new_new_n224__ & new_new_n255__;
  assign new_new_n257__ = ~G13 & ~new_new_n172__;
  assign new_new_n258__ = G20 & ~G107;
  assign new_new_n259__ = ~new_new_n257__ & new_new_n258__;
  assign new_new_n260__ = ~G33 & G87;
  assign new_new_n261__ = ~new_new_n205__ & ~new_new_n260__;
  assign new_new_n262__ = ~G20 & ~new_new_n261__;
  assign new_new_n263__ = ~new_new_n173__ & new_new_n262__;
  assign new_new_n264__ = G107 & ~new_new_n171__;
  assign new_new_n265__ = new_new_n175__ & new_new_n264__;
  assign new_new_n266__ = ~new_new_n259__ & ~new_new_n263__;
  assign new_new_n267__ = ~new_new_n265__ & new_new_n266__;
  assign new_new_n268__ = G250 & new_new_n152__;
  assign new_new_n269__ = G257 & new_new_n150__;
  assign new_new_n270__ = G33 & G294;
  assign new_new_n271__ = ~new_new_n268__ & ~new_new_n270__;
  assign new_new_n272__ = ~new_new_n269__ & new_new_n271__;
  assign new_new_n273__ = new_new_n148__ & ~new_new_n272__;
  assign new_new_n274__ = G264 & new_new_n161__;
  assign new_new_n275__ = ~new_new_n160__ & ~new_new_n274__;
  assign new_new_n276__ = ~new_new_n273__ & new_new_n275__;
  assign new_new_n277__ = ~G169 & ~new_new_n276__;
  assign new_new_n278__ = ~G179 & new_new_n276__;
  assign new_new_n279__ = ~new_new_n267__ & ~new_new_n277__;
  assign new_new_n280__ = ~new_new_n278__ & new_new_n279__;
  assign new_new_n281__ = G190 & new_new_n276__;
  assign new_new_n282__ = G200 & ~new_new_n276__;
  assign new_new_n283__ = new_new_n267__ & ~new_new_n281__;
  assign new_new_n284__ = ~new_new_n282__ & new_new_n283__;
  assign new_new_n285__ = ~new_new_n280__ & ~new_new_n284__;
  assign new_new_n286__ = new_new_n191__ & new_new_n285__;
  assign new_new_n287__ = new_new_n256__ & new_new_n286__;
  assign new_new_n288__ = G20 & ~G77;
  assign new_new_n289__ = new_new_n168__ & new_new_n288__;
  assign new_new_n290__ = ~G1 & G20;
  assign new_new_n291__ = G77 & ~new_new_n290__;
  assign new_new_n292__ = new_new_n175__ & new_new_n291__;
  assign new_new_n293__ = G33 & G87;
  assign new_new_n294__ = ~G33 & G58;
  assign new_new_n295__ = ~G20 & ~new_new_n293__;
  assign new_new_n296__ = ~new_new_n294__ & new_new_n295__;
  assign new_new_n297__ = ~new_new_n173__ & ~new_new_n288__;
  assign new_new_n298__ = ~new_new_n296__ & new_new_n297__;
  assign new_new_n299__ = ~new_new_n289__ & ~new_new_n292__;
  assign new_new_n300__ = ~new_new_n298__ & new_new_n299__;
  assign new_new_n301__ = ~G41 & ~G45;
  assign new_new_n302__ = ~G1 & ~new_new_n301__;
  assign new_new_n303__ = ~new_new_n148__ & ~new_new_n302__;
  assign new_new_n304__ = G244 & new_new_n303__;
  assign new_new_n305__ = new_new_n157__ & new_new_n302__;
  assign new_new_n306__ = G238 & new_new_n150__;
  assign new_new_n307__ = G232 & new_new_n152__;
  assign new_new_n308__ = ~new_new_n226__ & ~new_new_n306__;
  assign new_new_n309__ = ~new_new_n307__ & new_new_n308__;
  assign new_new_n310__ = new_new_n148__ & ~new_new_n309__;
  assign new_new_n311__ = ~new_new_n304__ & ~new_new_n305__;
  assign new_new_n312__ = ~new_new_n310__ & new_new_n311__;
  assign new_new_n313__ = ~G169 & ~new_new_n312__;
  assign new_new_n314__ = ~G179 & new_new_n312__;
  assign new_new_n315__ = ~new_new_n300__ & ~new_new_n313__;
  assign new_new_n316__ = ~new_new_n314__ & new_new_n315__;
  assign new_new_n317__ = G200 & ~new_new_n312__;
  assign new_new_n318__ = G190 & new_new_n312__;
  assign new_new_n319__ = new_new_n300__ & ~new_new_n317__;
  assign new_new_n320__ = ~new_new_n318__ & new_new_n319__;
  assign new_new_n321__ = ~new_new_n316__ & ~new_new_n320__;
  assign new_new_n322__ = ~G50 & new_new_n174__;
  assign new_new_n323__ = ~G20 & ~G33;
  assign new_new_n324__ = G150 & new_new_n323__;
  assign new_new_n325__ = G20 & ~new_new_n74__;
  assign new_new_n326__ = ~G20 & G33;
  assign new_new_n327__ = G58 & new_new_n326__;
  assign new_new_n328__ = ~new_new_n324__ & ~new_new_n327__;
  assign new_new_n329__ = ~new_new_n325__ & new_new_n328__;
  assign new_new_n330__ = ~new_new_n173__ & ~new_new_n329__;
  assign new_new_n331__ = G50 & ~new_new_n290__;
  assign new_new_n332__ = new_new_n175__ & new_new_n331__;
  assign new_new_n333__ = ~new_new_n322__ & ~new_new_n330__;
  assign new_new_n334__ = ~new_new_n332__ & new_new_n333__;
  assign new_new_n335__ = G226 & new_new_n303__;
  assign new_new_n336__ = G33 & G77;
  assign new_new_n337__ = G223 & new_new_n150__;
  assign new_new_n338__ = G222 & new_new_n152__;
  assign new_new_n339__ = ~new_new_n336__ & ~new_new_n337__;
  assign new_new_n340__ = ~new_new_n338__ & new_new_n339__;
  assign new_new_n341__ = new_new_n148__ & ~new_new_n340__;
  assign new_new_n342__ = ~new_new_n305__ & ~new_new_n335__;
  assign new_new_n343__ = ~new_new_n341__ & new_new_n342__;
  assign new_new_n344__ = ~G169 & ~new_new_n343__;
  assign new_new_n345__ = ~G179 & new_new_n343__;
  assign new_new_n346__ = ~new_new_n334__ & ~new_new_n344__;
  assign new_new_n347__ = ~new_new_n345__ & new_new_n346__;
  assign new_new_n348__ = G190 & new_new_n343__;
  assign new_new_n349__ = G200 & ~new_new_n343__;
  assign new_new_n350__ = new_new_n334__ & ~new_new_n348__;
  assign new_new_n351__ = ~new_new_n349__ & new_new_n350__;
  assign new_new_n352__ = ~new_new_n347__ & ~new_new_n351__;
  assign new_new_n353__ = ~G58 & new_new_n174__;
  assign new_new_n354__ = G159 & new_new_n323__;
  assign new_new_n355__ = G20 & ~new_new_n128__;
  assign new_new_n356__ = G68 & new_new_n326__;
  assign new_new_n357__ = ~new_new_n354__ & ~new_new_n356__;
  assign new_new_n358__ = ~new_new_n355__ & new_new_n357__;
  assign new_new_n359__ = ~new_new_n173__ & ~new_new_n358__;
  assign new_new_n360__ = G58 & ~new_new_n290__;
  assign new_new_n361__ = new_new_n175__ & new_new_n360__;
  assign new_new_n362__ = ~new_new_n353__ & ~new_new_n359__;
  assign new_new_n363__ = ~new_new_n361__ & new_new_n362__;
  assign new_new_n364__ = G232 & new_new_n303__;
  assign new_new_n365__ = G223 & new_new_n152__;
  assign new_new_n366__ = G226 & new_new_n150__;
  assign new_new_n367__ = ~new_new_n293__ & ~new_new_n365__;
  assign new_new_n368__ = ~new_new_n366__ & new_new_n367__;
  assign new_new_n369__ = new_new_n148__ & ~new_new_n368__;
  assign new_new_n370__ = ~new_new_n305__ & ~new_new_n364__;
  assign new_new_n371__ = ~new_new_n369__ & new_new_n370__;
  assign new_new_n372__ = ~G169 & ~new_new_n371__;
  assign new_new_n373__ = ~G179 & new_new_n371__;
  assign new_new_n374__ = ~new_new_n363__ & ~new_new_n372__;
  assign new_new_n375__ = ~new_new_n373__ & new_new_n374__;
  assign new_new_n376__ = G190 & new_new_n371__;
  assign new_new_n377__ = G200 & ~new_new_n371__;
  assign new_new_n378__ = new_new_n363__ & ~new_new_n376__;
  assign new_new_n379__ = ~new_new_n377__ & new_new_n378__;
  assign new_new_n380__ = ~new_new_n375__ & ~new_new_n379__;
  assign new_new_n381__ = G20 & ~G68;
  assign new_new_n382__ = ~new_new_n257__ & new_new_n381__;
  assign new_new_n383__ = ~G33 & G50;
  assign new_new_n384__ = ~new_new_n336__ & ~new_new_n383__;
  assign new_new_n385__ = ~G20 & ~new_new_n384__;
  assign new_new_n386__ = ~new_new_n173__ & new_new_n385__;
  assign new_new_n387__ = G68 & ~new_new_n290__;
  assign new_new_n388__ = new_new_n175__ & new_new_n387__;
  assign new_new_n389__ = ~new_new_n382__ & ~new_new_n386__;
  assign new_new_n390__ = ~new_new_n388__ & new_new_n389__;
  assign new_new_n391__ = G238 & new_new_n303__;
  assign new_new_n392__ = G232 & new_new_n150__;
  assign new_new_n393__ = G226 & new_new_n152__;
  assign new_new_n394__ = ~new_new_n193__ & ~new_new_n392__;
  assign new_new_n395__ = ~new_new_n393__ & new_new_n394__;
  assign new_new_n396__ = new_new_n148__ & ~new_new_n395__;
  assign new_new_n397__ = ~new_new_n305__ & ~new_new_n391__;
  assign new_new_n398__ = ~new_new_n396__ & new_new_n397__;
  assign new_new_n399__ = ~G169 & ~new_new_n398__;
  assign new_new_n400__ = ~G179 & new_new_n398__;
  assign new_new_n401__ = ~new_new_n390__ & ~new_new_n399__;
  assign new_new_n402__ = ~new_new_n400__ & new_new_n401__;
  assign new_new_n403__ = G190 & new_new_n398__;
  assign new_new_n404__ = G200 & ~new_new_n398__;
  assign new_new_n405__ = new_new_n390__ & ~new_new_n403__;
  assign new_new_n406__ = ~new_new_n404__ & new_new_n405__;
  assign new_new_n407__ = ~new_new_n402__ & ~new_new_n406__;
  assign new_new_n408__ = new_new_n321__ & new_new_n352__;
  assign new_new_n409__ = new_new_n380__ & new_new_n407__;
  assign new_new_n410__ = new_new_n408__ & new_new_n409__;
  assign G372 = new_new_n287__ & new_new_n410__;
  assign new_new_n412__ = new_new_n186__ & ~new_new_n284__;
  assign new_new_n413__ = ~new_new_n280__ & ~new_new_n412__;
  assign new_new_n414__ = new_new_n256__ & ~new_new_n413__;
  assign new_new_n415__ = ~new_new_n223__ & new_new_n250__;
  assign new_new_n416__ = ~new_new_n219__ & ~new_new_n415__;
  assign new_new_n417__ = ~new_new_n414__ & new_new_n416__;
  assign new_new_n418__ = new_new_n410__ & ~new_new_n417__;
  assign new_new_n419__ = ~new_new_n316__ & ~new_new_n402__;
  assign new_new_n420__ = ~new_new_n406__ & ~new_new_n419__;
  assign new_new_n421__ = ~new_new_n375__ & ~new_new_n420__;
  assign new_new_n422__ = ~new_new_n379__ & ~new_new_n421__;
  assign new_new_n423__ = ~new_new_n347__ & ~new_new_n422__;
  assign new_new_n424__ = ~new_new_n351__ & ~new_new_n423__;
  assign G369 = new_new_n418__ | new_new_n424__;
  assign new_new_n426__ = ~G20 & G213;
  assign new_new_n427__ = new_new_n168__ & new_new_n426__;
  assign new_new_n428__ = G343 & new_new_n427__;
  assign new_new_n429__ = new_new_n280__ & ~new_new_n428__;
  assign new_new_n430__ = new_new_n186__ & ~new_new_n428__;
  assign new_new_n431__ = ~new_new_n267__ & new_new_n428__;
  assign new_new_n432__ = new_new_n285__ & ~new_new_n431__;
  assign new_new_n433__ = new_new_n280__ & new_new_n431__;
  assign new_new_n434__ = ~new_new_n432__ & ~new_new_n433__;
  assign new_new_n435__ = new_new_n430__ & ~new_new_n434__;
  assign new_new_n436__ = ~new_new_n429__ & ~new_new_n435__;
  assign new_new_n437__ = ~new_new_n185__ & new_new_n428__;
  assign new_new_n438__ = new_new_n191__ & ~new_new_n437__;
  assign new_new_n439__ = new_new_n186__ & new_new_n428__;
  assign new_new_n440__ = ~new_new_n438__ & ~new_new_n439__;
  assign new_new_n441__ = G330 & ~new_new_n440__;
  assign new_new_n442__ = ~new_new_n434__ & new_new_n441__;
  assign G399 = ~new_new_n436__ | new_new_n442__;
  assign new_new_n444__ = ~new_new_n417__ & ~new_new_n428__;
  assign new_new_n445__ = ~G179 & ~new_new_n164__;
  assign new_new_n446__ = ~new_new_n215__ & ~new_new_n246__;
  assign new_new_n447__ = ~new_new_n276__ & new_new_n446__;
  assign new_new_n448__ = new_new_n445__ & new_new_n447__;
  assign new_new_n449__ = new_new_n215__ & new_new_n246__;
  assign new_new_n450__ = new_new_n276__ & new_new_n449__;
  assign new_new_n451__ = new_new_n166__ & new_new_n450__;
  assign new_new_n452__ = ~new_new_n448__ & ~new_new_n451__;
  assign new_new_n453__ = new_new_n428__ & ~new_new_n452__;
  assign new_new_n454__ = new_new_n287__ & ~new_new_n428__;
  assign new_new_n455__ = ~new_new_n453__ & ~new_new_n454__;
  assign new_new_n456__ = G330 & ~new_new_n455__;
  assign new_new_n457__ = ~new_new_n444__ & ~new_new_n456__;
  assign new_new_n458__ = ~G1 & ~new_new_n457__;
  assign new_new_n459__ = ~G41 & new_new_n100__;
  assign new_new_n460__ = new_new_n80__ & new_new_n459__;
  assign new_new_n461__ = ~G116 & new_new_n197__;
  assign new_new_n462__ = G1 & ~new_new_n459__;
  assign new_new_n463__ = new_new_n461__ & new_new_n462__;
  assign new_new_n464__ = ~new_new_n460__ & ~new_new_n463__;
  assign G364 = new_new_n458__ | ~new_new_n464__;
  assign new_new_n466__ = G13 & ~G20;
  assign new_new_n467__ = G45 & new_new_n466__;
  assign new_new_n468__ = G1 & ~new_new_n467__;
  assign new_new_n469__ = ~new_new_n459__ & new_new_n468__;
  assign new_new_n470__ = ~G330 & new_new_n440__;
  assign new_new_n471__ = ~new_new_n441__ & ~new_new_n469__;
  assign new_new_n472__ = ~new_new_n470__ & new_new_n471__;
  assign new_new_n473__ = ~G13 & ~G20;
  assign new_new_n474__ = ~G33 & new_new_n473__;
  assign new_new_n475__ = new_new_n440__ & new_new_n474__;
  assign new_new_n476__ = G20 & ~G169;
  assign new_new_n477__ = new_new_n78__ & ~new_new_n476__;
  assign new_new_n478__ = G20 & G179;
  assign new_new_n479__ = G200 & new_new_n478__;
  assign new_new_n480__ = ~G190 & new_new_n479__;
  assign new_new_n481__ = G317 & new_new_n480__;
  assign new_new_n482__ = G20 & ~G190;
  assign new_new_n483__ = G20 & G200;
  assign new_new_n484__ = ~new_new_n478__ & ~new_new_n483__;
  assign new_new_n485__ = new_new_n482__ & new_new_n484__;
  assign new_new_n486__ = G329 & new_new_n485__;
  assign new_new_n487__ = G190 & new_new_n479__;
  assign new_new_n488__ = G326 & new_new_n487__;
  assign new_new_n489__ = ~G200 & new_new_n478__;
  assign new_new_n490__ = ~G190 & new_new_n489__;
  assign new_new_n491__ = G311 & new_new_n490__;
  assign new_new_n492__ = ~new_new_n478__ & new_new_n483__;
  assign new_new_n493__ = G190 & new_new_n492__;
  assign new_new_n494__ = G303 & new_new_n493__;
  assign new_new_n495__ = ~G190 & new_new_n492__;
  assign new_new_n496__ = G283 & new_new_n495__;
  assign new_new_n497__ = ~new_new_n482__ & new_new_n484__;
  assign new_new_n498__ = G294 & new_new_n497__;
  assign new_new_n499__ = G190 & new_new_n489__;
  assign new_new_n500__ = G322 & new_new_n499__;
  assign new_new_n501__ = G33 & ~new_new_n481__;
  assign new_new_n502__ = ~new_new_n486__ & ~new_new_n488__;
  assign new_new_n503__ = ~new_new_n491__ & ~new_new_n494__;
  assign new_new_n504__ = ~new_new_n496__ & ~new_new_n498__;
  assign new_new_n505__ = ~new_new_n500__ & new_new_n504__;
  assign new_new_n506__ = new_new_n502__ & new_new_n503__;
  assign new_new_n507__ = new_new_n501__ & new_new_n506__;
  assign new_new_n508__ = new_new_n505__ & new_new_n507__;
  assign new_new_n509__ = G68 & new_new_n480__;
  assign new_new_n510__ = G77 & new_new_n490__;
  assign new_new_n511__ = G87 & new_new_n493__;
  assign new_new_n512__ = G50 & new_new_n487__;
  assign new_new_n513__ = G107 & new_new_n495__;
  assign new_new_n514__ = G159 & new_new_n485__;
  assign new_new_n515__ = G97 & new_new_n497__;
  assign new_new_n516__ = G58 & new_new_n499__;
  assign new_new_n517__ = ~G33 & ~new_new_n509__;
  assign new_new_n518__ = ~new_new_n510__ & ~new_new_n511__;
  assign new_new_n519__ = ~new_new_n512__ & ~new_new_n513__;
  assign new_new_n520__ = ~new_new_n514__ & ~new_new_n515__;
  assign new_new_n521__ = ~new_new_n516__ & new_new_n520__;
  assign new_new_n522__ = new_new_n518__ & new_new_n519__;
  assign new_new_n523__ = new_new_n517__ & new_new_n522__;
  assign new_new_n524__ = new_new_n521__ & new_new_n523__;
  assign new_new_n525__ = ~new_new_n508__ & ~new_new_n524__;
  assign new_new_n526__ = new_new_n477__ & ~new_new_n525__;
  assign new_new_n527__ = ~new_new_n474__ & ~new_new_n477__;
  assign new_new_n528__ = ~G116 & ~new_new_n100__;
  assign new_new_n529__ = ~G33 & new_new_n100__;
  assign new_new_n530__ = G355 & new_new_n529__;
  assign new_new_n531__ = ~G45 & new_new_n80__;
  assign new_new_n532__ = G33 & new_new_n100__;
  assign new_new_n533__ = G45 & new_new_n134__;
  assign new_new_n534__ = ~new_new_n531__ & new_new_n532__;
  assign new_new_n535__ = ~new_new_n533__ & new_new_n534__;
  assign new_new_n536__ = ~new_new_n528__ & ~new_new_n530__;
  assign new_new_n537__ = ~new_new_n535__ & new_new_n536__;
  assign new_new_n538__ = new_new_n527__ & ~new_new_n537__;
  assign new_new_n539__ = new_new_n469__ & ~new_new_n538__;
  assign new_new_n540__ = ~new_new_n526__ & new_new_n539__;
  assign new_new_n541__ = ~new_new_n475__ & new_new_n540__;
  assign G396 = new_new_n472__ | new_new_n541__;
  assign new_new_n543__ = ~new_new_n300__ & new_new_n428__;
  assign new_new_n544__ = new_new_n321__ & ~new_new_n543__;
  assign new_new_n545__ = new_new_n316__ & new_new_n543__;
  assign new_new_n546__ = ~new_new_n544__ & ~new_new_n545__;
  assign new_new_n547__ = new_new_n444__ & ~new_new_n546__;
  assign new_new_n548__ = ~new_new_n444__ & new_new_n546__;
  assign new_new_n549__ = ~new_new_n547__ & ~new_new_n548__;
  assign new_new_n550__ = new_new_n456__ & new_new_n549__;
  assign new_new_n551__ = ~new_new_n456__ & ~new_new_n549__;
  assign new_new_n552__ = ~new_new_n469__ & ~new_new_n550__;
  assign new_new_n553__ = ~new_new_n551__ & new_new_n552__;
  assign new_new_n554__ = ~G13 & ~G33;
  assign new_new_n555__ = ~new_new_n477__ & ~new_new_n554__;
  assign new_new_n556__ = ~G77 & new_new_n555__;
  assign new_new_n557__ = G150 & new_new_n480__;
  assign new_new_n558__ = G50 & new_new_n493__;
  assign new_new_n559__ = G68 & new_new_n495__;
  assign new_new_n560__ = G159 & new_new_n490__;
  assign new_new_n561__ = G132 & new_new_n485__;
  assign new_new_n562__ = G137 & new_new_n487__;
  assign new_new_n563__ = G58 & new_new_n497__;
  assign new_new_n564__ = G143 & new_new_n499__;
  assign new_new_n565__ = ~G33 & ~new_new_n557__;
  assign new_new_n566__ = ~new_new_n558__ & ~new_new_n559__;
  assign new_new_n567__ = ~new_new_n560__ & ~new_new_n561__;
  assign new_new_n568__ = ~new_new_n562__ & ~new_new_n563__;
  assign new_new_n569__ = ~new_new_n564__ & new_new_n568__;
  assign new_new_n570__ = new_new_n566__ & new_new_n567__;
  assign new_new_n571__ = new_new_n565__ & new_new_n570__;
  assign new_new_n572__ = new_new_n569__ & new_new_n571__;
  assign new_new_n573__ = G107 & new_new_n493__;
  assign new_new_n574__ = G303 & new_new_n487__;
  assign new_new_n575__ = G283 & new_new_n480__;
  assign new_new_n576__ = G294 & new_new_n499__;
  assign new_new_n577__ = G116 & new_new_n490__;
  assign new_new_n578__ = G311 & new_new_n485__;
  assign new_new_n579__ = G87 & new_new_n495__;
  assign new_new_n580__ = G33 & ~new_new_n515__;
  assign new_new_n581__ = ~new_new_n573__ & ~new_new_n574__;
  assign new_new_n582__ = ~new_new_n575__ & ~new_new_n576__;
  assign new_new_n583__ = ~new_new_n577__ & ~new_new_n578__;
  assign new_new_n584__ = ~new_new_n579__ & new_new_n583__;
  assign new_new_n585__ = new_new_n581__ & new_new_n582__;
  assign new_new_n586__ = new_new_n580__ & new_new_n585__;
  assign new_new_n587__ = new_new_n584__ & new_new_n586__;
  assign new_new_n588__ = ~new_new_n572__ & ~new_new_n587__;
  assign new_new_n589__ = new_new_n477__ & ~new_new_n588__;
  assign new_new_n590__ = new_new_n546__ & new_new_n554__;
  assign new_new_n591__ = new_new_n469__ & ~new_new_n556__;
  assign new_new_n592__ = ~new_new_n589__ & new_new_n591__;
  assign new_new_n593__ = ~new_new_n590__ & new_new_n592__;
  assign G384 = new_new_n553__ | new_new_n593__;
  assign new_new_n595__ = new_new_n375__ & ~new_new_n427__;
  assign new_new_n596__ = new_new_n402__ & ~new_new_n428__;
  assign new_new_n597__ = ~new_new_n363__ & new_new_n427__;
  assign new_new_n598__ = new_new_n380__ & ~new_new_n597__;
  assign new_new_n599__ = new_new_n375__ & new_new_n597__;
  assign new_new_n600__ = ~new_new_n598__ & ~new_new_n599__;
  assign new_new_n601__ = new_new_n596__ & ~new_new_n600__;
  assign new_new_n602__ = ~new_new_n390__ & new_new_n428__;
  assign new_new_n603__ = new_new_n407__ & ~new_new_n602__;
  assign new_new_n604__ = new_new_n402__ & new_new_n602__;
  assign new_new_n605__ = ~new_new_n603__ & ~new_new_n604__;
  assign new_new_n606__ = ~new_new_n600__ & ~new_new_n605__;
  assign new_new_n607__ = new_new_n316__ & ~new_new_n428__;
  assign new_new_n608__ = ~new_new_n547__ & ~new_new_n607__;
  assign new_new_n609__ = new_new_n606__ & ~new_new_n608__;
  assign new_new_n610__ = ~new_new_n595__ & ~new_new_n601__;
  assign new_new_n611__ = ~new_new_n609__ & new_new_n610__;
  assign new_new_n612__ = ~new_new_n546__ & new_new_n606__;
  assign new_new_n613__ = ~new_new_n410__ & ~new_new_n612__;
  assign new_new_n614__ = new_new_n410__ & new_new_n612__;
  assign new_new_n615__ = new_new_n456__ & ~new_new_n613__;
  assign new_new_n616__ = ~new_new_n614__ & new_new_n615__;
  assign new_new_n617__ = ~new_new_n611__ & ~new_new_n616__;
  assign new_new_n618__ = new_new_n611__ & new_new_n616__;
  assign new_new_n619__ = ~new_new_n617__ & ~new_new_n618__;
  assign new_new_n620__ = new_new_n410__ & new_new_n444__;
  assign new_new_n621__ = ~new_new_n424__ & ~new_new_n620__;
  assign new_new_n622__ = new_new_n619__ & new_new_n621__;
  assign new_new_n623__ = ~new_new_n619__ & ~new_new_n621__;
  assign new_new_n624__ = ~new_new_n79__ & ~new_new_n99__;
  assign new_new_n625__ = ~new_new_n622__ & new_new_n624__;
  assign new_new_n626__ = ~new_new_n623__ & new_new_n625__;
  assign new_new_n627__ = new_new_n128__ & new_new_n130__;
  assign new_new_n628__ = ~G50 & G68;
  assign new_new_n629__ = ~new_new_n627__ & ~new_new_n628__;
  assign new_new_n630__ = new_new_n99__ & ~new_new_n629__;
  assign new_new_n631__ = G116 & new_new_n78__;
  assign new_new_n632__ = new_new_n232__ & new_new_n631__;
  assign new_new_n633__ = ~new_new_n630__ & ~new_new_n632__;
  assign G367 = new_new_n626__ | ~new_new_n633__;
  assign new_new_n635__ = ~new_new_n204__ & new_new_n428__;
  assign new_new_n636__ = new_new_n224__ & ~new_new_n635__;
  assign new_new_n637__ = new_new_n219__ & new_new_n635__;
  assign new_new_n638__ = ~new_new_n636__ & ~new_new_n637__;
  assign new_new_n639__ = new_new_n474__ & new_new_n638__;
  assign new_new_n640__ = G159 & new_new_n480__;
  assign new_new_n641__ = G50 & new_new_n490__;
  assign new_new_n642__ = G137 & new_new_n485__;
  assign new_new_n643__ = G143 & new_new_n487__;
  assign new_new_n644__ = G58 & new_new_n493__;
  assign new_new_n645__ = G77 & new_new_n495__;
  assign new_new_n646__ = G68 & new_new_n497__;
  assign new_new_n647__ = G150 & new_new_n499__;
  assign new_new_n648__ = ~G33 & ~new_new_n640__;
  assign new_new_n649__ = ~new_new_n641__ & ~new_new_n642__;
  assign new_new_n650__ = ~new_new_n643__ & ~new_new_n644__;
  assign new_new_n651__ = ~new_new_n645__ & ~new_new_n646__;
  assign new_new_n652__ = ~new_new_n647__ & new_new_n651__;
  assign new_new_n653__ = new_new_n649__ & new_new_n650__;
  assign new_new_n654__ = new_new_n648__ & new_new_n653__;
  assign new_new_n655__ = new_new_n652__ & new_new_n654__;
  assign new_new_n656__ = G294 & new_new_n480__;
  assign new_new_n657__ = G116 & new_new_n493__;
  assign new_new_n658__ = G97 & new_new_n495__;
  assign new_new_n659__ = G283 & new_new_n490__;
  assign new_new_n660__ = G317 & new_new_n485__;
  assign new_new_n661__ = G311 & new_new_n487__;
  assign new_new_n662__ = G107 & new_new_n497__;
  assign new_new_n663__ = G303 & new_new_n499__;
  assign new_new_n664__ = G33 & ~new_new_n656__;
  assign new_new_n665__ = ~new_new_n657__ & ~new_new_n658__;
  assign new_new_n666__ = ~new_new_n659__ & ~new_new_n660__;
  assign new_new_n667__ = ~new_new_n661__ & ~new_new_n662__;
  assign new_new_n668__ = ~new_new_n663__ & new_new_n667__;
  assign new_new_n669__ = new_new_n665__ & new_new_n666__;
  assign new_new_n670__ = new_new_n664__ & new_new_n669__;
  assign new_new_n671__ = new_new_n668__ & new_new_n670__;
  assign new_new_n672__ = ~new_new_n655__ & ~new_new_n671__;
  assign new_new_n673__ = new_new_n477__ & ~new_new_n672__;
  assign new_new_n674__ = new_new_n114__ & new_new_n532__;
  assign new_new_n675__ = G87 & ~new_new_n100__;
  assign new_new_n676__ = new_new_n527__ & ~new_new_n675__;
  assign new_new_n677__ = ~new_new_n674__ & new_new_n676__;
  assign new_new_n678__ = new_new_n469__ & ~new_new_n677__;
  assign new_new_n679__ = ~new_new_n673__ & new_new_n678__;
  assign new_new_n680__ = ~new_new_n639__ & new_new_n679__;
  assign new_new_n681__ = ~new_new_n238__ & new_new_n428__;
  assign new_new_n682__ = new_new_n255__ & ~new_new_n681__;
  assign new_new_n683__ = new_new_n250__ & new_new_n681__;
  assign new_new_n684__ = ~new_new_n682__ & ~new_new_n683__;
  assign new_new_n685__ = ~new_new_n436__ & ~new_new_n684__;
  assign new_new_n686__ = new_new_n250__ & ~new_new_n428__;
  assign new_new_n687__ = ~new_new_n685__ & ~new_new_n686__;
  assign new_new_n688__ = new_new_n442__ & ~new_new_n684__;
  assign new_new_n689__ = new_new_n687__ & ~new_new_n688__;
  assign new_new_n690__ = ~new_new_n687__ & new_new_n688__;
  assign new_new_n691__ = ~new_new_n689__ & ~new_new_n690__;
  assign new_new_n692__ = new_new_n638__ & new_new_n691__;
  assign new_new_n693__ = ~new_new_n638__ & ~new_new_n691__;
  assign new_new_n694__ = ~new_new_n692__ & ~new_new_n693__;
  assign new_new_n695__ = ~new_new_n430__ & new_new_n434__;
  assign new_new_n696__ = ~new_new_n435__ & ~new_new_n695__;
  assign new_new_n697__ = new_new_n441__ & new_new_n696__;
  assign new_new_n698__ = ~new_new_n441__ & ~new_new_n696__;
  assign new_new_n699__ = ~new_new_n697__ & ~new_new_n698__;
  assign new_new_n700__ = new_new_n457__ & new_new_n699__;
  assign new_new_n701__ = ~new_new_n436__ & new_new_n442__;
  assign new_new_n702__ = G399 & ~new_new_n701__;
  assign new_new_n703__ = new_new_n684__ & new_new_n702__;
  assign new_new_n704__ = ~new_new_n684__ & ~new_new_n702__;
  assign new_new_n705__ = ~new_new_n703__ & ~new_new_n704__;
  assign new_new_n706__ = new_new_n700__ & ~new_new_n705__;
  assign new_new_n707__ = new_new_n457__ & ~new_new_n706__;
  assign new_new_n708__ = new_new_n459__ & ~new_new_n707__;
  assign new_new_n709__ = new_new_n468__ & ~new_new_n708__;
  assign new_new_n710__ = ~new_new_n694__ & ~new_new_n709__;
  assign G387 = new_new_n680__ | new_new_n710__;
  assign new_new_n712__ = ~new_new_n468__ & new_new_n699__;
  assign new_new_n713__ = ~G107 & ~new_new_n100__;
  assign new_new_n714__ = ~new_new_n461__ & new_new_n529__;
  assign new_new_n715__ = G68 & G77;
  assign new_new_n716__ = ~G45 & ~G50;
  assign new_new_n717__ = G58 & new_new_n716__;
  assign new_new_n718__ = ~new_new_n715__ & new_new_n717__;
  assign new_new_n719__ = new_new_n461__ & new_new_n718__;
  assign new_new_n720__ = G45 & new_new_n123__;
  assign new_new_n721__ = new_new_n532__ & ~new_new_n719__;
  assign new_new_n722__ = ~new_new_n720__ & new_new_n721__;
  assign new_new_n723__ = ~new_new_n713__ & ~new_new_n714__;
  assign new_new_n724__ = ~new_new_n722__ & new_new_n723__;
  assign new_new_n725__ = new_new_n527__ & ~new_new_n724__;
  assign new_new_n726__ = new_new_n434__ & new_new_n474__;
  assign new_new_n727__ = G311 & new_new_n480__;
  assign new_new_n728__ = G326 & new_new_n485__;
  assign new_new_n729__ = G322 & new_new_n487__;
  assign new_new_n730__ = G303 & new_new_n490__;
  assign new_new_n731__ = G294 & new_new_n493__;
  assign new_new_n732__ = G116 & new_new_n495__;
  assign new_new_n733__ = G283 & new_new_n497__;
  assign new_new_n734__ = G317 & new_new_n499__;
  assign new_new_n735__ = G33 & ~new_new_n727__;
  assign new_new_n736__ = ~new_new_n728__ & ~new_new_n729__;
  assign new_new_n737__ = ~new_new_n730__ & ~new_new_n731__;
  assign new_new_n738__ = ~new_new_n732__ & ~new_new_n733__;
  assign new_new_n739__ = ~new_new_n734__ & new_new_n738__;
  assign new_new_n740__ = new_new_n736__ & new_new_n737__;
  assign new_new_n741__ = new_new_n735__ & new_new_n740__;
  assign new_new_n742__ = new_new_n739__ & new_new_n741__;
  assign new_new_n743__ = G68 & new_new_n490__;
  assign new_new_n744__ = G159 & new_new_n487__;
  assign new_new_n745__ = G77 & new_new_n493__;
  assign new_new_n746__ = G58 & new_new_n480__;
  assign new_new_n747__ = G50 & new_new_n499__;
  assign new_new_n748__ = G87 & new_new_n497__;
  assign new_new_n749__ = G150 & new_new_n485__;
  assign new_new_n750__ = ~G33 & ~new_new_n658__;
  assign new_new_n751__ = ~new_new_n743__ & ~new_new_n744__;
  assign new_new_n752__ = ~new_new_n745__ & ~new_new_n746__;
  assign new_new_n753__ = ~new_new_n747__ & ~new_new_n748__;
  assign new_new_n754__ = ~new_new_n749__ & new_new_n753__;
  assign new_new_n755__ = new_new_n751__ & new_new_n752__;
  assign new_new_n756__ = new_new_n750__ & new_new_n755__;
  assign new_new_n757__ = new_new_n754__ & new_new_n756__;
  assign new_new_n758__ = ~new_new_n742__ & ~new_new_n757__;
  assign new_new_n759__ = new_new_n477__ & ~new_new_n758__;
  assign new_new_n760__ = new_new_n469__ & ~new_new_n725__;
  assign new_new_n761__ = ~new_new_n759__ & new_new_n760__;
  assign new_new_n762__ = ~new_new_n726__ & new_new_n761__;
  assign new_new_n763__ = ~new_new_n457__ & ~new_new_n699__;
  assign new_new_n764__ = new_new_n459__ & ~new_new_n700__;
  assign new_new_n765__ = ~new_new_n763__ & new_new_n764__;
  assign new_new_n766__ = ~new_new_n712__ & ~new_new_n762__;
  assign G393 = new_new_n765__ | ~new_new_n766__;
  assign new_new_n768__ = ~new_new_n468__ & ~new_new_n705__;
  assign new_new_n769__ = new_new_n474__ & new_new_n684__;
  assign new_new_n770__ = G294 & new_new_n490__;
  assign new_new_n771__ = G283 & new_new_n493__;
  assign new_new_n772__ = G116 & new_new_n497__;
  assign new_new_n773__ = G317 & new_new_n487__;
  assign new_new_n774__ = G303 & new_new_n480__;
  assign new_new_n775__ = G311 & new_new_n499__;
  assign new_new_n776__ = G322 & new_new_n485__;
  assign new_new_n777__ = G33 & ~new_new_n513__;
  assign new_new_n778__ = ~new_new_n770__ & ~new_new_n771__;
  assign new_new_n779__ = ~new_new_n772__ & ~new_new_n773__;
  assign new_new_n780__ = ~new_new_n774__ & ~new_new_n775__;
  assign new_new_n781__ = ~new_new_n776__ & new_new_n780__;
  assign new_new_n782__ = new_new_n778__ & new_new_n779__;
  assign new_new_n783__ = new_new_n777__ & new_new_n782__;
  assign new_new_n784__ = new_new_n781__ & new_new_n783__;
  assign new_new_n785__ = G58 & new_new_n490__;
  assign new_new_n786__ = G68 & new_new_n493__;
  assign new_new_n787__ = G77 & new_new_n497__;
  assign new_new_n788__ = G150 & new_new_n487__;
  assign new_new_n789__ = G50 & new_new_n480__;
  assign new_new_n790__ = G159 & new_new_n499__;
  assign new_new_n791__ = G143 & new_new_n485__;
  assign new_new_n792__ = ~G33 & ~new_new_n579__;
  assign new_new_n793__ = ~new_new_n785__ & ~new_new_n786__;
  assign new_new_n794__ = ~new_new_n787__ & ~new_new_n788__;
  assign new_new_n795__ = ~new_new_n789__ & ~new_new_n790__;
  assign new_new_n796__ = ~new_new_n791__ & new_new_n795__;
  assign new_new_n797__ = new_new_n793__ & new_new_n794__;
  assign new_new_n798__ = new_new_n792__ & new_new_n797__;
  assign new_new_n799__ = new_new_n796__ & new_new_n798__;
  assign new_new_n800__ = ~new_new_n784__ & ~new_new_n799__;
  assign new_new_n801__ = new_new_n477__ & ~new_new_n800__;
  assign new_new_n802__ = new_new_n143__ & new_new_n532__;
  assign new_new_n803__ = G97 & ~new_new_n100__;
  assign new_new_n804__ = new_new_n527__ & ~new_new_n803__;
  assign new_new_n805__ = ~new_new_n802__ & new_new_n804__;
  assign new_new_n806__ = new_new_n469__ & ~new_new_n805__;
  assign new_new_n807__ = ~new_new_n801__ & new_new_n806__;
  assign new_new_n808__ = ~new_new_n769__ & new_new_n807__;
  assign new_new_n809__ = ~new_new_n700__ & new_new_n705__;
  assign new_new_n810__ = new_new_n459__ & ~new_new_n706__;
  assign new_new_n811__ = ~new_new_n809__ & new_new_n810__;
  assign new_new_n812__ = ~new_new_n768__ & ~new_new_n808__;
  assign G390 = new_new_n811__ | ~new_new_n812__;
  assign new_new_n814__ = ~new_new_n605__ & ~new_new_n608__;
  assign new_new_n815__ = ~new_new_n596__ & ~new_new_n814__;
  assign new_new_n816__ = new_new_n456__ & ~new_new_n546__;
  assign new_new_n817__ = ~new_new_n605__ & new_new_n816__;
  assign new_new_n818__ = new_new_n815__ & ~new_new_n817__;
  assign new_new_n819__ = ~new_new_n815__ & new_new_n817__;
  assign new_new_n820__ = ~new_new_n818__ & ~new_new_n819__;
  assign new_new_n821__ = new_new_n600__ & new_new_n820__;
  assign new_new_n822__ = ~new_new_n600__ & ~new_new_n820__;
  assign new_new_n823__ = ~new_new_n821__ & ~new_new_n822__;
  assign new_new_n824__ = ~new_new_n468__ & ~new_new_n823__;
  assign new_new_n825__ = ~G58 & new_new_n555__;
  assign new_new_n826__ = G137 & new_new_n480__;
  assign new_new_n827__ = G125 & new_new_n485__;
  assign new_new_n828__ = G143 & new_new_n490__;
  assign new_new_n829__ = G150 & new_new_n493__;
  assign new_new_n830__ = G50 & new_new_n495__;
  assign new_new_n831__ = G128 & new_new_n487__;
  assign new_new_n832__ = G159 & new_new_n497__;
  assign new_new_n833__ = G132 & new_new_n499__;
  assign new_new_n834__ = ~G33 & ~new_new_n826__;
  assign new_new_n835__ = ~new_new_n827__ & ~new_new_n828__;
  assign new_new_n836__ = ~new_new_n829__ & ~new_new_n830__;
  assign new_new_n837__ = ~new_new_n831__ & ~new_new_n832__;
  assign new_new_n838__ = ~new_new_n833__ & new_new_n837__;
  assign new_new_n839__ = new_new_n835__ & new_new_n836__;
  assign new_new_n840__ = new_new_n834__ & new_new_n839__;
  assign new_new_n841__ = new_new_n838__ & new_new_n840__;
  assign new_new_n842__ = G107 & new_new_n480__;
  assign new_new_n843__ = G283 & new_new_n487__;
  assign new_new_n844__ = G97 & new_new_n490__;
  assign new_new_n845__ = G294 & new_new_n485__;
  assign new_new_n846__ = G116 & new_new_n499__;
  assign new_new_n847__ = G33 & ~new_new_n511__;
  assign new_new_n848__ = ~new_new_n559__ & ~new_new_n787__;
  assign new_new_n849__ = ~new_new_n842__ & ~new_new_n843__;
  assign new_new_n850__ = ~new_new_n844__ & ~new_new_n845__;
  assign new_new_n851__ = ~new_new_n846__ & new_new_n850__;
  assign new_new_n852__ = new_new_n848__ & new_new_n849__;
  assign new_new_n853__ = new_new_n847__ & new_new_n852__;
  assign new_new_n854__ = new_new_n851__ & new_new_n853__;
  assign new_new_n855__ = ~new_new_n841__ & ~new_new_n854__;
  assign new_new_n856__ = new_new_n477__ & ~new_new_n855__;
  assign new_new_n857__ = new_new_n554__ & new_new_n600__;
  assign new_new_n858__ = new_new_n469__ & ~new_new_n825__;
  assign new_new_n859__ = ~new_new_n856__ & new_new_n858__;
  assign new_new_n860__ = ~new_new_n857__ & new_new_n859__;
  assign new_new_n861__ = new_new_n410__ & ~new_new_n457__;
  assign new_new_n862__ = ~new_new_n424__ & ~new_new_n861__;
  assign new_new_n863__ = new_new_n605__ & ~new_new_n816__;
  assign new_new_n864__ = ~new_new_n817__ & ~new_new_n863__;
  assign new_new_n865__ = new_new_n608__ & new_new_n864__;
  assign new_new_n866__ = ~new_new_n608__ & ~new_new_n864__;
  assign new_new_n867__ = ~new_new_n865__ & ~new_new_n866__;
  assign new_new_n868__ = new_new_n862__ & ~new_new_n867__;
  assign new_new_n869__ = ~new_new_n823__ & new_new_n868__;
  assign new_new_n870__ = new_new_n823__ & ~new_new_n868__;
  assign new_new_n871__ = new_new_n459__ & ~new_new_n869__;
  assign new_new_n872__ = ~new_new_n870__ & new_new_n871__;
  assign new_new_n873__ = ~new_new_n824__ & ~new_new_n860__;
  assign G378 = new_new_n872__ | ~new_new_n873__;
  assign new_new_n875__ = new_new_n862__ & ~new_new_n869__;
  assign new_new_n876__ = new_new_n456__ & new_new_n612__;
  assign new_new_n877__ = new_new_n611__ & ~new_new_n876__;
  assign new_new_n878__ = ~new_new_n611__ & new_new_n876__;
  assign new_new_n879__ = ~new_new_n877__ & ~new_new_n878__;
  assign new_new_n880__ = ~new_new_n334__ & new_new_n427__;
  assign new_new_n881__ = new_new_n352__ & ~new_new_n880__;
  assign new_new_n882__ = new_new_n347__ & new_new_n880__;
  assign new_new_n883__ = ~new_new_n881__ & ~new_new_n882__;
  assign new_new_n884__ = new_new_n879__ & new_new_n883__;
  assign new_new_n885__ = ~new_new_n879__ & ~new_new_n883__;
  assign new_new_n886__ = ~new_new_n884__ & ~new_new_n885__;
  assign new_new_n887__ = new_new_n459__ & ~new_new_n886__;
  assign new_new_n888__ = ~new_new_n875__ & new_new_n887__;
  assign new_new_n889__ = ~new_new_n468__ & ~new_new_n886__;
  assign new_new_n890__ = ~G50 & new_new_n555__;
  assign new_new_n891__ = G41 & ~G50;
  assign new_new_n892__ = G125 & new_new_n487__;
  assign new_new_n893__ = G159 & new_new_n495__;
  assign new_new_n894__ = G128 & new_new_n499__;
  assign new_new_n895__ = G150 & new_new_n497__;
  assign new_new_n896__ = G132 & new_new_n480__;
  assign new_new_n897__ = G124 & new_new_n485__;
  assign new_new_n898__ = G143 & new_new_n493__;
  assign new_new_n899__ = G137 & new_new_n490__;
  assign new_new_n900__ = ~G33 & ~G41;
  assign new_new_n901__ = ~new_new_n892__ & new_new_n900__;
  assign new_new_n902__ = ~new_new_n893__ & ~new_new_n894__;
  assign new_new_n903__ = ~new_new_n895__ & ~new_new_n896__;
  assign new_new_n904__ = ~new_new_n897__ & ~new_new_n898__;
  assign new_new_n905__ = ~new_new_n899__ & new_new_n904__;
  assign new_new_n906__ = new_new_n902__ & new_new_n903__;
  assign new_new_n907__ = new_new_n901__ & new_new_n906__;
  assign new_new_n908__ = new_new_n905__ & new_new_n907__;
  assign new_new_n909__ = G283 & new_new_n485__;
  assign new_new_n910__ = G107 & new_new_n499__;
  assign new_new_n911__ = G58 & new_new_n495__;
  assign new_new_n912__ = G97 & new_new_n480__;
  assign new_new_n913__ = G87 & new_new_n490__;
  assign new_new_n914__ = G116 & new_new_n487__;
  assign new_new_n915__ = G33 & ~G41;
  assign new_new_n916__ = ~new_new_n646__ & new_new_n915__;
  assign new_new_n917__ = ~new_new_n745__ & ~new_new_n909__;
  assign new_new_n918__ = ~new_new_n910__ & ~new_new_n911__;
  assign new_new_n919__ = ~new_new_n912__ & ~new_new_n913__;
  assign new_new_n920__ = ~new_new_n914__ & new_new_n919__;
  assign new_new_n921__ = new_new_n917__ & new_new_n918__;
  assign new_new_n922__ = new_new_n916__ & new_new_n921__;
  assign new_new_n923__ = new_new_n920__ & new_new_n922__;
  assign new_new_n924__ = ~new_new_n891__ & ~new_new_n908__;
  assign new_new_n925__ = ~new_new_n923__ & new_new_n924__;
  assign new_new_n926__ = new_new_n477__ & ~new_new_n925__;
  assign new_new_n927__ = new_new_n554__ & new_new_n883__;
  assign new_new_n928__ = new_new_n469__ & ~new_new_n890__;
  assign new_new_n929__ = ~new_new_n926__ & new_new_n928__;
  assign new_new_n930__ = ~new_new_n927__ & new_new_n929__;
  assign new_new_n931__ = ~new_new_n889__ & ~new_new_n930__;
  assign G375 = new_new_n888__ | ~new_new_n931__;
  assign new_new_n933__ = ~new_new_n468__ & ~new_new_n867__;
  assign new_new_n934__ = ~G68 & new_new_n555__;
  assign new_new_n935__ = G150 & new_new_n490__;
  assign new_new_n936__ = G159 & new_new_n493__;
  assign new_new_n937__ = G132 & new_new_n487__;
  assign new_new_n938__ = G143 & new_new_n480__;
  assign new_new_n939__ = G137 & new_new_n499__;
  assign new_new_n940__ = G50 & new_new_n497__;
  assign new_new_n941__ = G128 & new_new_n485__;
  assign new_new_n942__ = ~G33 & ~new_new_n911__;
  assign new_new_n943__ = ~new_new_n935__ & ~new_new_n936__;
  assign new_new_n944__ = ~new_new_n937__ & ~new_new_n938__;
  assign new_new_n945__ = ~new_new_n939__ & ~new_new_n940__;
  assign new_new_n946__ = ~new_new_n941__ & new_new_n945__;
  assign new_new_n947__ = new_new_n943__ & new_new_n944__;
  assign new_new_n948__ = new_new_n942__ & new_new_n947__;
  assign new_new_n949__ = new_new_n946__ & new_new_n948__;
  assign new_new_n950__ = G283 & new_new_n499__;
  assign new_new_n951__ = G303 & new_new_n485__;
  assign new_new_n952__ = G97 & new_new_n493__;
  assign new_new_n953__ = G116 & new_new_n480__;
  assign new_new_n954__ = G107 & new_new_n490__;
  assign new_new_n955__ = G294 & new_new_n487__;
  assign new_new_n956__ = G33 & ~new_new_n645__;
  assign new_new_n957__ = ~new_new_n748__ & ~new_new_n950__;
  assign new_new_n958__ = ~new_new_n951__ & ~new_new_n952__;
  assign new_new_n959__ = ~new_new_n953__ & ~new_new_n954__;
  assign new_new_n960__ = ~new_new_n955__ & new_new_n959__;
  assign new_new_n961__ = new_new_n957__ & new_new_n958__;
  assign new_new_n962__ = new_new_n956__ & new_new_n961__;
  assign new_new_n963__ = new_new_n960__ & new_new_n962__;
  assign new_new_n964__ = ~new_new_n949__ & ~new_new_n963__;
  assign new_new_n965__ = new_new_n477__ & ~new_new_n964__;
  assign new_new_n966__ = new_new_n554__ & new_new_n605__;
  assign new_new_n967__ = new_new_n469__ & ~new_new_n934__;
  assign new_new_n968__ = ~new_new_n965__ & new_new_n967__;
  assign new_new_n969__ = ~new_new_n966__ & new_new_n968__;
  assign new_new_n970__ = ~new_new_n862__ & new_new_n867__;
  assign new_new_n971__ = new_new_n459__ & ~new_new_n868__;
  assign new_new_n972__ = ~new_new_n970__ & new_new_n971__;
  assign new_new_n973__ = ~new_new_n933__ & ~new_new_n969__;
  assign G381 = new_new_n972__ | ~new_new_n973__;
  assign new_new_n975__ = ~G396 & ~G393;
  assign new_new_n976__ = ~G384 & ~G381;
  assign new_new_n977__ = ~G378 & ~G375;
  assign new_new_n978__ = ~G390 & new_new_n975__;
  assign new_new_n979__ = ~G387 & new_new_n978__;
  assign new_new_n980__ = new_new_n976__ & new_new_n979__;
  assign G407 = ~new_new_n977__ | ~new_new_n980__;
  assign new_new_n982__ = G213 & ~G343;
  assign new_new_n983__ = new_new_n977__ & new_new_n982__;
  assign new_new_n984__ = G213 & G407;
  assign G409 = new_new_n983__ | ~new_new_n984__;
  assign new_new_n986__ = G384 & G381;
  assign new_new_n987__ = ~new_new_n976__ & ~new_new_n986__;
  assign new_new_n988__ = G396 & G393;
  assign new_new_n989__ = ~new_new_n975__ & ~new_new_n988__;
  assign new_new_n990__ = G390 & new_new_n989__;
  assign new_new_n991__ = ~G390 & ~new_new_n989__;
  assign new_new_n992__ = ~new_new_n990__ & ~new_new_n991__;
  assign new_new_n993__ = ~G387 & ~new_new_n992__;
  assign new_new_n994__ = G387 & new_new_n992__;
  assign new_new_n995__ = ~new_new_n993__ & ~new_new_n994__;
  assign new_new_n996__ = new_new_n987__ & new_new_n995__;
  assign new_new_n997__ = ~new_new_n987__ & ~new_new_n995__;
  assign new_new_n998__ = ~new_new_n996__ & ~new_new_n997__;
  assign new_new_n999__ = G378 & G375;
  assign new_new_n1000__ = ~new_new_n977__ & ~new_new_n999__;
  assign new_new_n1001__ = ~new_new_n982__ & ~new_new_n1000__;
  assign new_new_n1002__ = ~G2897 & new_new_n982__;
  assign new_new_n1003__ = ~new_new_n1001__ & ~new_new_n1002__;
  assign new_new_n1004__ = new_new_n998__ & new_new_n1003__;
  assign new_new_n1005__ = ~new_new_n998__ & ~new_new_n1003__;
  assign G405 = new_new_n1004__ | new_new_n1005__;
  assign new_new_n1007__ = new_new_n998__ & new_new_n1000__;
  assign new_new_n1008__ = ~new_new_n998__ & ~new_new_n1000__;
  assign G402 = new_new_n1007__ | new_new_n1008__;
endmodule


