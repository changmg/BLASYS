module mult16_35(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , po0 , po1 , po2 , po3 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ;
  output po0 , po1 , po2 , po3 ;
  wire new_n9, new_n10, new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36, new_n37, new_n38;
  assign new_n9 = pi0 & pi1 ;
  assign new_n10 = ~pi0 & ~pi1 ;
  assign new_n11 = ~new_n9 & ~new_n10 ;
  assign new_n12 = pi2 & new_n11 ;
  assign new_n13 = ~pi2 & ~new_n11 ;
  assign new_n14 = ~new_n12 & ~new_n13 ;
  assign new_n15 = ~new_n9 & ~new_n12 ;
  assign new_n16 = pi5 & ~new_n15 ;
  assign new_n17 = ~pi5 & new_n15 ;
  assign new_n18 = ~new_n16 & ~new_n17 ;
  assign new_n19 = ~pi4 & new_n18 ;
  assign new_n20 = pi4 & ~new_n18 ;
  assign new_n21 = ~new_n19 & ~new_n20 ;
  assign new_n22 = ~pi3 & new_n21 ;
  assign new_n23 = pi3 & ~new_n21 ;
  assign new_n24 = ~new_n22 & ~new_n23 ;
  assign new_n25 = ~pi6 & new_n24 ;
  assign new_n26 = pi6 & ~new_n24 ;
  assign new_n27 = ~new_n25 & ~new_n26 ;
  assign new_n28 = ~new_n16 & ~new_n19 ;
  assign new_n29 = ~pi7 & new_n28 ;
  assign new_n30 = pi7 & ~new_n28 ;
  assign new_n31 = ~new_n29 & ~new_n30 ;
  assign new_n32 = ~new_n22 & ~new_n25 ;
  assign new_n33 = ~new_n31 & ~new_n32 ;
  assign new_n34 = new_n31 & new_n32 ;
  assign new_n35 = ~new_n33 & ~new_n34 ;
  assign new_n36 = ~new_n22 & ~new_n30 ;
  assign new_n37 = ~new_n25 & new_n36 ;
  assign new_n38 = ~new_n29 & ~new_n37 ;
  assign po0 = new_n14 ;
  assign po1 = new_n27 ;
  assign po2 = new_n35 ;
  assign po3 = new_n38 ;
endmodule
