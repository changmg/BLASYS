// Benchmark "ex" written by ABC on Fri Jul  1 14:11:17 2022

module ex ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m,
    F  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m;
  output F;
  assign F = b & e;
endmodule


