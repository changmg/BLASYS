module mult16_49(pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 , pi11 , po00 , po01 , po02 , po03 , po04 , po05 , po06 , po07 , po08 , po09 , po10 , po11 );
  input pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 , pi11 ;
  output po00 , po01 , po02 , po03 , po04 , po05 , po06 , po07 , po08 , po09 , po10 , po11 ;
  wire new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36, new_n37, new_n38, new_n39, new_n40, new_n41, new_n42, new_n43, new_n44, new_n45, new_n46, new_n47, new_n48, new_n49, new_n50, new_n51, new_n52, new_n53, new_n54, new_n55, new_n56, new_n57, new_n58;
  assign new_n13 = pi02 & pi06 ;
  assign new_n14 = pi02 & pi07 ;
  assign new_n15 = pi03 & pi08 ;
  assign new_n16 = pi09 & new_n15 ;
  assign new_n17 = pi03 & pi06 ;
  assign new_n18 = pi00 & pi08 ;
  assign new_n19 = ~new_n17 & ~new_n18 ;
  assign new_n20 = ~new_n16 & ~new_n19 ;
  assign new_n21 = new_n14 & new_n20 ;
  assign new_n22 = ~new_n14 & ~new_n20 ;
  assign new_n23 = ~new_n21 & ~new_n22 ;
  assign new_n24 = pi03 & pi07 ;
  assign new_n25 = pi04 & pi08 ;
  assign new_n26 = pi04 & pi06 ;
  assign new_n27 = pi01 & pi08 ;
  assign new_n28 = ~new_n26 & ~new_n27 ;
  assign new_n29 = ~new_n16 & ~new_n21 ;
  assign new_n30 = pi05 & pi08 ;
  assign new_n31 = pi04 & pi07 ;
  assign new_n32 = new_n13 & new_n30 ;
  assign new_n33 = pi05 & pi06 ;
  assign new_n34 = pi02 & pi08 ;
  assign new_n35 = ~new_n33 & ~new_n34 ;
  assign new_n36 = ~new_n32 & ~new_n35 ;
  assign new_n37 = new_n31 & new_n36 ;
  assign new_n38 = ~new_n31 & ~new_n36 ;
  assign new_n39 = ~new_n37 & ~new_n38 ;
  assign new_n40 = ~new_n32 & ~new_n37 ;
  assign new_n41 = new_n24 & new_n30 ;
  assign new_n42 = pi05 & pi07 ;
  assign new_n43 = ~new_n15 & ~new_n42 ;
  assign new_n44 = ~new_n41 & ~new_n43 ;
  assign new_n45 = ~new_n40 & new_n44 ;
  assign new_n46 = new_n40 & ~new_n44 ;
  assign new_n47 = ~new_n45 & ~new_n46 ;
  assign new_n48 = pi10 & new_n47 ;
  assign new_n49 = ~pi10 & ~new_n47 ;
  assign new_n50 = ~new_n48 & ~new_n49 ;
  assign new_n51 = ~new_n45 & ~new_n48 ;
  assign new_n52 = pi04 & new_n41 ;
  assign new_n53 = ~new_n25 & ~new_n41 ;
  assign new_n54 = ~new_n52 & ~new_n53 ;
  assign new_n55 = pi11 & new_n54 ;
  assign new_n56 = ~pi11 & ~new_n54 ;
  assign new_n57 = ~new_n55 & ~new_n56 ;
  assign new_n58 = ~new_n52 & ~new_n55 ;
  assign po00 = new_n13 ;
  assign po01 = new_n23 ;
  assign po02 = new_n24 ;
  assign po03 = new_n25 ;
  assign po04 = new_n28 ;
  assign po05 = new_n29 ;
  assign po06 = new_n30 ;
  assign po07 = new_n39 ;
  assign po08 = new_n50 ;
  assign po09 = new_n51 ;
  assign po10 = new_n57 ;
  assign po11 = new_n58 ;
endmodule
