module max_10(pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 , pi11 , pi12 , po0 , po1 , po2 , po3 , po4 , po5 , po6 );
  input pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 , pi11 , pi12 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 ;
  wire new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36, new_n37, new_n38, new_n39, new_n40, new_n41, new_n42, new_n43, new_n44;
  assign new_n14 = pi02 & ~pi06 ;
  assign new_n15 = ~pi01 & pi05 ;
  assign new_n16 = ~pi00 & pi04 ;
  assign new_n17 = ~pi09 & ~new_n16 ;
  assign new_n18 = ~pi08 & new_n17 ;
  assign new_n19 = pi01 & ~pi05 ;
  assign new_n20 = pi00 & ~pi04 ;
  assign new_n21 = ~new_n19 & ~new_n20 ;
  assign new_n22 = ~new_n18 & new_n21 ;
  assign new_n23 = ~new_n15 & ~new_n22 ;
  assign new_n24 = ~new_n14 & ~new_n23 ;
  assign new_n25 = ~pi03 & pi07 ;
  assign new_n26 = ~pi02 & pi06 ;
  assign new_n27 = ~new_n25 & ~new_n26 ;
  assign new_n28 = ~new_n24 & new_n27 ;
  assign new_n29 = pi03 & ~pi07 ;
  assign new_n30 = pi00 & pi10 ;
  assign new_n31 = pi04 & ~pi10 ;
  assign new_n32 = ~new_n30 & ~new_n31 ;
  assign new_n33 = pi01 & pi10 ;
  assign new_n34 = pi05 & ~pi10 ;
  assign new_n35 = ~new_n33 & ~new_n34 ;
  assign new_n36 = pi02 & pi10 ;
  assign new_n37 = pi06 & ~pi10 ;
  assign new_n38 = ~new_n36 & ~new_n37 ;
  assign new_n39 = pi03 & pi10 ;
  assign new_n40 = pi07 & ~pi10 ;
  assign new_n41 = ~new_n39 & ~new_n40 ;
  assign new_n42 = ~pi11 & ~pi12 ;
  assign new_n43 = ~pi10 & pi12 ;
  assign new_n44 = ~new_n42 & ~new_n43 ;
  assign po0 = new_n28 ;
  assign po1 = new_n29 ;
  assign po2 = new_n32 ;
  assign po3 = new_n35 ;
  assign po4 = new_n38 ;
  assign po5 = new_n41 ;
  assign po6 = new_n44 ;
endmodule
