module buttfly(\in_0[0] , \in_0[1] , \in_0[2] , \in_0[3] , \in_0[4] , \in_0[5] , \in_0[6] , \in_0[7] , \in_0[8] , \in_0[9] , \in_0[10] , \in_0[11] , \in_0[12] , \in_0[13] , \in_0[14] , \in_0[15] , \in_1[0] , \in_1[1] , \in_1[2] , \in_1[3] , \in_1[4] 
, \in_1[5] , \in_1[6] , \in_1[7] , \in_1[8] , \in_1[9] , \in_1[10] , \in_1[11] , \in_1[12] , \in_1[13] , \in_1[14] , \in_1[15] , \res_0[0] , \res_0[1] , \res_0[2] , \res_0[3] , \res_0[4] , \res_0[5] , \res_0[6] , \res_0[7] , \res_0[8] , \res_0[9] 
, \res_0[10] , \res_0[11] , \res_0[12] , \res_0[13] , \res_0[14] , \res_0[15] , \res_0[16] , \res_1[0] , \res_1[1] , \res_1[2] , \res_1[3] , \res_1[4] , \res_1[5] , \res_1[6] , \res_1[7] , \res_1[8] , \res_1[9] , \res_1[10] , \res_1[11] , \res_1[12] , \res_1[13] 
, \res_1[14] , \res_1[15] , \res_1[16] );
  input \in_0[0] ;
  input \in_0[10] ;
  input \in_0[11] ;
  input \in_0[12] ;
  input \in_0[13] ;
  input \in_0[14] ;
  input \in_0[15] ;
  input \in_0[1] ;
  input \in_0[2] ;
  input \in_0[3] ;
  input \in_0[4] ;
  input \in_0[5] ;
  input \in_0[6] ;
  input \in_0[7] ;
  input \in_0[8] ;
  input \in_0[9] ;
  input \in_1[0] ;
  input \in_1[10] ;
  input \in_1[11] ;
  input \in_1[12] ;
  input \in_1[13] ;
  input \in_1[14] ;
  input \in_1[15] ;
  input \in_1[1] ;
  input \in_1[2] ;
  input \in_1[3] ;
  input \in_1[4] ;
  input \in_1[5] ;
  input \in_1[6] ;
  input \in_1[7] ;
  input \in_1[8] ;
  input \in_1[9] ;
  output \res_0[0] ;
  output \res_0[10] ;
  output \res_0[11] ;
  output \res_0[12] ;
  output \res_0[13] ;
  output \res_0[14] ;
  output \res_0[15] ;
  output \res_0[16] ;
  output \res_0[1] ;
  output \res_0[2] ;
  output \res_0[3] ;
  output \res_0[4] ;
  output \res_0[5] ;
  output \res_0[6] ;
  output \res_0[7] ;
  output \res_0[8] ;
  output \res_0[9] ;
  output \res_1[0] ;
  output \res_1[10] ;
  output \res_1[11] ;
  output \res_1[12] ;
  output \res_1[13] ;
  output \res_1[14] ;
  output \res_1[15] ;
  output \res_1[16] ;
  output \res_1[1] ;
  output \res_1[2] ;
  output \res_1[3] ;
  output \res_1[4] ;
  output \res_1[5] ;
  output \res_1[6] ;
  output \res_1[7] ;
  output \res_1[8] ;
  output \res_1[9] ;
  top U0 ( .pi00( \in_0[0] ) , .pi01( \in_0[1] ) , .pi02( \in_0[2] ) , .pi03( \in_0[3] ) , .pi04( \in_0[4] ) , .pi05( \in_0[5] ) , .pi06( \in_0[6] ) , .pi07( \in_0[7] ) , .pi08( \in_0[8] ) , .pi09( \in_0[9] ) , .pi10( \in_0[10] ) , .pi11( \in_0[11] ) , .pi12( \in_0[12] ) , .pi13( \in_0[13] ) , .pi14( \in_0[14] ) , .pi15( \in_0[15] ) , .pi16( \in_1[0] ) , .pi17( \in_1[1] ) , .pi18( \in_1[2] ) , .pi19( \in_1[3] ) , .pi20( \in_1[4] ) , .pi21( \in_1[5] ) , .pi22( \in_1[6] ) , .pi23( \in_1[7] ) , .pi24( \in_1[8] ) , .pi25( \in_1[9] ) , .pi26( \in_1[10] ) , .pi27( \in_1[11] ) , .pi28( \in_1[12] ) , .pi29( \in_1[13] ) , .pi30( \in_1[14] ) , .pi31( \in_1[15] ) , .po01( \res_0[1] ) , .po02( \res_0[2] ) , .po03( \res_0[3] ) , .po04( \res_0[4] ) , .po05( \res_0[5] ) , .po06( \res_0[6] ) , .po07( \res_0[7] ) , .po08( \res_0[8] ) , .po09( \res_0[9] ) , .po10( \res_0[10] ) , .po11( \res_0[11] ) , .po12( \res_0[12] ) , .po13( \res_0[13] ) , .po14( \res_0[14] ) , .po15( \res_0[15] ) , .po16( \res_0[16] ) , .po17( \res_0[0] ) , .po00( \res_1[0] ) , .po18( \res_1[1] ) , .po19( \res_1[2] ) , .po20( \res_1[3] ) , .po21( \res_1[4] ) , .po22( \res_1[5] ) , .po23( \res_1[6] ) , .po24( \res_1[7] ) , .po25( \res_1[8] ) , .po26( \res_1[9] ) , .po27( \res_1[10] ) , .po28( \res_1[11] ) , .po29( \res_1[12] ) , .po30( \res_1[13] ) , .po31( \res_1[14] ) , .po32( \res_1[15] ) , .po33( \res_1[16] ) );
endmodule

module top(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33;
  wire n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, tpo00, tpo01, tpo02, tpo03, tpo04, tpo05, tpo06, tpo07, tpo08, tpo09, tpo10, tpo11, tpo12, tpo13, tpo14, tpo15, tpo16, tpo18, tpo19, tpo20, tpo21, tpo22, tpo23, tpo24, tpo25, tpo26, tpo27, tpo28, tpo29, tpo30, tpo31, tpo32, tpo33;
  assign po00 = ~tpo00;
  assign po01 = ~tpo01;
  assign po02 = ~tpo02;
  assign po03 = ~tpo03;
  assign po04 = ~tpo04;
  assign po05 = ~tpo05;
  assign po06 = ~tpo06;
  assign po07 = ~tpo07;
  assign po08 = ~tpo08;
  assign po09 = ~tpo09;
  assign po10 = ~tpo10;
  assign po11 = ~tpo11;
  assign po12 = ~tpo12;
  assign po13 = ~tpo13;
  assign po14 = ~tpo14;
  assign po15 = ~tpo15;
  assign po16 = ~tpo16;
  assign po17 = ~tpo00;
  assign po18 = ~tpo18;
  assign po19 = ~tpo19;
  assign po20 = ~tpo20;
  assign po21 = ~tpo21;
  assign po22 = ~tpo22;
  assign po23 = ~tpo23;
  assign po24 = ~tpo24;
  assign po25 = ~tpo25;
  assign po26 = ~tpo26;
  assign po27 = ~tpo27;
  assign po28 = ~tpo28;
  assign po29 = ~tpo29;
  assign po30 = ~tpo30;
  assign po31 = tpo31;
  assign po32 = ~tpo32;
  assign po33 = ~tpo33;
  buttfly_0 U0 ( .pi00( pi13 ), .pi01( pi14 ), .pi02( pi15 ), .pi03( pi29 ), .pi04( pi30 ), .pi05( pi31 ), .pi06( n8 ), .pi07( n9 ), .pi08( n18 ), .pi09( n19 ), .po0( tpo13 ), .po1( tpo14 ), .po2( tpo15 ), .po3( tpo16 ), .po4( tpo30 ), .po5( tpo31 ), .po6( tpo32 ), .po7( tpo33 ) );
  buttfly_1 U1 ( .pi0( pi11 ), .pi1( pi12 ), .pi2( pi27 ), .pi3( pi28 ), .pi4( n6 ), .pi5( n7 ), .pi6( n16 ), .pi7( n17 ), .po0( tpo11 ), .po1( tpo12 ), .po2( n8 ), .po3( n9 ), .po4( tpo28 ), .po5( tpo29 ), .po6( n18 ), .po7( n19 ) );
  buttfly_2 U2 ( .pi00( pi08 ), .pi01( pi09 ), .pi02( pi10 ), .pi03( pi24 ), .pi04( pi25 ), .pi05( pi26 ), .pi06( n4 ), .pi07( n5 ), .pi08( n14 ), .pi09( n15 ), .po00( tpo08 ), .po01( tpo09 ), .po02( tpo10 ), .po03( n6 ), .po04( n7 ), .po05( tpo25 ), .po06( tpo26 ), .po07( tpo27 ), .po08( n16 ), .po09( n17 ) );
  buttfly_3 U3 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi02 ), .pi3( pi16 ), .pi4( pi17 ), .pi5( pi18 ), .po0( tpo00 ), .po1( tpo01 ), .po2( tpo02 ), .po3( n0 ), .po4( n1 ), .po5( tpo18 ), .po6( tpo19 ), .po7( n10 ), .po8( n11 ) );
  buttfly_4 U4 ( .pi00( pi03 ), .pi01( pi04 ), .pi02( pi05 ), .pi03( pi19 ), .pi04( pi20 ), .pi05( pi21 ), .pi06( n0 ), .pi07( n1 ), .pi08( n10 ), .pi09( n11 ), .po00( tpo03 ), .po01( tpo04 ), .po02( tpo05 ), .po03( n2 ), .po04( n3 ), .po05( tpo20 ), .po06( tpo21 ), .po07( tpo22 ), .po08( n12 ), .po09( n13 ) );
  buttfly_5 U5 ( .pi0( pi06 ), .pi1( pi07 ), .pi2( pi22 ), .pi3( pi23 ), .pi4( n2 ), .pi5( n3 ), .pi6( n12 ), .pi7( n13 ), .po0( tpo06 ), .po1( tpo07 ), .po2( n4 ), .po3( n5 ), .po4( tpo23 ), .po5( tpo24 ), .po6( n14 ), .po7( n15 ) );
endmodule
