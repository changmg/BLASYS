module mult8(\A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \B[0] , \B[1] , \B[2] , \B[3] , \B[4] , \B[5] , \B[6] , \B[7] , \O[0] , \O[1] , \O[2] , \O[3] , \O[4] 
, \O[5] , \O[6] , \O[7] , \O[8] , \O[9] , \O[10] , \O[11] , \O[12] , \O[13] , \O[14] , \O[15] );
  input \A[0] ;
  input \A[1] ;
  input \A[2] ;
  input \A[3] ;
  input \A[4] ;
  input \A[5] ;
  input \A[6] ;
  input \A[7] ;
  input \B[0] ;
  input \B[1] ;
  input \B[2] ;
  input \B[3] ;
  input \B[4] ;
  input \B[5] ;
  input \B[6] ;
  input \B[7] ;
  output \O[0] ;
  output \O[10] ;
  output \O[11] ;
  output \O[12] ;
  output \O[13] ;
  output \O[14] ;
  output \O[15] ;
  output \O[1] ;
  output \O[2] ;
  output \O[3] ;
  output \O[4] ;
  output \O[5] ;
  output \O[6] ;
  output \O[7] ;
  output \O[8] ;
  output \O[9] ;
  top U0 ( .pi00( \A[0] ) , .pi01( \A[1] ) , .pi02( \A[2] ) , .pi03( \A[3] ) , .pi04( \A[4] ) , .pi05( \A[5] ) , .pi06( \A[6] ) , .pi07( \A[7] ) , .pi08( \B[0] ) , .pi09( \B[1] ) , .pi10( \B[2] ) , .pi11( \B[3] ) , .pi12( \B[4] ) , .pi13( \B[5] ) , .pi14( \B[6] ) , .pi15( \B[7] ) , .po00( \O[0] ) , .po01( \O[1] ) , .po02( \O[2] ) , .po03( \O[3] ) , .po04( \O[4] ) , .po05( \O[5] ) , .po06( \O[6] ) , .po07( \O[7] ) , .po08( \O[8] ) , .po09( \O[9] ) , .po10( \O[10] ) , .po11( \O[11] ) , .po12( \O[12] ) , .po13( \O[13] ) , .po14( \O[14] ) , .po15( \O[15] ) );
endmodule

module top(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15;
  wire n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, tpo00, tpo01, tpo02, tpo03, tpo04, tpo05, tpo06, tpo07, tpo08, tpo09, tpo10, tpo11, tpo12, tpo13, tpo14, tpo15;
  assign po00 = tpo00;
  assign po01 = tpo01;
  assign po02 = ~tpo02;
  assign po03 = ~tpo03;
  assign po04 = ~tpo04;
  assign po05 = ~tpo05;
  assign po06 = ~tpo06;
  assign po07 = ~tpo07;
  assign po08 = tpo08;
  assign po09 = ~tpo09;
  assign po10 = ~tpo10;
  assign po11 = ~tpo11;
  assign po12 = tpo12;
  assign po13 = ~tpo13;
  assign po14 = tpo14;
  assign po15 = tpo15;
  mult8_0 U0 ( .pi0( n28 ), .pi1( n29 ), .pi2( n30 ), .pi3( n31 ), .pi4( n37 ), .pi5( n38 ), .po0( n32 ), .po1( n33 ), .po2( n39 ), .po3( n40 ), .po4( n41 ) );
  mult8_1 U1 ( .pi0( pi03 ), .pi1( pi04 ), .pi2( pi08 ), .pi3( pi09 ), .pi4( pi10 ), .pi5( pi11 ), .pi6( n7 ), .pi7( n18 ), .po00(  ), .po01(  ), .po02(  ), .po03(  ), .po04( n0 ), .po05( n3 ), .po06( n4 ), .po07( n8 ), .po08( n9 ), .po09( n11 ), .po10( n17 ), .po11( n19 ), .po12( n21 ), .po13( n30 ), .po14( n31 ) );
  mult8_2 U2 ( .pi0( pi05 ), .pi1( pi06 ), .pi2( pi07 ), .pi3( pi08 ), .pi4( pi09 ), .pi5( pi10 ), .pi6( pi11 ), .pi7( n8 ), .pi8( n17 ), .po00(  ), .po01( n7 ), .po02( n18 ), .po03( n28 ), .po04( n29 ), .po05( n37 ), .po06( n38 ), .po07( n51 ), .po08( n52 ), .po09( n59 ), .po10( n60 ) );
  mult8_3 U3 ( .pi0( n13 ), .pi1( n14 ), .pi2( n15 ), .pi3( n16 ), .pi4( n19 ), .pi5( n20 ), .pi6( n21 ), .pi7( n22 ), .pi8( n23 ), .po0( tpo05 ), .po1( n24 ), .po2( n25 ), .po3( n26 ), .po4( n27 ) );
  mult8_4 U4 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi02 ), .pi3( pi08 ), .pi4( pi09 ), .pi5( pi10 ), .pi6( n0 ), .pi7( n3 ), .pi8( n4 ), .po00(  ), .po01(  ), .po02( tpo00 ), .po03( tpo01 ), .po04( tpo02 ), .po05( n1 ), .po06( n2 ), .po07( n5 ), .po08( n6 ), .po09( n10 ), .po10( n12 ) );
  mult8_5 U5 ( .pi00( pi00 ), .pi01( pi01 ), .pi02( pi02 ), .pi03( pi11 ), .pi04( pi12 ), .pi05( pi13 ), .pi06( n1 ), .pi07( n2 ), .pi08( n5 ), .pi09( n6 ), .pi10( n9 ), .pi11( n10 ), .pi12( n11 ), .pi13( n12 ), .po00(  ), .po01(  ), .po02( tpo03 ), .po03( tpo04 ), .po04( n13 ), .po05( n14 ), .po06( n15 ), .po07( n16 ), .po08( n20 ), .po09( n22 ), .po10( n23 ) );
  mult8_6 U6 ( .pi0( n27 ), .pi1( n32 ), .pi2( n33 ), .pi3( n34 ), .pi4( n41 ), .pi5( n42 ), .pi6( n44 ), .po0( n35 ), .po1( n36 ), .po2( n43 ), .po3( n50 ) );
  mult8_7 U7 ( .pi00( pi00 ), .pi01( pi01 ), .pi02( pi02 ), .pi03( pi03 ), .pi04( pi13 ), .pi05( pi14 ), .pi06( pi15 ), .pi07( n24 ), .pi08( n25 ), .pi09( n26 ), .pi10( n35 ), .pi11( n36 ), .pi12( n43 ), .po00(  ), .po01(  ), .po02(  ), .po03(  ), .po04( tpo06 ), .po05( tpo07 ), .po06( n44 ), .po07( n45 ), .po08( n46 ), .po09( n47 ), .po10( n48 ), .po11( n49 ), .po12( n55 ), .po13( n56 ) );
  mult8_8 U8 ( .pi00( n45 ), .pi01( n46 ), .pi02( n47 ), .pi03( n48 ), .pi04( n49 ), .pi05( n50 ), .pi06( n53 ), .pi07( n54 ), .pi08( n55 ), .pi09( n56 ), .po0( tpo08 ), .po1( tpo09 ), .po2( n57 ), .po3( n58 ), .po4( n68 ) );
  mult8_9 U9 ( .pi00( pi03 ), .pi01( pi04 ), .pi02( pi05 ), .pi03( pi06 ), .pi04( pi07 ), .pi05( pi12 ), .pi06( pi13 ), .pi07( pi14 ), .pi08( pi15 ), .pi09( n39 ), .pi10( n40 ), .pi11( n51 ), .pi12( n52 ), .pi13( n59 ), .pi14( n60 ), .po00(  ), .po01( n34 ), .po02( n42 ), .po03( n53 ), .po04( n54 ), .po05( n61 ), .po06( n62 ), .po07( n63 ), .po08( n64 ), .po09( n67 ), .po10( n70 ), .po11( n71 ), .po12( n72 ), .po13( n73 ), .po14( n74 ), .po15( n75 ) );
  mult8_10 U10 ( .pi0( pi05 ), .pi1( pi06 ), .pi2( pi07 ), .pi3( pi14 ), .pi4( pi15 ), .pi5( n70 ), .pi6( n74 ), .pi7( n75 ), .pi8( n78 ), .po0(  ), .po1(  ), .po2( n76 ), .po3( n77 ), .po4( tpo13 ), .po5( tpo14 ), .po6( tpo15 ) );
  mult8_11 U11 ( .pi00( n57 ), .pi01( n65 ), .pi02( n66 ), .pi03( n67 ), .pi04( n68 ), .pi05( n69 ), .pi06( n71 ), .pi07( n72 ), .pi08( n73 ), .pi09( n76 ), .pi10( n77 ), .po0( tpo10 ), .po1( tpo11 ), .po2( n78 ), .po3( tpo12 ) );
  mult8_12 U12 ( .pi0( n58 ), .pi1( n61 ), .pi2( n62 ), .pi3( n63 ), .pi4( n64 ), .po0( n65 ), .po1( n66 ), .po2( n69 ) );
endmodule
