module max_50_2(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , po0 , po1 , po2 , po3 , po4 , po5 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 ;
  output po0 , po1 , po2 , po3 , po4 , po5 ;
  wire new_n7, new_n8, new_n9, new_n10, new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18;
  assign new_n7 = pi0 & ~pi2 ;
  assign new_n8 = pi1 & ~pi3 ;
  assign new_n9 = ~pi0 & pi2 ;
  assign new_n10 = ~pi5 & ~new_n9 ;
  assign new_n11 = ~new_n8 & ~new_n10 ;
  assign new_n12 = ~pi1 & pi3 ;
  assign new_n13 = pi0 & pi4 ;
  assign new_n14 = pi2 & ~pi4 ;
  assign new_n15 = ~new_n13 & ~new_n14 ;
  assign new_n16 = pi1 & pi4 ;
  assign new_n17 = pi3 & ~pi4 ;
  assign new_n18 = ~new_n16 & ~new_n17 ;
  assign po0 = pi4 ;
  assign po1 = new_n7 ;
  assign po2 = new_n11 ;
  assign po3 = new_n12 ;
  assign po4 = new_n15 ;
  assign po5 = new_n18 ;
endmodule
