module mult8_9(pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 , pi11 , pi12 , pi13 , pi14 , po00 , po01 , po02 , po03 , po04 , po05 , po06 , po07 , po08 , po09 , po10 , po11 , po12 , po13 , po14 , po15 );
  input pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 , pi11 , pi12 , pi13 , pi14 ;
  output po00 , po01 , po02 , po03 , po04 , po05 , po06 , po07 , po08 , po09 , po10 , po11 , po12 , po13 , po14 , po15 ;
  wire new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36, new_n37, new_n38, new_n39, new_n40, new_n41, new_n42, new_n43, new_n44, new_n45, new_n46, new_n47, new_n48, new_n49, new_n50, new_n51, new_n52, new_n53, new_n54, new_n55, new_n56, new_n57, new_n58, new_n59, new_n60, new_n61, new_n62, new_n63, new_n64, new_n65, new_n66, new_n67, new_n68, new_n69, new_n70, new_n71, new_n72, new_n73, new_n74, new_n75, new_n76, new_n77, new_n78, new_n79;
  assign new_n16 = pi00 & pi05 ;
  assign new_n17 = pi01 & pi05 ;
  assign new_n18 = ~pi10 & new_n17 ;
  assign new_n19 = ~pi09 & ~new_n18 ;
  assign new_n20 = pi11 & ~pi12 ;
  assign new_n21 = ~pi11 & pi12 ;
  assign new_n22 = ~new_n20 & ~new_n21 ;
  assign new_n23 = pi02 & pi05 ;
  assign new_n24 = new_n22 & ~new_n23 ;
  assign new_n25 = ~new_n22 & new_n23 ;
  assign new_n26 = ~new_n24 & ~new_n25 ;
  assign new_n27 = ~new_n19 & ~new_n26 ;
  assign new_n28 = ~new_n22 & ~new_n23 ;
  assign new_n29 = new_n22 & new_n23 ;
  assign new_n30 = ~new_n28 & ~new_n29 ;
  assign new_n31 = new_n19 & ~new_n30 ;
  assign new_n32 = ~new_n27 & ~new_n31 ;
  assign new_n33 = pi01 & pi06 ;
  assign new_n34 = new_n32 & ~new_n33 ;
  assign new_n35 = ~new_n32 & new_n33 ;
  assign new_n36 = ~new_n34 & ~new_n35 ;
  assign new_n37 = ~new_n32 & ~new_n33 ;
  assign new_n38 = new_n32 & new_n33 ;
  assign new_n39 = ~new_n37 & ~new_n38 ;
  assign new_n40 = ~pi13 & ~pi14 ;
  assign new_n41 = pi03 & pi05 ;
  assign new_n42 = ~new_n40 & ~new_n41 ;
  assign new_n43 = new_n40 & new_n41 ;
  assign new_n44 = ~new_n42 & ~new_n43 ;
  assign new_n45 = ~new_n21 & new_n23 ;
  assign new_n46 = ~new_n20 & ~new_n45 ;
  assign new_n47 = ~new_n44 & new_n46 ;
  assign new_n48 = new_n40 & ~new_n41 ;
  assign new_n49 = ~new_n40 & new_n41 ;
  assign new_n50 = ~new_n48 & ~new_n49 ;
  assign new_n51 = ~new_n46 & ~new_n50 ;
  assign new_n52 = ~new_n47 & ~new_n51 ;
  assign new_n53 = pi02 & pi06 ;
  assign new_n54 = ~new_n31 & new_n33 ;
  assign new_n55 = ~new_n27 & ~new_n54 ;
  assign new_n56 = pi01 & pi07 ;
  assign new_n57 = pi00 & pi08 ;
  assign new_n58 = pi04 & pi05 ;
  assign new_n59 = ~pi13 & ~new_n58 ;
  assign new_n60 = pi03 & pi06 ;
  assign new_n61 = ~new_n59 & new_n60 ;
  assign new_n62 = ~pi14 & new_n41 ;
  assign new_n63 = ~new_n59 & ~new_n62 ;
  assign new_n64 = ~new_n60 & ~new_n63 ;
  assign new_n65 = new_n61 & ~new_n62 ;
  assign new_n66 = ~new_n64 & ~new_n65 ;
  assign new_n67 = ~new_n47 & new_n53 ;
  assign new_n68 = ~new_n51 & ~new_n67 ;
  assign new_n69 = new_n66 & ~new_n68 ;
  assign new_n70 = ~new_n51 & ~new_n53 ;
  assign new_n71 = ~new_n47 & ~new_n70 ;
  assign new_n72 = ~new_n66 & ~new_n71 ;
  assign new_n73 = ~new_n69 & ~new_n72 ;
  assign new_n74 = pi02 & pi07 ;
  assign new_n75 = pi01 & pi08 ;
  assign new_n76 = pi04 & pi06 ;
  assign new_n77 = ~new_n62 & ~new_n76 ;
  assign new_n78 = ~new_n72 & new_n74 ;
  assign new_n79 = ~new_n69 & ~new_n78 ;
  assign po00 = pi01 ;
  assign po01 = new_n16 ;
  assign po02 = new_n17 ;
  assign po03 = new_n36 ;
  assign po04 = new_n39 ;
  assign po05 = new_n52 ;
  assign po06 = new_n53 ;
  assign po07 = new_n55 ;
  assign po08 = new_n56 ;
  assign po09 = new_n57 ;
  assign po10 = new_n61 ;
  assign po11 = new_n73 ;
  assign po12 = new_n74 ;
  assign po13 = new_n75 ;
  assign po14 = new_n77 ;
  assign po15 = new_n79 ;
endmodule
