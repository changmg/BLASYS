module mac_2(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 , po0 , po1 , po2 , po3 , po4 , po5 , po6 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 ;
  wire new_n10, new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36, new_n37, new_n38, new_n39, new_n40, new_n41, new_n42, new_n43, new_n44, new_n45, new_n46, new_n47, new_n48, new_n49, new_n50, new_n51, new_n52;
  assign new_n10 = pi0 & pi2 ;
  assign new_n11 = pi5 & new_n10 ;
  assign new_n12 = ~pi5 & ~new_n10 ;
  assign new_n13 = ~new_n11 & ~new_n12 ;
  assign new_n14 = pi1 & pi2 ;
  assign new_n15 = pi6 & new_n14 ;
  assign new_n16 = ~pi6 & ~new_n14 ;
  assign new_n17 = ~new_n15 & ~new_n16 ;
  assign new_n18 = ~new_n11 & ~new_n17 ;
  assign new_n19 = new_n11 & new_n17 ;
  assign new_n20 = ~new_n18 & ~new_n19 ;
  assign new_n21 = pi0 & pi3 ;
  assign new_n22 = new_n20 & new_n21 ;
  assign new_n23 = ~new_n20 & ~new_n21 ;
  assign new_n24 = ~new_n22 & ~new_n23 ;
  assign new_n25 = pi1 & pi3 ;
  assign new_n26 = ~new_n19 & ~new_n22 ;
  assign new_n27 = pi7 & new_n15 ;
  assign new_n28 = ~pi7 & ~new_n15 ;
  assign new_n29 = ~new_n27 & ~new_n28 ;
  assign new_n30 = new_n25 & new_n29 ;
  assign new_n31 = ~new_n25 & ~new_n29 ;
  assign new_n32 = ~new_n30 & ~new_n31 ;
  assign new_n33 = new_n26 & ~new_n32 ;
  assign new_n34 = ~new_n26 & new_n32 ;
  assign new_n35 = ~new_n33 & ~new_n34 ;
  assign new_n36 = pi0 & pi4 ;
  assign new_n37 = new_n35 & new_n36 ;
  assign new_n38 = ~new_n35 & ~new_n36 ;
  assign new_n39 = ~new_n37 & ~new_n38 ;
  assign new_n40 = pi1 & pi4 ;
  assign new_n41 = ~new_n27 & ~new_n30 ;
  assign new_n42 = pi8 & ~new_n41 ;
  assign new_n43 = ~pi8 & new_n41 ;
  assign new_n44 = ~new_n42 & ~new_n43 ;
  assign new_n45 = ~new_n40 & ~new_n44 ;
  assign new_n46 = new_n40 & new_n44 ;
  assign new_n47 = ~new_n45 & ~new_n46 ;
  assign new_n48 = ~new_n34 & ~new_n37 ;
  assign new_n49 = new_n47 & ~new_n48 ;
  assign new_n50 = ~new_n47 & new_n48 ;
  assign new_n51 = ~new_n49 & ~new_n50 ;
  assign new_n52 = ~new_n42 & ~new_n46 ;
  assign po0 = new_n13 ;
  assign po1 = new_n24 ;
  assign po2 = new_n25 ;
  assign po3 = new_n39 ;
  assign po4 = new_n49 ;
  assign po5 = new_n51 ;
  assign po6 = new_n52 ;
endmodule
