module max_31_1(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , po0 , po1 , po2 , po3 , po4 , po5 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ;
  output po0 , po1 , po2 , po3 , po4 , po5 ;
  wire new_n9, new_n10, new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27;
  assign new_n9 = pi0 & ~pi3 ;
  assign new_n10 = ~pi0 & pi3 ;
  assign new_n11 = ~pi1 & pi4 ;
  assign new_n12 = ~new_n10 & ~new_n11 ;
  assign new_n13 = ~pi6 & new_n12 ;
  assign new_n14 = pi2 & ~pi5 ;
  assign new_n15 = pi1 & ~pi4 ;
  assign new_n16 = ~new_n14 & ~new_n15 ;
  assign new_n17 = ~new_n13 & new_n16 ;
  assign new_n18 = ~pi2 & pi5 ;
  assign new_n19 = pi0 & pi7 ;
  assign new_n20 = pi3 & ~pi7 ;
  assign new_n21 = ~new_n19 & ~new_n20 ;
  assign new_n22 = pi1 & pi7 ;
  assign new_n23 = pi4 & ~pi7 ;
  assign new_n24 = ~new_n22 & ~new_n23 ;
  assign new_n25 = pi2 & pi7 ;
  assign new_n26 = pi5 & ~pi7 ;
  assign new_n27 = ~new_n25 & ~new_n26 ;
  assign po0 = new_n9 ;
  assign po1 = new_n17 ;
  assign po2 = new_n18 ;
  assign po3 = new_n21 ;
  assign po4 = new_n24 ;
  assign po5 = new_n27 ;
endmodule
