// Benchmark "c2670" written by ABC on Sat Jul 16 14:42:52 2022

module c2670 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35;
  wire new_n192_, new_n193_, new_n195_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n208_, new_n209_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n218_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n248_, new_n249_, new_n251_, new_n252_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n327_,
    new_n328_, new_n330_, new_n332_, new_n333_, new_n334_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n769_;
  assign new_n192_ = pi136 & pi137;
  assign new_n193_ = pi138 & pi139;
  assign po00 = ~new_n192_ | ~new_n193_;
  assign new_n195_ = pi001 & pi010;
  assign po01 = ~pi120 | ~new_n195_;
  assign po02 = pi073 & pi114;
  assign po03 = ~pi006 | ~pi120;
  assign po04 = ~pi118 | po03;
  assign po05 = ~pi144 | po03;
  assign new_n201_ = pi042 & pi052;
  assign new_n202_ = pi085 & pi095;
  assign new_n203_ = new_n201_ & new_n202_;
  assign new_n204_ = pi031 & pi063;
  assign new_n205_ = pi075 & pi105;
  assign new_n206_ = new_n204_ & new_n205_;
  assign po06 = new_n203_ & new_n206_;
  assign new_n208_ = pi144 & ~new_n206_;
  assign new_n209_ = pi118 & ~new_n203_;
  assign po07 = ~new_n208_ & ~new_n209_;
  assign new_n211_ = pi088 & pi142;
  assign new_n212_ = pi098 & ~pi142;
  assign new_n213_ = pi143 & ~new_n212_;
  assign new_n214_ = ~new_n211_ & new_n213_;
  assign new_n215_ = pi078 & pi142;
  assign new_n216_ = pi108 & ~pi142;
  assign new_n217_ = ~pi143 & ~new_n216_;
  assign new_n218_ = ~new_n215_ & new_n217_;
  assign po08 = new_n214_ | new_n218_;
  assign new_n220_ = pi087 & pi142;
  assign new_n221_ = pi097 & ~pi142;
  assign new_n222_ = pi143 & ~new_n221_;
  assign new_n223_ = ~new_n220_ & new_n222_;
  assign new_n224_ = pi077 & pi142;
  assign new_n225_ = pi107 & ~pi142;
  assign new_n226_ = ~pi143 & ~new_n225_;
  assign new_n227_ = ~new_n224_ & new_n226_;
  assign po09 = new_n223_ | new_n227_;
  assign new_n229_ = pi089 & pi142;
  assign new_n230_ = pi099 & ~pi142;
  assign new_n231_ = pi143 & ~new_n230_;
  assign new_n232_ = ~new_n229_ & new_n231_;
  assign new_n233_ = pi079 & pi142;
  assign new_n234_ = pi109 & ~pi142;
  assign new_n235_ = ~pi143 & ~new_n234_;
  assign new_n236_ = ~new_n233_ & new_n235_;
  assign po10 = new_n232_ | new_n236_;
  assign new_n238_ = pi051 & pi116;
  assign new_n239_ = pi041 & ~pi116;
  assign new_n240_ = pi119 & ~new_n239_;
  assign new_n241_ = ~new_n238_ & new_n240_;
  assign new_n242_ = pi030 & pi116;
  assign new_n243_ = pi062 & ~pi116;
  assign new_n244_ = ~pi119 & ~new_n243_;
  assign new_n245_ = ~new_n242_ & new_n244_;
  assign new_n246_ = ~new_n241_ & ~new_n245_;
  assign po11 = ~pi121 | new_n246_;
  assign new_n248_ = pi115 & pi120;
  assign new_n249_ = pi027 & new_n248_;
  assign po12 = ~po07 | ~new_n249_;
  assign new_n251_ = pi000 & pi002;
  assign new_n252_ = new_n248_ & ~new_n251_;
  assign po13 = ~po07 | ~new_n252_;
  assign new_n254_ = pi059 & pi116;
  assign new_n255_ = pi048 & ~pi116;
  assign new_n256_ = pi119 & ~new_n255_;
  assign new_n257_ = ~new_n254_ & new_n256_;
  assign new_n258_ = pi038 & pi116;
  assign new_n259_ = pi070 & ~pi116;
  assign new_n260_ = ~pi119 & ~new_n259_;
  assign new_n261_ = ~new_n258_ & new_n260_;
  assign po14 = ~new_n257_ & ~new_n261_;
  assign new_n263_ = pi058 & pi116;
  assign new_n264_ = pi047 & ~pi116;
  assign new_n265_ = pi119 & ~new_n264_;
  assign new_n266_ = ~new_n263_ & new_n265_;
  assign new_n267_ = pi037 & pi116;
  assign new_n268_ = pi069 & ~pi116;
  assign new_n269_ = ~pi119 & ~new_n268_;
  assign new_n270_ = ~new_n267_ & new_n269_;
  assign po15 = ~new_n266_ & ~new_n270_;
  assign new_n272_ = pi057 & pi116;
  assign new_n273_ = pi046 & ~pi116;
  assign new_n274_ = pi119 & ~new_n273_;
  assign new_n275_ = ~new_n272_ & new_n274_;
  assign new_n276_ = pi036 & pi116;
  assign new_n277_ = pi068 & ~pi116;
  assign new_n278_ = ~pi119 & ~new_n277_;
  assign new_n279_ = ~new_n276_ & new_n278_;
  assign po16 = ~new_n275_ & ~new_n279_;
  assign new_n281_ = pi056 & pi116;
  assign new_n282_ = pi045 & ~pi116;
  assign new_n283_ = pi119 & ~new_n282_;
  assign new_n284_ = ~new_n281_ & new_n283_;
  assign new_n285_ = pi035 & pi116;
  assign new_n286_ = pi067 & ~pi116;
  assign new_n287_ = ~pi119 & ~new_n286_;
  assign new_n288_ = ~new_n285_ & new_n287_;
  assign po17 = ~new_n284_ & ~new_n288_;
  assign new_n290_ = pi055 & pi119;
  assign new_n291_ = pi034 & ~pi119;
  assign new_n292_ = pi116 & ~new_n291_;
  assign new_n293_ = ~new_n290_ & new_n292_;
  assign new_n294_ = ~pi066 & ~pi116;
  assign new_n295_ = ~pi119 & new_n294_;
  assign po18 = ~new_n293_ & ~new_n295_;
  assign new_n297_ = pi054 & pi116;
  assign new_n298_ = pi044 & ~pi116;
  assign new_n299_ = pi119 & ~new_n298_;
  assign new_n300_ = ~new_n297_ & new_n299_;
  assign new_n301_ = pi033 & pi116;
  assign new_n302_ = pi065 & ~pi116;
  assign new_n303_ = ~pi119 & ~new_n302_;
  assign new_n304_ = ~new_n301_ & new_n303_;
  assign po19 = ~new_n300_ & ~new_n304_;
  assign new_n306_ = pi053 & pi116;
  assign new_n307_ = pi043 & ~pi116;
  assign new_n308_ = pi119 & ~new_n307_;
  assign new_n309_ = ~new_n306_ & new_n308_;
  assign new_n310_ = pi032 & pi116;
  assign new_n311_ = pi064 & ~pi116;
  assign new_n312_ = ~pi119 & ~new_n311_;
  assign new_n313_ = ~new_n310_ & new_n312_;
  assign po20 = ~new_n309_ & ~new_n313_;
  assign new_n315_ = pi122 & ~po15;
  assign new_n316_ = pi060 & pi116;
  assign new_n317_ = pi049 & ~pi116;
  assign new_n318_ = pi119 & ~new_n317_;
  assign new_n319_ = ~new_n316_ & new_n318_;
  assign new_n320_ = pi039 & pi116;
  assign new_n321_ = pi071 & ~pi116;
  assign new_n322_ = ~pi119 & ~new_n321_;
  assign new_n323_ = ~new_n320_ & new_n322_;
  assign new_n324_ = ~new_n319_ & ~new_n323_;
  assign new_n325_ = ~pi122 & ~new_n324_;
  assign po21 = ~new_n315_ & ~new_n325_;
  assign new_n327_ = pi122 & ~po16;
  assign new_n328_ = ~pi122 & ~po14;
  assign po22 = ~new_n327_ & ~new_n328_;
  assign new_n330_ = pi117 & ~pi121;
  assign po23 = new_n324_ | new_n330_;
  assign new_n332_ = ~pi117 & ~new_n324_;
  assign new_n333_ = pi122 & ~new_n332_;
  assign new_n334_ = ~pi122 & new_n246_;
  assign po24 = new_n333_ | new_n334_;
  assign new_n336_ = pi086 & pi142;
  assign new_n337_ = pi096 & ~pi142;
  assign new_n338_ = pi143 & ~new_n337_;
  assign new_n339_ = ~new_n336_ & new_n338_;
  assign new_n340_ = pi076 & pi142;
  assign new_n341_ = pi106 & ~pi142;
  assign new_n342_ = ~pi143 & ~new_n341_;
  assign new_n343_ = ~new_n340_ & new_n342_;
  assign new_n344_ = ~new_n339_ & ~new_n343_;
  assign new_n345_ = pi140 & new_n344_;
  assign new_n346_ = ~pi140 & ~new_n344_;
  assign new_n347_ = ~pi141 & ~new_n346_;
  assign po25 = new_n345_ | ~new_n347_;
  assign new_n349_ = pi123 & ~pi124;
  assign new_n350_ = ~pi123 & pi124;
  assign new_n351_ = ~new_n349_ & ~new_n350_;
  assign new_n352_ = ~pi149 & ~pi150;
  assign new_n353_ = pi149 & pi150;
  assign new_n354_ = ~new_n352_ & ~new_n353_;
  assign new_n355_ = pi145 & new_n354_;
  assign new_n356_ = ~pi145 & ~new_n354_;
  assign new_n357_ = ~new_n355_ & ~new_n356_;
  assign new_n358_ = ~pi151 & ~pi152;
  assign new_n359_ = pi151 & pi152;
  assign new_n360_ = ~new_n358_ & ~new_n359_;
  assign new_n361_ = ~pi147 & ~pi148;
  assign new_n362_ = pi147 & pi148;
  assign new_n363_ = ~new_n361_ & ~new_n362_;
  assign new_n364_ = pi146 & new_n363_;
  assign new_n365_ = ~pi146 & ~new_n363_;
  assign new_n366_ = ~new_n364_ & ~new_n365_;
  assign new_n367_ = new_n360_ & ~new_n366_;
  assign new_n368_ = ~new_n360_ & new_n366_;
  assign new_n369_ = ~new_n367_ & ~new_n368_;
  assign new_n370_ = ~new_n357_ & new_n369_;
  assign new_n371_ = new_n357_ & ~new_n369_;
  assign new_n372_ = ~new_n370_ & ~new_n371_;
  assign new_n373_ = ~new_n351_ & ~new_n372_;
  assign new_n374_ = new_n351_ & new_n372_;
  assign new_n375_ = pi009 & ~new_n374_;
  assign po26 = ~new_n373_ & new_n375_;
  assign new_n377_ = pi140 & ~pi141;
  assign new_n378_ = ~pi140 & pi141;
  assign new_n379_ = ~new_n377_ & ~new_n378_;
  assign new_n380_ = ~pi138 & ~pi139;
  assign new_n381_ = ~new_n193_ & ~new_n380_;
  assign new_n382_ = ~pi136 & ~pi137;
  assign new_n383_ = ~new_n192_ & ~new_n382_;
  assign new_n384_ = pi135 & ~pi154;
  assign new_n385_ = ~pi135 & pi154;
  assign new_n386_ = ~new_n384_ & ~new_n385_;
  assign new_n387_ = new_n383_ & new_n386_;
  assign new_n388_ = ~new_n383_ & ~new_n386_;
  assign new_n389_ = ~new_n387_ & ~new_n388_;
  assign new_n390_ = new_n381_ & ~new_n389_;
  assign new_n391_ = ~new_n381_ & new_n389_;
  assign new_n392_ = ~new_n390_ & ~new_n391_;
  assign new_n393_ = new_n379_ & new_n392_;
  assign new_n394_ = ~new_n379_ & ~new_n392_;
  assign po27 = ~new_n393_ & ~new_n394_;
  assign new_n396_ = ~pi131 & ~pi132;
  assign new_n397_ = pi131 & pi132;
  assign new_n398_ = ~new_n396_ & ~new_n397_;
  assign new_n399_ = ~pi129 & ~pi130;
  assign new_n400_ = pi129 & pi130;
  assign new_n401_ = ~new_n399_ & ~new_n400_;
  assign new_n402_ = pi126 & new_n401_;
  assign new_n403_ = ~pi126 & ~new_n401_;
  assign new_n404_ = ~new_n402_ & ~new_n403_;
  assign new_n405_ = new_n398_ & ~new_n404_;
  assign new_n406_ = ~new_n398_ & new_n404_;
  assign new_n407_ = ~new_n405_ & ~new_n406_;
  assign new_n408_ = ~pi127 & ~pi128;
  assign new_n409_ = pi127 & pi128;
  assign new_n410_ = ~new_n408_ & ~new_n409_;
  assign new_n411_ = pi153 & new_n410_;
  assign new_n412_ = ~pi153 & ~new_n410_;
  assign new_n413_ = ~new_n411_ & ~new_n412_;
  assign new_n414_ = pi133 & ~pi134;
  assign new_n415_ = ~pi133 & pi134;
  assign new_n416_ = ~new_n414_ & ~new_n415_;
  assign new_n417_ = new_n413_ & ~new_n416_;
  assign new_n418_ = ~new_n413_ & new_n416_;
  assign new_n419_ = ~new_n417_ & ~new_n418_;
  assign new_n420_ = new_n407_ & new_n419_;
  assign new_n421_ = ~new_n407_ & ~new_n419_;
  assign po28 = ~new_n420_ & ~new_n421_;
  assign new_n423_ = ~pi019 & ~pi022;
  assign new_n424_ = pi091 & pi142;
  assign new_n425_ = pi101 & ~pi142;
  assign new_n426_ = pi143 & ~new_n425_;
  assign new_n427_ = ~new_n424_ & new_n426_;
  assign new_n428_ = pi081 & pi142;
  assign new_n429_ = pi111 & ~pi142;
  assign new_n430_ = ~pi143 & ~new_n429_;
  assign new_n431_ = ~new_n428_ & new_n430_;
  assign new_n432_ = ~new_n427_ & ~new_n431_;
  assign new_n433_ = pi022 & ~new_n432_;
  assign new_n434_ = ~new_n423_ & ~new_n433_;
  assign new_n435_ = pi135 & new_n434_;
  assign new_n436_ = ~pi022 & ~pi026;
  assign new_n437_ = pi022 & po09;
  assign new_n438_ = ~new_n436_ & ~new_n437_;
  assign new_n439_ = ~pi139 & ~new_n438_;
  assign new_n440_ = ~pi005 & ~pi011;
  assign new_n441_ = pi011 & ~po19;
  assign new_n442_ = ~new_n440_ & ~new_n441_;
  assign new_n443_ = pi131 & new_n442_;
  assign new_n444_ = ~new_n439_ & ~new_n443_;
  assign new_n445_ = ~new_n435_ & new_n444_;
  assign new_n446_ = pi139 & new_n438_;
  assign new_n447_ = ~pi003 & ~pi011;
  assign new_n448_ = pi011 & ~new_n324_;
  assign new_n449_ = ~new_n447_ & ~new_n448_;
  assign new_n450_ = pi124 & new_n449_;
  assign new_n451_ = ~new_n446_ & ~new_n450_;
  assign new_n452_ = ~pi011 & ~pi012;
  assign new_n453_ = pi011 & ~new_n246_;
  assign new_n454_ = ~new_n452_ & ~new_n453_;
  assign new_n455_ = ~pi123 & ~new_n454_;
  assign new_n456_ = ~pi022 & ~pi025;
  assign new_n457_ = pi022 & po08;
  assign new_n458_ = ~new_n456_ & ~new_n457_;
  assign new_n459_ = pi138 & new_n458_;
  assign new_n460_ = ~new_n455_ & ~new_n459_;
  assign new_n461_ = new_n451_ & new_n460_;
  assign new_n462_ = ~pi022 & ~pi024;
  assign new_n463_ = pi090 & pi142;
  assign new_n464_ = pi100 & ~pi142;
  assign new_n465_ = pi143 & ~new_n464_;
  assign new_n466_ = ~new_n463_ & new_n465_;
  assign new_n467_ = pi080 & pi142;
  assign new_n468_ = pi110 & ~pi142;
  assign new_n469_ = ~pi143 & ~new_n468_;
  assign new_n470_ = ~new_n467_ & new_n469_;
  assign new_n471_ = ~new_n466_ & ~new_n470_;
  assign new_n472_ = pi022 & ~new_n471_;
  assign new_n473_ = ~new_n462_ & ~new_n472_;
  assign new_n474_ = pi136 & new_n473_;
  assign new_n475_ = ~pi135 & ~new_n434_;
  assign new_n476_ = ~new_n474_ & ~new_n475_;
  assign new_n477_ = ~pi131 & ~new_n442_;
  assign new_n478_ = pi123 & new_n454_;
  assign new_n479_ = ~new_n477_ & ~new_n478_;
  assign new_n480_ = new_n476_ & new_n479_;
  assign new_n481_ = new_n461_ & new_n480_;
  assign new_n482_ = new_n445_ & new_n481_;
  assign new_n483_ = ~pi011 & ~pi016;
  assign new_n484_ = pi011 & ~po18;
  assign new_n485_ = ~new_n483_ & ~new_n484_;
  assign new_n486_ = pi130 & ~new_n485_;
  assign new_n487_ = ~pi130 & new_n485_;
  assign new_n488_ = ~new_n486_ & ~new_n487_;
  assign new_n489_ = ~pi020 & ~pi022;
  assign new_n490_ = pi022 & po10;
  assign new_n491_ = ~new_n489_ & ~new_n490_;
  assign new_n492_ = pi137 & ~new_n491_;
  assign new_n493_ = ~pi137 & new_n491_;
  assign new_n494_ = ~new_n492_ & ~new_n493_;
  assign new_n495_ = ~pi018 & ~pi022;
  assign new_n496_ = pi084 & pi142;
  assign new_n497_ = pi094 & ~pi142;
  assign new_n498_ = pi143 & ~new_n497_;
  assign new_n499_ = ~new_n496_ & new_n498_;
  assign new_n500_ = pi074 & pi142;
  assign new_n501_ = pi104 & ~pi142;
  assign new_n502_ = ~pi143 & ~new_n501_;
  assign new_n503_ = ~new_n500_ & new_n502_;
  assign new_n504_ = ~new_n499_ & ~new_n503_;
  assign new_n505_ = pi022 & ~new_n504_;
  assign new_n506_ = ~new_n495_ & ~new_n505_;
  assign new_n507_ = pi133 & ~new_n506_;
  assign new_n508_ = ~pi133 & new_n506_;
  assign new_n509_ = ~new_n507_ & ~new_n508_;
  assign new_n510_ = ~new_n494_ & ~new_n509_;
  assign new_n511_ = ~new_n488_ & new_n510_;
  assign new_n512_ = ~pi136 & ~new_n473_;
  assign new_n513_ = pi022 & ~new_n344_;
  assign new_n514_ = ~pi021 & ~pi022;
  assign new_n515_ = pi008 & ~new_n514_;
  assign new_n516_ = ~new_n513_ & new_n515_;
  assign new_n517_ = ~new_n512_ & new_n516_;
  assign new_n518_ = ~pi022 & ~pi023;
  assign new_n519_ = pi092 & pi142;
  assign new_n520_ = pi102 & ~pi142;
  assign new_n521_ = pi143 & ~new_n520_;
  assign new_n522_ = ~new_n519_ & new_n521_;
  assign new_n523_ = pi082 & pi142;
  assign new_n524_ = pi112 & ~pi142;
  assign new_n525_ = ~pi143 & ~new_n524_;
  assign new_n526_ = ~new_n523_ & new_n525_;
  assign new_n527_ = ~new_n522_ & ~new_n526_;
  assign new_n528_ = pi022 & ~new_n527_;
  assign new_n529_ = ~new_n518_ & ~new_n528_;
  assign new_n530_ = pi134 & new_n529_;
  assign new_n531_ = ~pi124 & ~new_n449_;
  assign new_n532_ = ~new_n530_ & ~new_n531_;
  assign new_n533_ = new_n517_ & new_n532_;
  assign new_n534_ = ~pi011 & ~pi015;
  assign new_n535_ = pi011 & ~po17;
  assign new_n536_ = ~new_n534_ & ~new_n535_;
  assign new_n537_ = pi129 & ~new_n536_;
  assign new_n538_ = ~pi129 & new_n536_;
  assign new_n539_ = ~new_n537_ & ~new_n538_;
  assign new_n540_ = ~pi004 & ~pi011;
  assign new_n541_ = pi011 & ~po15;
  assign new_n542_ = ~new_n540_ & ~new_n541_;
  assign new_n543_ = pi127 & ~new_n542_;
  assign new_n544_ = ~pi127 & new_n542_;
  assign new_n545_ = ~new_n543_ & ~new_n544_;
  assign new_n546_ = ~new_n539_ & ~new_n545_;
  assign new_n547_ = new_n533_ & new_n546_;
  assign new_n548_ = ~pi011 & ~pi017;
  assign new_n549_ = pi011 & ~po20;
  assign new_n550_ = ~new_n548_ & ~new_n549_;
  assign new_n551_ = pi132 & new_n550_;
  assign new_n552_ = ~pi134 & ~new_n529_;
  assign new_n553_ = ~new_n551_ & ~new_n552_;
  assign new_n554_ = ~pi138 & ~new_n458_;
  assign new_n555_ = ~pi011 & ~pi014;
  assign new_n556_ = pi011 & ~po16;
  assign new_n557_ = ~new_n555_ & ~new_n556_;
  assign new_n558_ = pi128 & new_n557_;
  assign new_n559_ = ~new_n554_ & ~new_n558_;
  assign new_n560_ = new_n553_ & new_n559_;
  assign new_n561_ = ~pi132 & ~new_n550_;
  assign new_n562_ = ~pi011 & ~pi013;
  assign new_n563_ = pi011 & ~po14;
  assign new_n564_ = ~new_n562_ & ~new_n563_;
  assign new_n565_ = pi126 & new_n564_;
  assign new_n566_ = ~new_n561_ & ~new_n565_;
  assign new_n567_ = ~pi128 & ~new_n557_;
  assign new_n568_ = ~pi126 & ~new_n564_;
  assign new_n569_ = ~new_n567_ & ~new_n568_;
  assign new_n570_ = new_n566_ & new_n569_;
  assign new_n571_ = new_n560_ & new_n570_;
  assign new_n572_ = new_n547_ & new_n571_;
  assign new_n573_ = new_n511_ & new_n572_;
  assign po29 = new_n482_ & new_n573_;
  assign new_n575_ = ~new_n324_ & new_n330_;
  assign new_n576_ = po11 & ~new_n575_;
  assign new_n577_ = pi061 & pi116;
  assign new_n578_ = pi050 & ~pi116;
  assign new_n579_ = pi119 & ~new_n578_;
  assign new_n580_ = ~new_n577_ & new_n579_;
  assign new_n581_ = pi040 & pi116;
  assign new_n582_ = pi072 & ~pi116;
  assign new_n583_ = ~pi119 & ~new_n582_;
  assign new_n584_ = ~new_n581_ & new_n583_;
  assign new_n585_ = ~new_n580_ & ~new_n584_;
  assign new_n586_ = ~new_n246_ & ~new_n585_;
  assign new_n587_ = new_n246_ & new_n585_;
  assign new_n588_ = ~new_n586_ & ~new_n587_;
  assign new_n589_ = ~new_n576_ & ~new_n588_;
  assign new_n590_ = new_n576_ & new_n588_;
  assign po30 = ~new_n589_ & ~new_n590_;
  assign new_n592_ = ~po08 & po09;
  assign new_n593_ = po08 & ~po09;
  assign new_n594_ = ~new_n592_ & ~new_n593_;
  assign new_n595_ = new_n344_ & new_n594_;
  assign new_n596_ = ~new_n344_ & ~new_n594_;
  assign new_n597_ = ~new_n595_ & ~new_n596_;
  assign new_n598_ = ~new_n432_ & new_n527_;
  assign new_n599_ = new_n432_ & ~new_n527_;
  assign new_n600_ = ~new_n598_ & ~new_n599_;
  assign new_n601_ = pi093 & pi142;
  assign new_n602_ = pi103 & ~pi142;
  assign new_n603_ = pi143 & ~new_n602_;
  assign new_n604_ = ~new_n601_ & new_n603_;
  assign new_n605_ = pi083 & pi142;
  assign new_n606_ = pi113 & ~pi142;
  assign new_n607_ = ~pi143 & ~new_n606_;
  assign new_n608_ = ~new_n605_ & new_n607_;
  assign new_n609_ = ~new_n604_ & ~new_n608_;
  assign new_n610_ = ~po10 & ~new_n504_;
  assign new_n611_ = po10 & new_n504_;
  assign new_n612_ = ~new_n610_ & ~new_n611_;
  assign new_n613_ = new_n471_ & new_n612_;
  assign new_n614_ = ~new_n471_ & ~new_n612_;
  assign new_n615_ = ~new_n613_ & ~new_n614_;
  assign new_n616_ = new_n609_ & ~new_n615_;
  assign new_n617_ = ~new_n609_ & new_n615_;
  assign new_n618_ = ~new_n616_ & ~new_n617_;
  assign new_n619_ = new_n600_ & new_n618_;
  assign new_n620_ = ~new_n600_ & ~new_n618_;
  assign new_n621_ = ~new_n619_ & ~new_n620_;
  assign new_n622_ = new_n597_ & new_n621_;
  assign new_n623_ = ~new_n597_ & ~new_n621_;
  assign new_n624_ = ~pi028 & ~new_n623_;
  assign po31 = ~new_n622_ & new_n624_;
  assign new_n626_ = po17 & ~po19;
  assign new_n627_ = ~po17 & po19;
  assign new_n628_ = ~new_n626_ & ~new_n627_;
  assign new_n629_ = ~po18 & po20;
  assign new_n630_ = po18 & ~po20;
  assign new_n631_ = ~new_n629_ & ~new_n630_;
  assign new_n632_ = new_n628_ & new_n631_;
  assign new_n633_ = ~new_n628_ & ~new_n631_;
  assign new_n634_ = ~new_n632_ & ~new_n633_;
  assign new_n635_ = ~po14 & ~new_n588_;
  assign new_n636_ = po14 & new_n588_;
  assign new_n637_ = ~new_n635_ & ~new_n636_;
  assign new_n638_ = new_n332_ & ~new_n637_;
  assign new_n639_ = new_n324_ & ~new_n637_;
  assign new_n640_ = ~new_n324_ & new_n637_;
  assign new_n641_ = ~new_n639_ & ~new_n640_;
  assign new_n642_ = ~new_n332_ & ~new_n641_;
  assign new_n643_ = ~new_n638_ & ~new_n642_;
  assign new_n644_ = new_n634_ & ~new_n643_;
  assign new_n645_ = ~new_n634_ & new_n643_;
  assign new_n646_ = ~new_n644_ & ~new_n645_;
  assign new_n647_ = pi122 & ~new_n646_;
  assign new_n648_ = ~pi122 & new_n585_;
  assign po32 = new_n647_ | new_n648_;
  assign new_n650_ = ~po15 & po16;
  assign new_n651_ = po15 & ~po16;
  assign new_n652_ = ~new_n650_ & ~new_n651_;
  assign new_n653_ = new_n641_ & new_n652_;
  assign new_n654_ = ~new_n641_ & ~new_n652_;
  assign new_n655_ = ~new_n653_ & ~new_n654_;
  assign new_n656_ = new_n634_ & ~new_n655_;
  assign new_n657_ = ~new_n634_ & new_n655_;
  assign new_n658_ = ~pi028 & ~new_n657_;
  assign po33 = ~new_n656_ & new_n658_;
  assign new_n660_ = ~pi125 & ~po10;
  assign new_n661_ = pi029 & po08;
  assign new_n662_ = new_n660_ & new_n661_;
  assign new_n663_ = pi128 & ~new_n662_;
  assign new_n664_ = pi138 & new_n662_;
  assign new_n665_ = pi007 & ~new_n664_;
  assign new_n666_ = ~new_n663_ & new_n665_;
  assign new_n667_ = ~po16 & new_n666_;
  assign new_n668_ = pi007 & po16;
  assign new_n669_ = ~new_n666_ & new_n668_;
  assign new_n670_ = ~new_n667_ & ~new_n669_;
  assign new_n671_ = pi129 & ~new_n662_;
  assign new_n672_ = pi139 & new_n662_;
  assign new_n673_ = pi007 & ~new_n672_;
  assign new_n674_ = ~new_n671_ & new_n673_;
  assign new_n675_ = pi007 & po17;
  assign new_n676_ = ~new_n674_ & new_n675_;
  assign new_n677_ = ~po17 & new_n674_;
  assign new_n678_ = ~new_n676_ & ~new_n677_;
  assign new_n679_ = pi127 & ~new_n662_;
  assign new_n680_ = pi137 & new_n662_;
  assign new_n681_ = ~new_n679_ & ~new_n680_;
  assign new_n682_ = ~po15 & new_n681_;
  assign new_n683_ = pi007 & ~pi131;
  assign new_n684_ = ~po19 & new_n683_;
  assign new_n685_ = ~new_n662_ & new_n684_;
  assign new_n686_ = pi007 & ~pi130;
  assign new_n687_ = pi007 & ~new_n686_;
  assign new_n688_ = po18 & new_n687_;
  assign new_n689_ = ~new_n662_ & new_n688_;
  assign new_n690_ = ~new_n685_ & ~new_n689_;
  assign new_n691_ = pi007 & ~new_n683_;
  assign new_n692_ = po19 & new_n691_;
  assign new_n693_ = ~new_n662_ & new_n692_;
  assign new_n694_ = ~po18 & new_n686_;
  assign new_n695_ = ~new_n662_ & new_n694_;
  assign new_n696_ = ~new_n693_ & ~new_n695_;
  assign new_n697_ = new_n690_ & new_n696_;
  assign new_n698_ = new_n682_ & new_n697_;
  assign new_n699_ = new_n678_ & new_n698_;
  assign new_n700_ = new_n670_ & new_n699_;
  assign new_n701_ = po15 & ~new_n681_;
  assign new_n702_ = ~new_n682_ & ~new_n701_;
  assign new_n703_ = pi126 & ~new_n662_;
  assign new_n704_ = pi136 & new_n662_;
  assign new_n705_ = ~new_n703_ & ~new_n704_;
  assign new_n706_ = po14 & ~new_n705_;
  assign new_n707_ = new_n697_ & ~new_n706_;
  assign new_n708_ = new_n702_ & new_n707_;
  assign new_n709_ = new_n678_ & new_n708_;
  assign new_n710_ = pi124 & ~new_n662_;
  assign new_n711_ = pi135 & new_n662_;
  assign new_n712_ = ~new_n710_ & ~new_n711_;
  assign new_n713_ = new_n324_ & ~new_n712_;
  assign new_n714_ = pi123 & ~new_n662_;
  assign new_n715_ = pi134 & new_n662_;
  assign new_n716_ = ~new_n246_ & ~new_n715_;
  assign new_n717_ = ~new_n714_ & new_n716_;
  assign new_n718_ = ~new_n713_ & new_n717_;
  assign new_n719_ = ~po14 & new_n705_;
  assign new_n720_ = ~new_n324_ & new_n712_;
  assign new_n721_ = ~new_n719_ & ~new_n720_;
  assign new_n722_ = ~new_n718_ & new_n721_;
  assign new_n723_ = new_n670_ & ~new_n722_;
  assign new_n724_ = new_n709_ & new_n723_;
  assign new_n725_ = new_n667_ & new_n697_;
  assign new_n726_ = new_n678_ & new_n725_;
  assign new_n727_ = new_n677_ & new_n697_;
  assign new_n728_ = ~new_n693_ & new_n695_;
  assign new_n729_ = ~new_n685_ & ~new_n728_;
  assign new_n730_ = ~new_n727_ & new_n729_;
  assign new_n731_ = ~new_n726_ & new_n730_;
  assign new_n732_ = ~new_n724_ & new_n731_;
  assign new_n733_ = ~new_n700_ & new_n732_;
  assign new_n734_ = ~new_n660_ & new_n661_;
  assign new_n735_ = pi135 & new_n432_;
  assign new_n736_ = new_n734_ & new_n735_;
  assign new_n737_ = ~pi134 & ~new_n527_;
  assign new_n738_ = new_n734_ & new_n737_;
  assign new_n739_ = ~new_n736_ & ~new_n738_;
  assign new_n740_ = pi132 & po20;
  assign new_n741_ = new_n734_ & new_n740_;
  assign new_n742_ = pi133 & new_n504_;
  assign new_n743_ = new_n734_ & new_n742_;
  assign new_n744_ = ~new_n741_ & ~new_n743_;
  assign new_n745_ = new_n739_ & new_n744_;
  assign new_n746_ = ~pi132 & ~po20;
  assign new_n747_ = new_n734_ & new_n746_;
  assign new_n748_ = ~pi133 & ~new_n504_;
  assign new_n749_ = new_n734_ & new_n748_;
  assign new_n750_ = ~new_n747_ & ~new_n749_;
  assign new_n751_ = ~pi135 & ~new_n432_;
  assign new_n752_ = new_n734_ & new_n751_;
  assign new_n753_ = pi134 & new_n527_;
  assign new_n754_ = new_n734_ & new_n753_;
  assign new_n755_ = ~new_n752_ & ~new_n754_;
  assign new_n756_ = new_n750_ & new_n755_;
  assign new_n757_ = new_n745_ & new_n756_;
  assign new_n758_ = ~new_n733_ & new_n757_;
  assign new_n759_ = new_n742_ & ~new_n749_;
  assign new_n760_ = ~new_n750_ & ~new_n754_;
  assign new_n761_ = ~new_n759_ & new_n760_;
  assign new_n762_ = ~new_n738_ & ~new_n761_;
  assign new_n763_ = ~new_n736_ & ~new_n762_;
  assign new_n764_ = ~new_n752_ & ~new_n763_;
  assign po34 = new_n758_ | ~new_n764_;
  assign new_n766_ = po07 & ~po27;
  assign new_n767_ = ~po28 & new_n766_;
  assign new_n768_ = ~po26 & new_n767_;
  assign new_n769_ = ~po31 & new_n768_;
  assign po35 = ~po33 & new_n769_;
endmodule


