// Benchmark "c2670" written by ABC on Thu Jul 14 21:14:08 2022

module c2670 ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
    G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
    G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
    G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
    G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
    G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
    G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136,
    G137, G138, G139, G140, G141, G142, _IN_G169 , _IN_G174 , _IN_G177 ,
    _IN_G178 , _IN_G179 , _IN_G180 , _IN_G181 , _IN_G182 , _IN_G183 ,
    _IN_G184 , _IN_G185 , _IN_G186 , _IN_G189 , _IN_G190 , _IN_G191 ,
    _IN_G192 , _IN_G193 , _IN_G194 , _IN_G195 , _IN_G196 , _IN_G197 ,
    _IN_G198 , _IN_G199 , _IN_G200 , _IN_G201 , _IN_G202 , _IN_G203 ,
    _IN_G204 , _IN_G205 , _IN_G206 , _IN_G207 , _IN_G208 , _IN_G209 ,
    _IN_G210 , _IN_G211 , _IN_G212 , _IN_G213 , _IN_G214 , _IN_G215 ,
    _IN_G239 , _IN_G240 , _IN_G241 , _IN_G242 , _IN_G243 , _IN_G244 ,
    _IN_G245 , _IN_G246 , _IN_G247 , _IN_G248 , _IN_G249 , _IN_G250 ,
    _IN_G251 , _IN_G252 , _IN_G253 , _IN_G254 , _IN_G255 , _IN_G256 ,
    _IN_G257 , _IN_G262 , _IN_G263 , _IN_G264 , _IN_G265 , _IN_G266 ,
    _IN_G267 , _IN_G268 , _IN_G269 , _IN_G270 , _IN_G271 , _IN_G272 ,
    _IN_G273 , _IN_G274 , _IN_G275 , _IN_G276 , _IN_G277 , _IN_G278 ,
    _IN_G279 , G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083,
    G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986,
    G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100,
    G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451,
    G2454, G2474, G2678,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    // G276, G277, G278, G279, G350, G335, G409, G369, G367, G411, G337, G384,
    G276, G277, G278, G279,
    // G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173,
    G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G173,
    G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171,
    // G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
    G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284,
    // G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145,
    G297, G148, G282, G156, G401, G227, G229, G311, G150, G145,
    // G395, G295, G331, G397, G329, G231, G308, G225  );
    G395, G295, G397, G329, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20,
    G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36,
    G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74,
    G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90,
    G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105,
    G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
    G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135,
    G136, G137, G138, G139, G140, G141, G142, _IN_G169 , _IN_G174 ,
    _IN_G177 , _IN_G178 , _IN_G179 , _IN_G180 , _IN_G181 , _IN_G182 ,
    _IN_G183 , _IN_G184 , _IN_G185 , _IN_G186 , _IN_G189 , _IN_G190 ,
    _IN_G191 , _IN_G192 , _IN_G193 , _IN_G194 , _IN_G195 , _IN_G196 ,
    _IN_G197 , _IN_G198 , _IN_G199 , _IN_G200 , _IN_G201 , _IN_G202 ,
    _IN_G203 , _IN_G204 , _IN_G205 , _IN_G206 , _IN_G207 , _IN_G208 ,
    _IN_G209 , _IN_G210 , _IN_G211 , _IN_G212 , _IN_G213 , _IN_G214 ,
    _IN_G215 , _IN_G239 , _IN_G240 , _IN_G241 , _IN_G242 , _IN_G243 ,
    _IN_G244 , _IN_G245 , _IN_G246 , _IN_G247 , _IN_G248 , _IN_G249 ,
    _IN_G250 , _IN_G251 , _IN_G252 , _IN_G253 , _IN_G254 , _IN_G255 ,
    _IN_G256 , _IN_G257 , _IN_G262 , _IN_G263 , _IN_G264 , _IN_G265 ,
    _IN_G266 , _IN_G267 , _IN_G268 , _IN_G269 , _IN_G270 , _IN_G271 ,
    _IN_G272 , _IN_G273 , _IN_G274 , _IN_G275 , _IN_G276 , _IN_G277 ,
    _IN_G278 , _IN_G279 , G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185,
    G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199,
    G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211,
    G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
    G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262,
    G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274,
    // G275, G276, G277, G278, G279, G350, G335, G409, G369, G367, G411, G337,
    G275, G276, G277, G278, G279, 
    // G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391,
    G218, G219, G220, G221, G235, G236, G237, G238, G158, G259,
    G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168,
    G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284,
    // G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
    G297, G148, G282, G156, G401, G227, G229, G311, G150,
    // G145, G395, G295, G331, G397, G329, G231, G308, G225;
    G145, G395, G295, G397, G329, G308, G225;
  wire new_new_n375__, new_new_n376__, new_new_n378__, new_new_n384__,
    new_new_n385__, new_new_n386__, new_new_n387__, new_new_n388__,
    new_new_n389__, new_new_n391__, new_new_n392__, new_new_n394__,
    new_new_n395__, new_new_n396__, new_new_n397__, new_new_n398__,
    new_new_n399__, new_new_n400__, new_new_n401__, new_new_n403__,
    new_new_n404__, new_new_n405__, new_new_n406__, new_new_n407__,
    new_new_n408__, new_new_n409__, new_new_n410__, new_new_n412__,
    new_new_n413__, new_new_n414__, new_new_n415__, new_new_n416__,
    new_new_n417__, new_new_n418__, new_new_n419__, new_new_n421__,
    new_new_n422__, new_new_n423__, new_new_n424__, new_new_n425__,
    new_new_n426__, new_new_n427__, new_new_n428__, new_new_n430__,
    new_new_n431__, new_new_n432__, new_new_n433__, new_new_n434__,
    new_new_n435__, new_new_n436__, new_new_n437__, new_new_n439__,
    new_new_n440__, new_new_n441__, new_new_n442__, new_new_n443__,
    new_new_n444__, new_new_n445__, new_new_n446__, new_new_n448__,
    new_new_n449__, new_new_n450__, new_new_n451__, new_new_n452__,
    new_new_n453__, new_new_n454__, new_new_n455__, new_new_n456__,
    new_new_n458__, new_new_n459__, new_new_n461__, new_new_n462__,
    new_new_n464__, new_new_n465__, new_new_n466__, new_new_n467__,
    new_new_n468__, new_new_n469__, new_new_n470__, new_new_n471__,
    new_new_n473__, new_new_n474__, new_new_n475__, new_new_n476__,
    new_new_n477__, new_new_n478__, new_new_n480__, new_new_n481__,
    new_new_n482__, new_new_n483__, new_new_n484__, new_new_n485__,
    new_new_n486__, new_new_n487__, new_new_n489__, new_new_n490__,
    new_new_n491__, new_new_n492__, new_new_n493__, new_new_n494__,
    new_new_n495__, new_new_n496__, new_new_n498__, new_new_n499__,
    new_new_n500__, new_new_n501__, new_new_n502__, new_new_n503__,
    new_new_n504__, new_new_n505__, new_new_n506__, new_new_n507__,
    new_new_n508__, new_new_n510__, new_new_n511__, new_new_n513__,
    new_new_n515__, new_new_n516__, new_new_n517__, new_new_n519__,
    new_new_n520__, new_new_n521__, new_new_n522__, new_new_n523__,
    new_new_n524__, new_new_n525__, new_new_n526__, new_new_n527__,
    new_new_n528__, new_new_n529__, new_new_n530__, new_new_n532__,
    new_new_n533__, new_new_n534__, new_new_n535__, new_new_n536__,
    new_new_n537__, new_new_n538__, new_new_n539__, new_new_n540__,
    new_new_n541__, new_new_n542__, new_new_n543__, new_new_n544__,
    new_new_n545__, new_new_n546__, new_new_n547__, new_new_n548__,
    new_new_n549__, new_new_n550__, new_new_n551__, new_new_n552__,
    new_new_n553__, new_new_n554__, new_new_n555__, new_new_n556__,
    new_new_n557__, new_new_n558__, new_new_n560__, new_new_n561__,
    new_new_n562__, new_new_n563__, new_new_n564__, new_new_n565__,
    new_new_n566__, new_new_n567__, new_new_n568__, new_new_n569__,
    new_new_n570__, new_new_n571__, new_new_n572__, new_new_n573__,
    new_new_n574__, new_new_n575__, new_new_n576__, new_new_n577__,
    new_new_n579__, new_new_n580__, new_new_n581__, new_new_n582__,
    new_new_n583__, new_new_n584__, new_new_n585__, new_new_n586__,
    new_new_n587__, new_new_n588__, new_new_n589__, new_new_n590__,
    new_new_n591__, new_new_n592__, new_new_n593__, new_new_n594__,
    new_new_n595__, new_new_n596__, new_new_n597__, new_new_n598__,
    new_new_n599__, new_new_n600__, new_new_n601__, new_new_n602__,
    new_new_n603__, new_new_n604__, new_new_n606__, new_new_n607__,
    new_new_n608__, new_new_n609__, new_new_n610__, new_new_n611__,
    new_new_n612__, new_new_n613__, new_new_n614__, new_new_n615__,
    new_new_n616__, new_new_n617__, new_new_n618__, new_new_n619__,
    new_new_n620__, new_new_n621__, new_new_n622__, new_new_n623__,
    new_new_n624__, new_new_n625__, new_new_n626__, new_new_n627__,
    new_new_n628__, new_new_n629__, new_new_n630__, new_new_n631__,
    new_new_n632__, new_new_n633__, new_new_n634__, new_new_n635__,
    new_new_n636__, new_new_n637__, new_new_n638__, new_new_n639__,
    new_new_n640__, new_new_n641__, new_new_n642__, new_new_n643__,
    new_new_n644__, new_new_n645__, new_new_n646__, new_new_n647__,
    new_new_n648__, new_new_n649__, new_new_n650__, new_new_n651__,
    new_new_n652__, new_new_n653__, new_new_n654__, new_new_n655__,
    new_new_n656__, new_new_n657__, new_new_n658__, new_new_n659__,
    new_new_n660__, new_new_n661__, new_new_n662__, new_new_n663__,
    new_new_n664__, new_new_n665__, new_new_n666__, new_new_n667__,
    new_new_n668__, new_new_n669__, new_new_n670__, new_new_n671__,
    new_new_n672__, new_new_n673__, new_new_n674__, new_new_n675__,
    new_new_n676__, new_new_n677__, new_new_n678__, new_new_n679__,
    new_new_n680__, new_new_n681__, new_new_n682__, new_new_n683__,
    new_new_n684__, new_new_n685__, new_new_n686__, new_new_n687__,
    new_new_n688__, new_new_n689__, new_new_n690__, new_new_n691__,
    new_new_n692__, new_new_n693__, new_new_n694__, new_new_n695__,
    new_new_n696__, new_new_n697__, new_new_n698__, new_new_n699__,
    new_new_n700__, new_new_n701__, new_new_n702__, new_new_n703__,
    new_new_n704__, new_new_n705__, new_new_n706__, new_new_n707__,
    new_new_n708__, new_new_n709__, new_new_n710__, new_new_n711__,
    new_new_n712__, new_new_n713__, new_new_n714__, new_new_n715__,
    new_new_n716__, new_new_n717__, new_new_n718__, new_new_n719__,
    new_new_n720__, new_new_n721__, new_new_n722__, new_new_n723__,
    new_new_n724__, new_new_n725__, new_new_n726__, new_new_n727__,
    new_new_n728__, new_new_n729__, new_new_n730__, new_new_n731__,
    new_new_n732__, new_new_n733__, new_new_n734__, new_new_n735__,
    new_new_n736__, new_new_n737__, new_new_n738__, new_new_n739__,
    new_new_n740__, new_new_n741__, new_new_n742__, new_new_n743__,
    new_new_n744__, new_new_n745__, new_new_n746__, new_new_n747__,
    new_new_n748__, new_new_n749__, new_new_n750__, new_new_n751__,
    new_new_n752__, new_new_n753__, new_new_n754__, new_new_n755__,
    new_new_n756__, new_new_n758__, new_new_n759__, new_new_n760__,
    new_new_n761__, new_new_n762__, new_new_n763__, new_new_n764__,
    new_new_n765__, new_new_n766__, new_new_n767__, new_new_n768__,
    new_new_n769__, new_new_n770__, new_new_n771__, new_new_n772__,
    new_new_n773__, new_new_n775__, new_new_n776__, new_new_n777__,
    new_new_n778__, new_new_n779__, new_new_n780__, new_new_n781__,
    new_new_n782__, new_new_n783__, new_new_n784__, new_new_n785__,
    new_new_n786__, new_new_n787__, new_new_n788__, new_new_n789__,
    new_new_n790__, new_new_n791__, new_new_n792__, new_new_n793__,
    new_new_n794__, new_new_n795__, new_new_n796__, new_new_n797__,
    new_new_n798__, new_new_n799__, new_new_n800__, new_new_n801__,
    new_new_n802__, new_new_n803__, new_new_n804__, new_new_n805__,
    new_new_n806__, new_new_n807__, new_new_n809__, new_new_n810__,
    new_new_n811__, new_new_n812__, new_new_n813__, new_new_n814__,
    new_new_n815__, new_new_n816__, new_new_n817__, new_new_n818__,
    new_new_n819__, new_new_n820__, new_new_n821__, new_new_n822__,
    new_new_n823__, new_new_n824__, new_new_n825__, new_new_n826__,
    new_new_n827__, new_new_n828__, new_new_n829__, new_new_n830__,
    new_new_n831__, new_new_n833__, new_new_n834__, new_new_n835__,
    new_new_n836__, new_new_n837__, new_new_n838__, new_new_n839__,
    new_new_n840__, new_new_n841__, new_new_n843__, new_new_n844__,
    new_new_n845__, new_new_n846__, new_new_n847__, new_new_n848__,
    new_new_n849__, new_new_n850__, new_new_n851__, new_new_n852__,
    new_new_n853__, new_new_n854__, new_new_n855__, new_new_n856__,
    new_new_n857__, new_new_n858__, new_new_n859__, new_new_n860__,
    new_new_n861__, new_new_n862__, new_new_n863__, new_new_n864__,
    new_new_n865__, new_new_n866__, new_new_n867__, new_new_n868__,
    new_new_n869__, new_new_n870__, new_new_n871__, new_new_n872__,
    new_new_n873__, new_new_n874__, new_new_n875__, new_new_n876__,
    new_new_n877__, new_new_n878__, new_new_n879__, new_new_n880__,
    new_new_n881__, new_new_n882__, new_new_n883__, new_new_n884__,
    new_new_n885__, new_new_n886__, new_new_n887__, new_new_n888__,
    new_new_n889__, new_new_n890__, new_new_n891__, new_new_n892__,
    new_new_n893__, new_new_n894__, new_new_n895__, new_new_n896__,
    new_new_n897__, new_new_n898__, new_new_n899__, new_new_n900__,
    new_new_n901__, new_new_n902__, new_new_n903__, new_new_n904__,
    new_new_n905__, new_new_n906__, new_new_n907__, new_new_n908__,
    new_new_n909__, new_new_n910__, new_new_n911__, new_new_n912__,
    new_new_n913__, new_new_n914__, new_new_n915__, new_new_n916__,
    new_new_n917__, new_new_n918__, new_new_n919__, new_new_n920__,
    new_new_n921__, new_new_n922__, new_new_n923__, new_new_n924__,
    new_new_n925__, new_new_n926__, new_new_n927__, new_new_n928__,
    new_new_n929__, new_new_n930__, new_new_n931__, new_new_n932__,
    new_new_n933__, new_new_n934__, new_new_n935__, new_new_n936__,
    new_new_n937__, new_new_n938__, new_new_n939__, new_new_n940__,
    new_new_n941__, new_new_n942__, new_new_n943__, new_new_n944__,
    new_new_n945__, new_new_n946__, new_new_n947__, new_new_n949__,
    new_new_n950__, new_new_n951__, new_new_n952__;
  assign new_new_n375__ = G2072 & G2078;
  assign new_new_n376__ = G2084 & G2090;
  assign G158 = ~new_new_n375__ | ~new_new_n376__;
  assign new_new_n378__ = G2 & G15;
  assign G259 = ~G661 | ~new_new_n378__;
  assign G173 = G94 & G452;
  assign G223 = ~G7 | ~G661;
  assign G234 = ~G567 | G223;
  assign G217 = ~G2106 | G223;
  assign new_new_n384__ = G57 & G69;
  assign new_new_n385__ = G108 & G120;
  assign new_new_n386__ = new_new_n384__ & new_new_n385__;
  assign new_new_n387__ = G44 & G82;
  assign new_new_n388__ = G96 & G132;
  assign new_new_n389__ = new_new_n387__ & new_new_n388__;
  assign G325 = new_new_n386__ & new_new_n389__;
  assign new_new_n391__ = G2106 & ~new_new_n389__;
  assign new_new_n392__ = G567 & ~new_new_n386__;
  assign G319 = ~new_new_n391__ & ~new_new_n392__;
  assign new_new_n394__ = G125 & ~G2104;
  assign new_new_n395__ = G113 & G2104;
  assign new_new_n396__ = G2105 & ~new_new_n394__;
  assign new_new_n397__ = ~new_new_n395__ & new_new_n396__;
  assign new_new_n398__ = G137 & ~G2104;
  assign new_new_n399__ = G101 & G2104;
  assign new_new_n400__ = ~G2105 & ~new_new_n398__;
  assign new_new_n401__ = ~new_new_n399__ & new_new_n400__;
  assign G160 = new_new_n397__ | new_new_n401__;
  assign new_new_n403__ = G124 & ~G2104;
  assign new_new_n404__ = G112 & G2104;
  assign new_new_n405__ = G2105 & ~new_new_n403__;
  assign new_new_n406__ = ~new_new_n404__ & new_new_n405__;
  assign new_new_n407__ = G136 & ~G2104;
  assign new_new_n408__ = G100 & G2104;
  assign new_new_n409__ = ~G2105 & ~new_new_n407__;
  assign new_new_n410__ = ~new_new_n408__ & new_new_n409__;
  assign G162 = new_new_n406__ | new_new_n410__;
  assign new_new_n412__ = G126 & ~G2104;
  assign new_new_n413__ = G114 & G2104;
  assign new_new_n414__ = G2105 & ~new_new_n412__;
  assign new_new_n415__ = ~new_new_n413__ & new_new_n414__;
  assign new_new_n416__ = G138 & ~G2104;
  assign new_new_n417__ = G102 & G2104;
  assign new_new_n418__ = ~G2105 & ~new_new_n416__;
  assign new_new_n419__ = ~new_new_n417__ & new_new_n418__;
  assign G164 = new_new_n415__ | new_new_n419__;
  assign new_new_n421__ = G62 & ~G543;
  assign new_new_n422__ = G75 & G543;
  assign new_new_n423__ = G651 & ~new_new_n421__;
  assign new_new_n424__ = ~new_new_n422__ & new_new_n423__;
  assign new_new_n425__ = G88 & ~G543;
  assign new_new_n426__ = G50 & G543;
  assign new_new_n427__ = ~G651 & ~new_new_n425__;
  assign new_new_n428__ = ~new_new_n426__ & new_new_n427__;
  assign G303 = ~new_new_n424__ & ~new_new_n428__;
  assign new_new_n430__ = G63 & ~G543;
  assign new_new_n431__ = G76 & G543;
  assign new_new_n432__ = G651 & ~new_new_n430__;
  assign new_new_n433__ = ~new_new_n431__ & new_new_n432__;
  assign new_new_n434__ = G89 & ~G543;
  assign new_new_n435__ = G51 & G543;
  assign new_new_n436__ = ~G651 & ~new_new_n434__;
  assign new_new_n437__ = ~new_new_n435__ & new_new_n436__;
  assign G286 = ~new_new_n433__ & ~new_new_n437__;
  assign new_new_n439__ = G64 & ~G543;
  assign new_new_n440__ = G77 & G543;
  assign new_new_n441__ = G651 & ~new_new_n439__;
  assign new_new_n442__ = ~new_new_n440__ & new_new_n441__;
  assign new_new_n443__ = G90 & ~G543;
  assign new_new_n444__ = G52 & G543;
  assign new_new_n445__ = ~G651 & ~new_new_n443__;
  assign new_new_n446__ = ~new_new_n444__ & new_new_n445__;
  assign G301 = ~new_new_n442__ & ~new_new_n446__;
  assign new_new_n448__ = G56 & ~G543;
  assign new_new_n449__ = G68 & G543;
  assign new_new_n450__ = G651 & ~new_new_n448__;
  assign new_new_n451__ = ~new_new_n449__ & new_new_n450__;
  assign new_new_n452__ = G81 & ~G543;
  assign new_new_n453__ = G43 & G543;
  assign new_new_n454__ = ~G651 & ~new_new_n452__;
  assign new_new_n455__ = ~new_new_n453__ & new_new_n454__;
  assign new_new_n456__ = ~new_new_n451__ & ~new_new_n455__;
  assign G153 = ~G860 | new_new_n456__;
  assign new_new_n458__ = G483 & G661;
  assign new_new_n459__ = G36 & new_new_n458__;
  assign G176 = ~G319 | ~new_new_n459__;
  assign new_new_n461__ = G1 & G3;
  assign new_new_n462__ = new_new_n458__ & ~new_new_n461__;
  assign G188 = ~G319 | ~new_new_n462__;
  assign new_new_n464__ = G65 & ~G543;
  assign new_new_n465__ = G78 & G543;
  assign new_new_n466__ = G651 & ~new_new_n464__;
  assign new_new_n467__ = ~new_new_n465__ & new_new_n466__;
  assign new_new_n468__ = G91 & ~G543;
  assign new_new_n469__ = G53 & G543;
  assign new_new_n470__ = ~G651 & ~new_new_n468__;
  assign new_new_n471__ = ~new_new_n469__ & new_new_n470__;
  assign G299 = ~new_new_n467__ & ~new_new_n471__;
  assign new_new_n473__ = G49 & ~G651;
  assign new_new_n474__ = G74 & G651;
  assign new_new_n475__ = G543 & ~new_new_n473__;
  assign new_new_n476__ = ~new_new_n474__ & new_new_n475__;
  assign new_new_n477__ = ~G87 & ~G543;
  assign new_new_n478__ = ~G651 & new_new_n477__;
  assign G288 = ~new_new_n476__ & ~new_new_n478__;
  assign new_new_n480__ = G61 & ~G543;
  assign new_new_n481__ = G73 & G543;
  assign new_new_n482__ = G651 & ~new_new_n480__;
  assign new_new_n483__ = ~new_new_n481__ & new_new_n482__;
  assign new_new_n484__ = G86 & ~G543;
  assign new_new_n485__ = G48 & G543;
  assign new_new_n486__ = ~G651 & ~new_new_n484__;
  assign new_new_n487__ = ~new_new_n485__ & new_new_n486__;
  assign G305 = ~new_new_n483__ & ~new_new_n487__;
  assign new_new_n489__ = G60 & ~G543;
  assign new_new_n490__ = G72 & G543;
  assign new_new_n491__ = G651 & ~new_new_n489__;
  assign new_new_n492__ = ~new_new_n490__ & new_new_n491__;
  assign new_new_n493__ = G85 & ~G543;
  assign new_new_n494__ = G47 & G543;
  assign new_new_n495__ = ~G651 & ~new_new_n493__;
  assign new_new_n496__ = ~new_new_n494__ & new_new_n495__;
  assign G290 = ~new_new_n492__ & ~new_new_n496__;
  assign new_new_n498__ = G868 & ~G301;
  assign new_new_n499__ = G66 & ~G543;
  assign new_new_n500__ = G79 & G543;
  assign new_new_n501__ = G651 & ~new_new_n499__;
  assign new_new_n502__ = ~new_new_n500__ & new_new_n501__;
  assign new_new_n503__ = G92 & ~G543;
  assign new_new_n504__ = G54 & G543;
  assign new_new_n505__ = ~G651 & ~new_new_n503__;
  assign new_new_n506__ = ~new_new_n504__ & new_new_n505__;
  assign new_new_n507__ = ~new_new_n502__ & ~new_new_n506__;
  assign new_new_n508__ = ~G868 & ~new_new_n507__;
  assign G284 = ~new_new_n498__ & ~new_new_n508__;
  assign new_new_n510__ = G868 & ~G286;
  assign new_new_n511__ = ~G868 & ~G299;
  assign G297 = ~new_new_n510__ & ~new_new_n511__;
  assign new_new_n513__ = G559 & ~G860;
  assign G148 = new_new_n507__ | new_new_n513__;
  assign new_new_n515__ = ~G559 & ~new_new_n507__;
  assign new_new_n516__ = G868 & ~new_new_n515__;
  assign new_new_n517__ = ~G868 & new_new_n456__;
  assign G282 = new_new_n516__ | new_new_n517__;
  assign new_new_n519__ = G123 & ~G2104;
  assign new_new_n520__ = G111 & G2104;
  assign new_new_n521__ = G2105 & ~new_new_n519__;
  assign new_new_n522__ = ~new_new_n520__ & new_new_n521__;
  assign new_new_n523__ = G135 & ~G2104;
  assign new_new_n524__ = G99 & G2104;
  assign new_new_n525__ = ~G2105 & ~new_new_n523__;
  assign new_new_n526__ = ~new_new_n524__ & new_new_n525__;
  assign new_new_n527__ = ~new_new_n522__ & ~new_new_n526__;
  assign new_new_n528__ = ~G2096 & ~new_new_n527__;
  assign new_new_n529__ = G2096 & new_new_n527__;
  assign new_new_n530__ = ~G2100 & ~new_new_n528__;
  assign G156 = new_new_n529__ | ~new_new_n530__;
  assign new_new_n532__ = G1341 & ~G1348;
  assign new_new_n533__ = ~G1341 & G1348;
  assign new_new_n534__ = ~new_new_n532__ & ~new_new_n533__;
  assign new_new_n535__ = ~G2443 & ~G2446;
  assign new_new_n536__ = G2443 & G2446;
  assign new_new_n537__ = ~new_new_n535__ & ~new_new_n536__;
  assign new_new_n538__ = G2427 & new_new_n537__;
  assign new_new_n539__ = ~G2427 & ~new_new_n537__;
  assign new_new_n540__ = ~new_new_n538__ & ~new_new_n539__;
  assign new_new_n541__ = ~G2451 & ~G2454;
  assign new_new_n542__ = G2451 & G2454;
  assign new_new_n543__ = ~new_new_n541__ & ~new_new_n542__;
  assign new_new_n544__ = ~G2435 & ~G2438;
  assign new_new_n545__ = G2435 & G2438;
  assign new_new_n546__ = ~new_new_n544__ & ~new_new_n545__;
  assign new_new_n547__ = G2430 & new_new_n546__;
  assign new_new_n548__ = ~G2430 & ~new_new_n546__;
  assign new_new_n549__ = ~new_new_n547__ & ~new_new_n548__;
  assign new_new_n550__ = new_new_n543__ & ~new_new_n549__;
  assign new_new_n551__ = ~new_new_n543__ & new_new_n549__;
  assign new_new_n552__ = ~new_new_n550__ & ~new_new_n551__;
  assign new_new_n553__ = ~new_new_n540__ & new_new_n552__;
  assign new_new_n554__ = new_new_n540__ & ~new_new_n552__;
  assign new_new_n555__ = ~new_new_n553__ & ~new_new_n554__;
  assign new_new_n556__ = new_new_n534__ & new_new_n555__;
  assign new_new_n557__ = ~new_new_n534__ & ~new_new_n555__;
  assign new_new_n558__ = G14 & ~new_new_n556__;
  assign G401 = ~new_new_n557__ & new_new_n558__;
  assign new_new_n560__ = G2096 & ~G2100;
  assign new_new_n561__ = ~G2096 & G2100;
  assign new_new_n562__ = ~new_new_n560__ & ~new_new_n561__;
  assign new_new_n563__ = ~G2084 & ~G2090;
  assign new_new_n564__ = ~new_new_n376__ & ~new_new_n563__;
  assign new_new_n565__ = ~G2072 & ~G2078;
  assign new_new_n566__ = ~new_new_n375__ & ~new_new_n565__;
  assign new_new_n567__ = G2067 & ~G2678;
  assign new_new_n568__ = ~G2067 & G2678;
  assign new_new_n569__ = ~new_new_n567__ & ~new_new_n568__;
  assign new_new_n570__ = new_new_n566__ & new_new_n569__;
  assign new_new_n571__ = ~new_new_n566__ & ~new_new_n569__;
  assign new_new_n572__ = ~new_new_n570__ & ~new_new_n571__;
  assign new_new_n573__ = new_new_n564__ & ~new_new_n572__;
  assign new_new_n574__ = ~new_new_n564__ & new_new_n572__;
  assign new_new_n575__ = ~new_new_n573__ & ~new_new_n574__;
  assign new_new_n576__ = new_new_n562__ & new_new_n575__;
  assign new_new_n577__ = ~new_new_n562__ & ~new_new_n575__;
  assign G227 = ~new_new_n576__ & ~new_new_n577__;
  assign new_new_n579__ = ~G1981 & ~G1986;
  assign new_new_n580__ = G1981 & G1986;
  assign new_new_n581__ = ~new_new_n579__ & ~new_new_n580__;
  assign new_new_n582__ = ~G1971 & ~G1976;
  assign new_new_n583__ = G1971 & G1976;
  assign new_new_n584__ = ~new_new_n582__ & ~new_new_n583__;
  assign new_new_n585__ = G1956 & new_new_n584__;
  assign new_new_n586__ = ~G1956 & ~new_new_n584__;
  assign new_new_n587__ = ~new_new_n585__ & ~new_new_n586__;
  assign new_new_n588__ = new_new_n581__ & ~new_new_n587__;
  assign new_new_n589__ = ~new_new_n581__ & new_new_n587__;
  assign new_new_n590__ = ~new_new_n588__ & ~new_new_n589__;
  assign new_new_n591__ = ~G1961 & ~G1966;
  assign new_new_n592__ = G1961 & G1966;
  assign new_new_n593__ = ~new_new_n591__ & ~new_new_n592__;
  assign new_new_n594__ = G2474 & new_new_n593__;
  assign new_new_n595__ = ~G2474 & ~new_new_n593__;
  assign new_new_n596__ = ~new_new_n594__ & ~new_new_n595__;
  assign new_new_n597__ = G1991 & ~G1996;
  assign new_new_n598__ = ~G1991 & G1996;
  assign new_new_n599__ = ~new_new_n597__ & ~new_new_n598__;
  assign new_new_n600__ = new_new_n596__ & ~new_new_n599__;
  assign new_new_n601__ = ~new_new_n596__ & new_new_n599__;
  assign new_new_n602__ = ~new_new_n600__ & ~new_new_n601__;
  assign new_new_n603__ = new_new_n590__ & new_new_n602__;
  assign new_new_n604__ = ~new_new_n590__ & ~new_new_n602__;
  assign G229 = ~new_new_n603__ & ~new_new_n604__;
  assign new_new_n606__ = ~G29 & ~G33;
  assign new_new_n607__ = G127 & ~G2104;
  assign new_new_n608__ = G115 & G2104;
  assign new_new_n609__ = G2105 & ~new_new_n607__;
  assign new_new_n610__ = ~new_new_n608__ & new_new_n609__;
  assign new_new_n611__ = G139 & ~G2104;
  assign new_new_n612__ = G103 & G2104;
  assign new_new_n613__ = ~G2105 & ~new_new_n611__;
  assign new_new_n614__ = ~new_new_n612__ & new_new_n613__;
  assign new_new_n615__ = ~new_new_n610__ & ~new_new_n614__;
  assign new_new_n616__ = G29 & ~new_new_n615__;
  assign new_new_n617__ = ~new_new_n606__ & ~new_new_n616__;
  assign new_new_n618__ = ~G2072 & ~new_new_n617__;
  assign new_new_n619__ = ~G29 & ~G32;
  assign new_new_n620__ = G129 & ~G2104;
  assign new_new_n621__ = G117 & G2104;
  assign new_new_n622__ = G2105 & ~new_new_n620__;
  assign new_new_n623__ = ~new_new_n621__ & new_new_n622__;
  assign new_new_n624__ = G141 & ~G2104;
  assign new_new_n625__ = G105 & G2104;
  assign new_new_n626__ = ~G2105 & ~new_new_n624__;
  assign new_new_n627__ = ~new_new_n625__ & new_new_n626__;
  assign new_new_n628__ = ~new_new_n623__ & ~new_new_n627__;
  assign new_new_n629__ = G29 & ~new_new_n628__;
  assign new_new_n630__ = ~new_new_n619__ & ~new_new_n629__;
  assign new_new_n631__ = G1996 & new_new_n630__;
  assign new_new_n632__ = G29 & ~new_new_n527__;
  assign new_new_n633__ = ~G4 & ~G16;
  assign new_new_n634__ = G16 & ~new_new_n507__;
  assign new_new_n635__ = ~new_new_n633__ & ~new_new_n634__;
  assign new_new_n636__ = ~G1348 & ~new_new_n635__;
  assign new_new_n637__ = ~G16 & ~G24;
  assign new_new_n638__ = G16 & ~G290;
  assign new_new_n639__ = ~new_new_n637__ & ~new_new_n638__;
  assign new_new_n640__ = ~G1986 & ~new_new_n639__;
  assign new_new_n641__ = ~G16 & ~G20;
  assign new_new_n642__ = G16 & ~G299;
  assign new_new_n643__ = ~new_new_n641__ & ~new_new_n642__;
  assign new_new_n644__ = G1956 & new_new_n643__;
  assign new_new_n645__ = ~G16 & ~G22;
  assign new_new_n646__ = G16 & ~G303;
  assign new_new_n647__ = ~new_new_n645__ & ~new_new_n646__;
  assign new_new_n648__ = G1971 & ~new_new_n647__;
  assign new_new_n649__ = ~G1971 & new_new_n647__;
  assign new_new_n650__ = ~new_new_n648__ & ~new_new_n649__;
  assign new_new_n651__ = ~G16 & ~G21;
  assign new_new_n652__ = G16 & ~G286;
  assign new_new_n653__ = ~new_new_n651__ & ~new_new_n652__;
  assign new_new_n654__ = ~G1966 & ~new_new_n653__;
  assign new_new_n655__ = ~G1956 & ~new_new_n643__;
  assign new_new_n656__ = ~G28 & ~G29;
  assign new_new_n657__ = G1986 & new_new_n639__;
  assign new_new_n658__ = ~G1996 & ~new_new_n630__;
  assign new_new_n659__ = ~G29 & ~G34;
  assign new_new_n660__ = G29 & G160;
  assign new_new_n661__ = ~new_new_n659__ & ~new_new_n660__;
  assign new_new_n662__ = ~G2084 & ~new_new_n661__;
  assign new_new_n663__ = G1966 & new_new_n653__;
  assign new_new_n664__ = G2072 & new_new_n617__;
  assign new_new_n665__ = ~G5 & ~G16;
  assign new_new_n666__ = G16 & ~G301;
  assign new_new_n667__ = ~new_new_n665__ & ~new_new_n666__;
  assign new_new_n668__ = G1961 & ~new_new_n667__;
  assign new_new_n669__ = ~G1961 & new_new_n667__;
  assign new_new_n670__ = ~new_new_n668__ & ~new_new_n669__;
  assign new_new_n671__ = ~G26 & ~G29;
  assign new_new_n672__ = G128 & ~G2104;
  assign new_new_n673__ = G116 & G2104;
  assign new_new_n674__ = G2105 & ~new_new_n672__;
  assign new_new_n675__ = ~new_new_n673__ & new_new_n674__;
  assign new_new_n676__ = G140 & ~G2104;
  assign new_new_n677__ = G104 & G2104;
  assign new_new_n678__ = ~G2105 & ~new_new_n676__;
  assign new_new_n679__ = ~new_new_n677__ & new_new_n678__;
  assign new_new_n680__ = ~new_new_n675__ & ~new_new_n679__;
  assign new_new_n681__ = G29 & ~new_new_n680__;
  assign new_new_n682__ = ~new_new_n671__ & ~new_new_n681__;
  assign new_new_n683__ = ~G2067 & ~new_new_n682__;
  assign new_new_n684__ = ~G27 & ~G29;
  assign new_new_n685__ = G29 & G164;
  assign new_new_n686__ = ~new_new_n684__ & ~new_new_n685__;
  assign new_new_n687__ = G2078 & ~new_new_n686__;
  assign new_new_n688__ = ~G2078 & new_new_n686__;
  assign new_new_n689__ = ~new_new_n687__ & ~new_new_n688__;
  assign new_new_n690__ = ~G6 & ~G16;
  assign new_new_n691__ = G16 & ~G305;
  assign new_new_n692__ = ~new_new_n690__ & ~new_new_n691__;
  assign new_new_n693__ = ~G1981 & ~new_new_n692__;
  assign new_new_n694__ = ~G16 & ~G19;
  assign new_new_n695__ = G16 & ~new_new_n456__;
  assign new_new_n696__ = ~new_new_n694__ & ~new_new_n695__;
  assign new_new_n697__ = G1341 & new_new_n696__;
  assign new_new_n698__ = ~G29 & ~G35;
  assign new_new_n699__ = G29 & G162;
  assign new_new_n700__ = ~new_new_n698__ & ~new_new_n699__;
  assign new_new_n701__ = G2090 & new_new_n700__;
  assign new_new_n702__ = ~G25 & ~G29;
  assign new_new_n703__ = G119 & ~G2104;
  assign new_new_n704__ = G107 & G2104;
  assign new_new_n705__ = G2105 & ~new_new_n703__;
  assign new_new_n706__ = ~new_new_n704__ & new_new_n705__;
  assign new_new_n707__ = G131 & ~G2104;
  assign new_new_n708__ = G95 & G2104;
  assign new_new_n709__ = ~G2105 & ~new_new_n707__;
  assign new_new_n710__ = ~new_new_n708__ & new_new_n709__;
  assign new_new_n711__ = ~new_new_n706__ & ~new_new_n710__;
  assign new_new_n712__ = G29 & ~new_new_n711__;
  assign new_new_n713__ = ~new_new_n702__ & ~new_new_n712__;
  assign new_new_n714__ = G1991 & ~new_new_n713__;
  assign new_new_n715__ = ~G1991 & new_new_n713__;
  assign new_new_n716__ = ~new_new_n714__ & ~new_new_n715__;
  assign new_new_n717__ = G1348 & new_new_n635__;
  assign new_new_n718__ = ~G1341 & ~new_new_n696__;
  assign new_new_n719__ = G2084 & new_new_n661__;
  assign new_new_n720__ = ~G2090 & ~new_new_n700__;
  assign new_new_n721__ = G1981 & new_new_n692__;
  assign new_new_n722__ = G2067 & new_new_n682__;
  assign new_new_n723__ = ~G16 & ~G23;
  assign new_new_n724__ = G16 & ~G288;
  assign new_new_n725__ = ~new_new_n723__ & ~new_new_n724__;
  assign new_new_n726__ = G1976 & ~new_new_n725__;
  assign new_new_n727__ = ~G1976 & new_new_n725__;
  assign new_new_n728__ = ~new_new_n726__ & ~new_new_n727__;
  assign new_new_n729__ = G11 & ~new_new_n656__;
  assign new_new_n730__ = ~new_new_n632__ & new_new_n729__;
  assign new_new_n731__ = ~new_new_n618__ & new_new_n730__;
  assign new_new_n732__ = ~new_new_n631__ & ~new_new_n636__;
  assign new_new_n733__ = ~new_new_n640__ & ~new_new_n644__;
  assign new_new_n734__ = ~new_new_n654__ & ~new_new_n655__;
  assign new_new_n735__ = ~new_new_n657__ & ~new_new_n658__;
  assign new_new_n736__ = ~new_new_n662__ & ~new_new_n663__;
  assign new_new_n737__ = ~new_new_n664__ & ~new_new_n683__;
  assign new_new_n738__ = ~new_new_n693__ & ~new_new_n697__;
  assign new_new_n739__ = ~new_new_n701__ & ~new_new_n717__;
  assign new_new_n740__ = ~new_new_n718__ & ~new_new_n719__;
  assign new_new_n741__ = ~new_new_n720__ & ~new_new_n721__;
  assign new_new_n742__ = ~new_new_n722__ & new_new_n741__;
  assign new_new_n743__ = new_new_n739__ & new_new_n740__;
  assign new_new_n744__ = new_new_n737__ & new_new_n738__;
  assign new_new_n745__ = new_new_n735__ & new_new_n736__;
  assign new_new_n746__ = new_new_n733__ & new_new_n734__;
  assign new_new_n747__ = new_new_n731__ & new_new_n732__;
  assign new_new_n748__ = ~new_new_n650__ & ~new_new_n670__;
  assign new_new_n749__ = ~new_new_n689__ & ~new_new_n716__;
  assign new_new_n750__ = ~new_new_n728__ & new_new_n749__;
  assign new_new_n751__ = new_new_n747__ & new_new_n748__;
  assign new_new_n752__ = new_new_n745__ & new_new_n746__;
  assign new_new_n753__ = new_new_n743__ & new_new_n744__;
  assign new_new_n754__ = new_new_n742__ & new_new_n753__;
  assign new_new_n755__ = new_new_n751__ & new_new_n752__;
  assign new_new_n756__ = new_new_n750__ & new_new_n755__;
  assign G311 = new_new_n754__ & new_new_n756__;
  assign new_new_n758__ = ~new_new_n507__ & new_new_n513__;
  assign new_new_n759__ = G153 & ~new_new_n758__;
  assign new_new_n760__ = G67 & ~G543;
  assign new_new_n761__ = G80 & G543;
  assign new_new_n762__ = G651 & ~new_new_n760__;
  assign new_new_n763__ = ~new_new_n761__ & new_new_n762__;
  assign new_new_n764__ = G93 & ~G543;
  assign new_new_n765__ = G55 & G543;
  assign new_new_n766__ = ~G651 & ~new_new_n764__;
  assign new_new_n767__ = ~new_new_n765__ & new_new_n766__;
  assign new_new_n768__ = ~new_new_n763__ & ~new_new_n767__;
  assign new_new_n769__ = ~new_new_n456__ & ~new_new_n768__;
  assign new_new_n770__ = new_new_n456__ & new_new_n768__;
  assign new_new_n771__ = ~new_new_n769__ & ~new_new_n770__;
  assign new_new_n772__ = ~new_new_n759__ & ~new_new_n771__;
  assign new_new_n773__ = new_new_n759__ & new_new_n771__;
  assign G145 = ~new_new_n772__ & ~new_new_n773__;
  assign new_new_n775__ = ~G160 & G162;
  assign new_new_n776__ = G160 & ~G162;
  assign new_new_n777__ = ~new_new_n775__ & ~new_new_n776__;
  assign new_new_n778__ = new_new_n527__ & new_new_n777__;
  assign new_new_n779__ = ~new_new_n527__ & ~new_new_n777__;
  assign new_new_n780__ = ~new_new_n778__ & ~new_new_n779__;
  assign new_new_n781__ = new_new_n628__ & ~new_new_n680__;
  assign new_new_n782__ = ~new_new_n628__ & new_new_n680__;
  assign new_new_n783__ = ~new_new_n781__ & ~new_new_n782__;
  assign new_new_n784__ = G130 & ~G2104;
  assign new_new_n785__ = G118 & G2104;
  assign new_new_n786__ = G2105 & ~new_new_n784__;
  assign new_new_n787__ = ~new_new_n785__ & new_new_n786__;
  assign new_new_n788__ = G142 & ~G2104;
  assign new_new_n789__ = G106 & G2104;
  assign new_new_n790__ = ~G2105 & ~new_new_n788__;
  assign new_new_n791__ = ~new_new_n789__ & new_new_n790__;
  assign new_new_n792__ = ~new_new_n787__ & ~new_new_n791__;
  assign new_new_n793__ = ~G164 & ~new_new_n711__;
  assign new_new_n794__ = G164 & new_new_n711__;
  assign new_new_n795__ = ~new_new_n793__ & ~new_new_n794__;
  assign new_new_n796__ = new_new_n615__ & new_new_n795__;
  assign new_new_n797__ = ~new_new_n615__ & ~new_new_n795__;
  assign new_new_n798__ = ~new_new_n796__ & ~new_new_n797__;
  assign new_new_n799__ = new_new_n792__ & ~new_new_n798__;
  assign new_new_n800__ = ~new_new_n792__ & new_new_n798__;
  assign new_new_n801__ = ~new_new_n799__ & ~new_new_n800__;
  assign new_new_n802__ = new_new_n783__ & new_new_n801__;
  assign new_new_n803__ = ~new_new_n783__ & ~new_new_n801__;
  assign new_new_n804__ = ~new_new_n802__ & ~new_new_n803__;
  assign new_new_n805__ = ~new_new_n780__ & ~new_new_n804__;
  assign new_new_n806__ = new_new_n780__ & new_new_n804__;
  assign new_new_n807__ = ~G37 & ~new_new_n805__;
  assign G395 = ~new_new_n806__ & new_new_n807__;
  assign new_new_n809__ = G303 & ~G305;
  assign new_new_n810__ = ~G303 & G305;
  assign new_new_n811__ = ~new_new_n809__ & ~new_new_n810__;
  assign new_new_n812__ = ~G288 & G290;
  assign new_new_n813__ = G288 & ~G290;
  assign new_new_n814__ = ~new_new_n812__ & ~new_new_n813__;
  assign new_new_n815__ = new_new_n811__ & new_new_n814__;
  assign new_new_n816__ = ~new_new_n811__ & ~new_new_n814__;
  assign new_new_n817__ = ~new_new_n815__ & ~new_new_n816__;
  assign new_new_n818__ = ~G299 & ~new_new_n771__;
  assign new_new_n819__ = G299 & new_new_n771__;
  assign new_new_n820__ = ~new_new_n818__ & ~new_new_n819__;
  assign new_new_n821__ = new_new_n515__ & ~new_new_n820__;
  assign new_new_n822__ = new_new_n507__ & ~new_new_n820__;
  assign new_new_n823__ = ~new_new_n507__ & new_new_n820__;
  assign new_new_n824__ = ~new_new_n822__ & ~new_new_n823__;
  assign new_new_n825__ = ~new_new_n515__ & ~new_new_n824__;
  assign new_new_n826__ = ~new_new_n821__ & ~new_new_n825__;
  assign new_new_n827__ = new_new_n817__ & ~new_new_n826__;
  assign new_new_n828__ = ~new_new_n817__ & new_new_n826__;
  assign new_new_n829__ = ~new_new_n827__ & ~new_new_n828__;
  assign new_new_n830__ = G868 & ~new_new_n829__;
  assign new_new_n831__ = ~G868 & new_new_n768__;
  assign G295 = new_new_n830__ | new_new_n831__;
  assign new_new_n833__ = G286 & ~G301;
  assign new_new_n834__ = ~G286 & G301;
  assign new_new_n835__ = ~new_new_n833__ & ~new_new_n834__;
  assign new_new_n836__ = new_new_n824__ & new_new_n835__;
  assign new_new_n837__ = ~new_new_n824__ & ~new_new_n835__;
  assign new_new_n838__ = ~new_new_n836__ & ~new_new_n837__;
  assign new_new_n839__ = ~new_new_n817__ & new_new_n838__;
  assign new_new_n840__ = new_new_n817__ & ~new_new_n838__;
  assign new_new_n841__ = ~G37 & ~new_new_n839__;
  assign G397 = ~new_new_n840__ & new_new_n841__;
  assign new_new_n843__ = ~G1384 & ~G164;
  assign new_new_n844__ = G40 & G160;
  assign new_new_n845__ = new_new_n843__ & new_new_n844__;
  assign new_new_n846__ = G2090 & new_new_n845__;
  assign new_new_n847__ = G1971 & ~new_new_n845__;
  assign new_new_n848__ = G8 & ~new_new_n846__;
  assign new_new_n849__ = ~new_new_n847__ & new_new_n848__;
  assign new_new_n850__ = G8 & G303;
  assign new_new_n851__ = ~new_new_n849__ & new_new_n850__;
  assign new_new_n852__ = ~G303 & new_new_n849__;
  assign new_new_n853__ = ~new_new_n851__ & ~new_new_n852__;
  assign new_new_n854__ = G1956 & ~new_new_n845__;
  assign new_new_n855__ = G2072 & new_new_n845__;
  assign new_new_n856__ = ~new_new_n854__ & ~new_new_n855__;
  assign new_new_n857__ = ~G299 & new_new_n856__;
  assign new_new_n858__ = G1348 & ~new_new_n845__;
  assign new_new_n859__ = G2067 & new_new_n845__;
  assign new_new_n860__ = ~new_new_n858__ & ~new_new_n859__;
  assign new_new_n861__ = ~new_new_n507__ & new_new_n860__;
  assign new_new_n862__ = G1996 & new_new_n845__;
  assign new_new_n863__ = new_new_n507__ & ~new_new_n860__;
  assign new_new_n864__ = G1341 & ~new_new_n845__;
  assign new_new_n865__ = ~new_new_n456__ & ~new_new_n862__;
  assign new_new_n866__ = ~new_new_n864__ & new_new_n865__;
  assign new_new_n867__ = ~new_new_n863__ & new_new_n866__;
  assign new_new_n868__ = ~new_new_n857__ & ~new_new_n861__;
  assign new_new_n869__ = ~new_new_n867__ & new_new_n868__;
  assign new_new_n870__ = G2084 & new_new_n845__;
  assign new_new_n871__ = G1966 & ~new_new_n845__;
  assign new_new_n872__ = G8 & ~new_new_n870__;
  assign new_new_n873__ = ~new_new_n871__ & new_new_n872__;
  assign new_new_n874__ = ~G286 & new_new_n873__;
  assign new_new_n875__ = G8 & G286;
  assign new_new_n876__ = ~new_new_n873__ & new_new_n875__;
  assign new_new_n877__ = ~new_new_n874__ & ~new_new_n876__;
  assign new_new_n878__ = G1961 & ~new_new_n845__;
  assign new_new_n879__ = G2078 & new_new_n845__;
  assign new_new_n880__ = ~new_new_n878__ & ~new_new_n879__;
  assign new_new_n881__ = G301 & ~new_new_n880__;
  assign new_new_n882__ = ~G301 & new_new_n880__;
  assign new_new_n883__ = G299 & ~new_new_n856__;
  assign new_new_n884__ = G8 & ~G1981;
  assign new_new_n885__ = ~G305 & new_new_n884__;
  assign new_new_n886__ = ~new_new_n845__ & new_new_n885__;
  assign new_new_n887__ = G8 & ~G1976;
  assign new_new_n888__ = G8 & ~new_new_n887__;
  assign new_new_n889__ = G288 & new_new_n888__;
  assign new_new_n890__ = ~new_new_n845__ & new_new_n889__;
  assign new_new_n891__ = G8 & ~new_new_n884__;
  assign new_new_n892__ = G305 & new_new_n891__;
  assign new_new_n893__ = ~new_new_n845__ & new_new_n892__;
  assign new_new_n894__ = ~G288 & new_new_n887__;
  assign new_new_n895__ = ~new_new_n845__ & new_new_n894__;
  assign new_new_n896__ = ~new_new_n886__ & ~new_new_n890__;
  assign new_new_n897__ = ~new_new_n893__ & ~new_new_n895__;
  assign new_new_n898__ = new_new_n896__ & new_new_n897__;
  assign new_new_n899__ = ~new_new_n881__ & ~new_new_n882__;
  assign new_new_n900__ = ~new_new_n883__ & new_new_n898__;
  assign new_new_n901__ = new_new_n899__ & new_new_n900__;
  assign new_new_n902__ = new_new_n853__ & new_new_n901__;
  assign new_new_n903__ = ~new_new_n869__ & new_new_n877__;
  assign new_new_n904__ = new_new_n902__ & new_new_n903__;
  assign new_new_n905__ = new_new_n874__ & new_new_n898__;
  assign new_new_n906__ = new_new_n853__ & new_new_n905__;
  assign new_new_n907__ = new_new_n852__ & new_new_n898__;
  assign new_new_n908__ = ~new_new_n893__ & new_new_n895__;
  assign new_new_n909__ = new_new_n882__ & new_new_n898__;
  assign new_new_n910__ = new_new_n853__ & new_new_n909__;
  assign new_new_n911__ = new_new_n877__ & new_new_n910__;
  assign new_new_n912__ = ~new_new_n886__ & ~new_new_n908__;
  assign new_new_n913__ = ~new_new_n907__ & new_new_n912__;
  assign new_new_n914__ = ~new_new_n906__ & new_new_n913__;
  assign new_new_n915__ = ~new_new_n904__ & new_new_n914__;
  assign new_new_n916__ = ~new_new_n911__ & new_new_n915__;
  assign new_new_n917__ = ~new_new_n843__ & new_new_n844__;
  assign new_new_n918__ = ~G2067 & ~new_new_n680__;
  assign new_new_n919__ = new_new_n917__ & new_new_n918__;
  assign new_new_n920__ = G1996 & new_new_n628__;
  assign new_new_n921__ = new_new_n917__ & new_new_n920__;
  assign new_new_n922__ = G2067 & new_new_n680__;
  assign new_new_n923__ = new_new_n917__ & new_new_n922__;
  assign new_new_n924__ = ~G1996 & ~new_new_n628__;
  assign new_new_n925__ = new_new_n917__ & new_new_n924__;
  assign new_new_n926__ = G1986 & G290;
  assign new_new_n927__ = new_new_n917__ & new_new_n926__;
  assign new_new_n928__ = ~G1986 & ~G290;
  assign new_new_n929__ = new_new_n917__ & new_new_n928__;
  assign new_new_n930__ = ~G1991 & ~new_new_n711__;
  assign new_new_n931__ = new_new_n917__ & new_new_n930__;
  assign new_new_n932__ = ~new_new_n929__ & ~new_new_n931__;
  assign new_new_n933__ = G1991 & new_new_n711__;
  assign new_new_n934__ = new_new_n917__ & new_new_n933__;
  assign new_new_n935__ = ~new_new_n919__ & ~new_new_n921__;
  assign new_new_n936__ = ~new_new_n923__ & ~new_new_n925__;
  assign new_new_n937__ = ~new_new_n927__ & ~new_new_n934__;
  assign new_new_n938__ = new_new_n936__ & new_new_n937__;
  assign new_new_n939__ = new_new_n932__ & new_new_n935__;
  assign new_new_n940__ = new_new_n938__ & new_new_n939__;
  assign new_new_n941__ = ~new_new_n916__ & new_new_n940__;
  assign new_new_n942__ = ~new_new_n931__ & new_new_n933__;
  assign new_new_n943__ = ~new_new_n921__ & ~new_new_n932__;
  assign new_new_n944__ = ~new_new_n942__ & new_new_n943__;
  assign new_new_n945__ = ~new_new_n925__ & ~new_new_n944__;
  assign new_new_n946__ = ~new_new_n923__ & ~new_new_n945__;
  assign new_new_n947__ = ~new_new_n919__ & ~new_new_n946__;
  assign G329 = new_new_n941__ | ~new_new_n947__;
  assign new_new_n949__ = G319 & ~G227;
  assign new_new_n950__ = ~G229 & new_new_n949__;
  assign new_new_n951__ = ~G401 & new_new_n950__;
  assign new_new_n952__ = ~G395 & new_new_n951__;
  assign G308 = ~G397 & new_new_n952__;
  assign G218 = ~G44;
  assign G219 = ~G132;
  assign G220 = ~G82;
  assign G221 = ~G96;
  assign G235 = ~G69;
  assign G236 = ~G120;
  assign G237 = ~G57;
  assign G238 = ~G108;
  assign G261 = ~G325;
  assign G166 = ~G303;
  assign G168 = ~G286;
  assign G171 = ~G301;
  assign G150 = ~G311;
  assign G225 = ~G308;
  assign G169 = _IN_G169 ;
  assign G174 = _IN_G174 ;
  assign G177 = _IN_G177 ;
  assign G178 = _IN_G178 ;
  assign G179 = _IN_G179 ;
  assign G180 = _IN_G180 ;
  assign G181 = _IN_G181 ;
  assign G182 = _IN_G182 ;
  assign G183 = _IN_G183 ;
  assign G184 = _IN_G184 ;
  assign G185 = _IN_G185 ;
  assign G186 = _IN_G186 ;
  assign G189 = _IN_G189 ;
  assign G190 = _IN_G190 ;
  assign G191 = _IN_G191 ;
  assign G192 = _IN_G192 ;
  assign G193 = _IN_G193 ;
  assign G194 = _IN_G194 ;
  assign G195 = _IN_G195 ;
  assign G196 = _IN_G196 ;
  assign G197 = _IN_G197 ;
  assign G198 = _IN_G198 ;
  assign G199 = _IN_G199 ;
  assign G200 = _IN_G200 ;
  assign G201 = _IN_G201 ;
  assign G202 = _IN_G202 ;
  assign G203 = _IN_G203 ;
  assign G204 = _IN_G204 ;
  assign G205 = _IN_G205 ;
  assign G206 = _IN_G206 ;
  assign G207 = _IN_G207 ;
  assign G208 = _IN_G208 ;
  assign G209 = _IN_G209 ;
  assign G210 = _IN_G210 ;
  assign G211 = _IN_G211 ;
  assign G212 = _IN_G212 ;
  assign G213 = _IN_G213 ;
  assign G214 = _IN_G214 ;
  assign G215 = _IN_G215 ;
  assign G239 = _IN_G239 ;
  assign G240 = _IN_G240 ;
  assign G241 = _IN_G241 ;
  assign G242 = _IN_G242 ;
  assign G243 = _IN_G243 ;
  assign G244 = _IN_G244 ;
  assign G245 = _IN_G245 ;
  assign G246 = _IN_G246 ;
  assign G247 = _IN_G247 ;
  assign G248 = _IN_G248 ;
  assign G249 = _IN_G249 ;
  assign G250 = _IN_G250 ;
  assign G251 = _IN_G251 ;
  assign G252 = _IN_G252 ;
  assign G253 = _IN_G253 ;
  assign G254 = _IN_G254 ;
  assign G255 = _IN_G255 ;
  assign G256 = _IN_G256 ;
  assign G257 = _IN_G257 ;
  assign G262 = _IN_G262 ;
  assign G263 = _IN_G263 ;
  assign G264 = _IN_G264 ;
  assign G265 = _IN_G265 ;
  assign G266 = _IN_G266 ;
  assign G267 = _IN_G267 ;
  assign G268 = _IN_G268 ;
  assign G269 = _IN_G269 ;
  assign G270 = _IN_G270 ;
  assign G271 = _IN_G271 ;
  assign G272 = _IN_G272 ;
  assign G273 = _IN_G273 ;
  assign G274 = _IN_G274 ;
  assign G275 = _IN_G275 ;
  assign G276 = _IN_G276 ;
  assign G277 = _IN_G277 ;
  assign G278 = _IN_G278 ;
  assign G279 = _IN_G279 ;
  // assign G350 = G452;
  // assign G335 = G452;
  // assign G409 = G452;
  // assign G369 = G1083;
  // assign G367 = G1083;
  // assign G411 = G2066;
  // assign G337 = G2066;
  // assign G384 = G2066;
  // assign G391 = G452;
  // assign G321 = G284;
  // assign G280 = G297;
  // assign G323 = G282;
  // assign G331 = G295;
  // assign G231 = 1'b0;
endmodule


