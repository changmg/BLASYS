// Benchmark "ex" written by ABC on Fri Jul  1 13:59:12 2022

module ex ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m,
    F  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m;
  output F;
  assign F = c & g;
endmodule


