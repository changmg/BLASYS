// Benchmark "ex" written by ABC on Thu Jul 14 00:20:05 2022

module ex ( 
    a, b, c, d, e, f,
    F  );
  input  a, b, c, d, e, f;
  output F;
  assign F = e;
endmodule


