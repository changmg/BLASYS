module adder8_1(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , po0 , po1 , po2 , po3 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 ;
  output po0 , po1 , po2 , po3 ;
  wire new_n8, new_n9, new_n10, new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31;
  assign new_n8 = ~pi0 & ~pi3 ;
  assign new_n9 = pi0 & pi3 ;
  assign new_n10 = ~new_n8 & ~new_n9 ;
  assign new_n11 = ~pi6 & ~new_n10 ;
  assign new_n12 = pi6 & new_n10 ;
  assign new_n13 = ~new_n11 & ~new_n12 ;
  assign new_n14 = pi1 & pi4 ;
  assign new_n15 = ~pi1 & ~pi4 ;
  assign new_n16 = ~new_n14 & ~new_n15 ;
  assign new_n17 = ~pi6 & ~new_n8 ;
  assign new_n18 = ~new_n9 & ~new_n17 ;
  assign new_n19 = ~new_n16 & ~new_n18 ;
  assign new_n20 = new_n16 & new_n18 ;
  assign new_n21 = ~new_n19 & ~new_n20 ;
  assign new_n22 = ~pi2 & ~pi5 ;
  assign new_n23 = pi2 & pi5 ;
  assign new_n24 = ~new_n22 & ~new_n23 ;
  assign new_n25 = ~new_n15 & ~new_n18 ;
  assign new_n26 = ~new_n14 & ~new_n25 ;
  assign new_n27 = ~new_n24 & ~new_n26 ;
  assign new_n28 = new_n24 & new_n26 ;
  assign new_n29 = ~new_n27 & ~new_n28 ;
  assign new_n30 = ~new_n22 & ~new_n26 ;
  assign new_n31 = ~new_n23 & ~new_n30 ;
  assign po0 = new_n13 ;
  assign po1 = new_n21 ;
  assign po2 = new_n29 ;
  assign po3 = new_n31 ;
endmodule
