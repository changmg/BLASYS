// Benchmark "c7552" written by ABC on Sat Jul 16 14:45:52 2022

module c7552 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52;
  wire new_n260_, new_n261_, new_n263_, new_n264_, new_n266_, new_n267_,
    new_n269_, new_n270_, new_n273_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n949_, new_n950_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_,
    new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_,
    new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_,
    new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1303_, new_n1304_, new_n1306_, new_n1307_,
    new_n1309_, new_n1310_, new_n1311_, new_n1313_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1330_,
    new_n1331_, new_n1332_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1343_, new_n1344_,
    new_n1345_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1353_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1369_, new_n1370_, new_n1371_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1378_, new_n1379_, new_n1381_, new_n1382_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1389_, new_n1390_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1401_, new_n1402_, new_n1403_, new_n1405_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1411_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1419_, new_n1420_,
    new_n1421_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1428_,
    new_n1429_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_,
    new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_,
    new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_,
    new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_,
    new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_,
    new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_;
  assign po00 = pi001 | pi019;
  assign new_n260_ = pi072 & pi106;
  assign new_n261_ = pi150 & pi162;
  assign po01 = ~new_n260_ | ~new_n261_;
  assign new_n263_ = pi074 & pi132;
  assign new_n264_ = pi140 & pi152;
  assign po02 = ~new_n263_ | ~new_n264_;
  assign new_n266_ = pi104 & pi105;
  assign new_n267_ = pi107 & pi108;
  assign po03 = ~new_n266_ | ~new_n267_;
  assign new_n269_ = pi084 & pi094;
  assign new_n270_ = pi110 & pi121;
  assign po04 = ~new_n269_ | ~new_n270_;
  assign po05 = pi001 | ~pi163;
  assign new_n273_ = ~pi001 & pi065;
  assign po06 = ~pi066 | ~new_n273_;
  assign po07 = pi000 & pi085;
  assign new_n276_ = ~pi004 & pi011;
  assign new_n277_ = ~pi184 & new_n276_;
  assign new_n278_ = pi004 & pi151;
  assign new_n279_ = ~new_n276_ & ~new_n278_;
  assign new_n280_ = ~pi004 & pi184;
  assign new_n281_ = new_n279_ & new_n280_;
  assign new_n282_ = ~new_n277_ & ~new_n281_;
  assign new_n283_ = pi203 & new_n282_;
  assign new_n284_ = ~pi203 & ~new_n282_;
  assign po08 = ~new_n283_ & ~new_n284_;
  assign new_n286_ = pi171 & pi204;
  assign new_n287_ = pi170 & new_n286_;
  assign new_n288_ = pi010 & ~new_n287_;
  assign new_n289_ = pi004 & pi157;
  assign new_n290_ = ~pi004 & pi051;
  assign new_n291_ = ~new_n289_ & ~new_n290_;
  assign new_n292_ = pi188 & new_n291_;
  assign new_n293_ = pi004 & pi158;
  assign new_n294_ = ~pi004 & pi005;
  assign new_n295_ = ~new_n293_ & ~new_n294_;
  assign new_n296_ = pi187 & new_n295_;
  assign new_n297_ = ~pi187 & ~new_n295_;
  assign new_n298_ = pi004 & pi159;
  assign new_n299_ = ~pi004 & pi006;
  assign new_n300_ = ~new_n298_ & ~new_n299_;
  assign new_n301_ = pi186 & new_n300_;
  assign new_n302_ = pi004 & pi160;
  assign new_n303_ = ~pi004 & pi007;
  assign new_n304_ = ~new_n302_ & ~new_n303_;
  assign new_n305_ = ~pi185 & ~new_n304_;
  assign new_n306_ = pi185 & new_n304_;
  assign new_n307_ = ~new_n305_ & ~new_n306_;
  assign new_n308_ = new_n277_ & new_n307_;
  assign new_n309_ = ~pi186 & ~new_n300_;
  assign new_n310_ = ~new_n305_ & ~new_n309_;
  assign new_n311_ = ~new_n308_ & new_n310_;
  assign new_n312_ = ~new_n301_ & ~new_n311_;
  assign new_n313_ = ~new_n297_ & ~new_n312_;
  assign new_n314_ = ~new_n296_ & ~new_n313_;
  assign new_n315_ = ~new_n292_ & new_n314_;
  assign new_n316_ = ~pi188 & ~new_n291_;
  assign new_n317_ = new_n282_ & new_n307_;
  assign new_n318_ = pi203 & new_n317_;
  assign new_n319_ = ~new_n301_ & ~new_n309_;
  assign new_n320_ = ~new_n296_ & ~new_n297_;
  assign new_n321_ = new_n319_ & new_n320_;
  assign new_n322_ = ~new_n292_ & new_n321_;
  assign new_n323_ = new_n318_ & new_n322_;
  assign new_n324_ = ~new_n316_ & ~new_n323_;
  assign new_n325_ = ~new_n315_ & new_n324_;
  assign new_n326_ = pi004 & pi155;
  assign new_n327_ = ~pi004 & pi063;
  assign new_n328_ = ~new_n326_ & ~new_n327_;
  assign new_n329_ = ~pi190 & ~new_n328_;
  assign new_n330_ = pi190 & new_n328_;
  assign new_n331_ = ~new_n329_ & ~new_n330_;
  assign new_n332_ = pi004 & pi156;
  assign new_n333_ = ~pi004 & pi064;
  assign new_n334_ = ~new_n332_ & ~new_n333_;
  assign new_n335_ = ~pi189 & ~new_n334_;
  assign new_n336_ = pi189 & new_n334_;
  assign new_n337_ = ~new_n335_ & ~new_n336_;
  assign new_n338_ = new_n331_ & new_n337_;
  assign new_n339_ = pi004 & pi154;
  assign new_n340_ = ~pi004 & pi062;
  assign new_n341_ = ~new_n339_ & ~new_n340_;
  assign new_n342_ = ~pi191 & ~new_n341_;
  assign new_n343_ = pi191 & new_n341_;
  assign new_n344_ = ~new_n342_ & ~new_n343_;
  assign new_n345_ = pi004 & pi153;
  assign new_n346_ = ~pi004 & pi050;
  assign new_n347_ = ~new_n345_ & ~new_n346_;
  assign new_n348_ = pi192 & new_n347_;
  assign new_n349_ = ~pi192 & ~new_n347_;
  assign new_n350_ = ~new_n348_ & ~new_n349_;
  assign new_n351_ = new_n344_ & new_n350_;
  assign new_n352_ = new_n338_ & new_n351_;
  assign new_n353_ = ~new_n325_ & new_n352_;
  assign new_n354_ = new_n331_ & new_n335_;
  assign new_n355_ = ~new_n329_ & ~new_n354_;
  assign new_n356_ = new_n351_ & ~new_n355_;
  assign new_n357_ = new_n342_ & ~new_n348_;
  assign new_n358_ = ~new_n349_ & ~new_n357_;
  assign new_n359_ = ~new_n356_ & new_n358_;
  assign new_n360_ = ~new_n353_ & new_n359_;
  assign new_n361_ = pi004 & pi148;
  assign new_n362_ = ~pi004 & pi049;
  assign new_n363_ = ~new_n361_ & ~new_n362_;
  assign new_n364_ = pi195 & new_n363_;
  assign new_n365_ = pi004 & pi139;
  assign new_n366_ = ~pi004 & pi060;
  assign new_n367_ = ~new_n365_ & ~new_n366_;
  assign new_n368_ = ~pi194 & ~new_n367_;
  assign new_n369_ = pi194 & new_n367_;
  assign new_n370_ = ~new_n368_ & ~new_n369_;
  assign new_n371_ = ~new_n364_ & new_n370_;
  assign new_n372_ = pi004 & pi147;
  assign new_n373_ = ~pi004 & pi048;
  assign new_n374_ = ~new_n372_ & ~new_n373_;
  assign new_n375_ = ~pi196 & ~new_n374_;
  assign new_n376_ = pi196 & new_n374_;
  assign new_n377_ = ~new_n375_ & ~new_n376_;
  assign new_n378_ = ~pi195 & ~new_n363_;
  assign new_n379_ = new_n377_ & ~new_n378_;
  assign new_n380_ = new_n371_ & new_n379_;
  assign new_n381_ = pi004 & pi145;
  assign new_n382_ = ~pi004 & pi013;
  assign new_n383_ = ~new_n381_ & ~new_n382_;
  assign new_n384_ = pi198 & new_n383_;
  assign new_n385_ = ~pi198 & ~new_n383_;
  assign new_n386_ = ~new_n384_ & ~new_n385_;
  assign new_n387_ = pi004 & pi146;
  assign new_n388_ = ~pi004 & pi061;
  assign new_n389_ = ~new_n387_ & ~new_n388_;
  assign new_n390_ = ~pi197 & ~new_n389_;
  assign new_n391_ = pi197 & new_n389_;
  assign new_n392_ = ~new_n390_ & ~new_n391_;
  assign new_n393_ = new_n386_ & new_n392_;
  assign new_n394_ = new_n380_ & new_n393_;
  assign new_n395_ = ~new_n360_ & new_n394_;
  assign new_n396_ = ~new_n364_ & ~new_n378_;
  assign new_n397_ = new_n368_ & new_n396_;
  assign new_n398_ = new_n377_ & new_n397_;
  assign new_n399_ = ~new_n375_ & ~new_n398_;
  assign new_n400_ = new_n393_ & ~new_n399_;
  assign new_n401_ = new_n377_ & new_n378_;
  assign new_n402_ = new_n393_ & new_n401_;
  assign new_n403_ = ~new_n384_ & new_n390_;
  assign new_n404_ = ~new_n385_ & ~new_n403_;
  assign new_n405_ = ~new_n402_ & new_n404_;
  assign new_n406_ = ~new_n400_ & new_n405_;
  assign new_n407_ = ~new_n395_ & new_n406_;
  assign new_n408_ = pi004 & pi143;
  assign new_n409_ = ~pi004 & pi008;
  assign new_n410_ = ~new_n408_ & ~new_n409_;
  assign new_n411_ = ~pi200 & ~new_n410_;
  assign new_n412_ = pi200 & new_n410_;
  assign new_n413_ = ~new_n411_ & ~new_n412_;
  assign new_n414_ = pi004 & pi144;
  assign new_n415_ = ~pi004 & pi009;
  assign new_n416_ = ~new_n414_ & ~new_n415_;
  assign new_n417_ = ~pi199 & ~new_n416_;
  assign new_n418_ = pi199 & new_n416_;
  assign new_n419_ = ~new_n417_ & ~new_n418_;
  assign new_n420_ = new_n413_ & new_n419_;
  assign new_n421_ = pi004 & pi141;
  assign new_n422_ = ~pi004 & pi028;
  assign new_n423_ = ~new_n421_ & ~new_n422_;
  assign new_n424_ = ~pi202 & ~new_n423_;
  assign new_n425_ = pi202 & new_n423_;
  assign new_n426_ = ~new_n424_ & ~new_n425_;
  assign new_n427_ = pi004 & pi142;
  assign new_n428_ = ~pi004 & pi014;
  assign new_n429_ = ~new_n427_ & ~new_n428_;
  assign new_n430_ = pi201 & new_n429_;
  assign new_n431_ = ~pi201 & ~new_n429_;
  assign new_n432_ = ~new_n430_ & ~new_n431_;
  assign new_n433_ = new_n426_ & new_n432_;
  assign new_n434_ = new_n420_ & new_n433_;
  assign new_n435_ = ~new_n407_ & new_n434_;
  assign new_n436_ = new_n413_ & new_n417_;
  assign new_n437_ = ~new_n411_ & ~new_n436_;
  assign new_n438_ = ~new_n430_ & ~new_n437_;
  assign new_n439_ = ~new_n431_ & ~new_n438_;
  assign new_n440_ = ~new_n424_ & new_n439_;
  assign new_n441_ = ~new_n425_ & ~new_n440_;
  assign new_n442_ = ~new_n435_ & ~new_n441_;
  assign new_n443_ = pi002 & pi003;
  assign new_n444_ = pi004 & ~pi079;
  assign new_n445_ = ~new_n443_ & ~new_n444_;
  assign new_n446_ = ~pi178 & new_n445_;
  assign new_n447_ = pi178 & ~new_n445_;
  assign new_n448_ = ~new_n446_ & ~new_n447_;
  assign new_n449_ = ~pi004 & pi067;
  assign new_n450_ = pi004 & pi080;
  assign new_n451_ = ~new_n449_ & ~new_n450_;
  assign new_n452_ = ~pi177 & ~new_n451_;
  assign new_n453_ = pi177 & new_n451_;
  assign new_n454_ = ~new_n452_ & ~new_n453_;
  assign new_n455_ = ~pi004 & pi070;
  assign new_n456_ = pi004 & pi081;
  assign new_n457_ = ~new_n455_ & ~new_n456_;
  assign new_n458_ = ~pi176 & ~new_n457_;
  assign new_n459_ = pi176 & new_n457_;
  assign new_n460_ = ~new_n458_ & ~new_n459_;
  assign new_n461_ = ~pi004 & pi068;
  assign new_n462_ = pi004 & pi082;
  assign new_n463_ = ~new_n461_ & ~new_n462_;
  assign new_n464_ = ~pi175 & ~new_n463_;
  assign new_n465_ = pi175 & new_n463_;
  assign new_n466_ = ~new_n464_ & ~new_n465_;
  assign new_n467_ = ~pi004 & pi071;
  assign new_n468_ = pi004 & pi073;
  assign new_n469_ = ~new_n467_ & ~new_n468_;
  assign new_n470_ = ~pi174 & ~new_n469_;
  assign new_n471_ = pi174 & new_n469_;
  assign new_n472_ = ~new_n470_ & ~new_n471_;
  assign new_n473_ = new_n466_ & new_n472_;
  assign new_n474_ = new_n460_ & new_n473_;
  assign new_n475_ = new_n454_ & new_n474_;
  assign new_n476_ = new_n448_ & new_n475_;
  assign new_n477_ = pi004 & ~pi077;
  assign new_n478_ = ~new_n443_ & ~new_n477_;
  assign new_n479_ = ~pi180 & new_n478_;
  assign new_n480_ = pi180 & ~new_n478_;
  assign new_n481_ = ~new_n479_ & ~new_n480_;
  assign new_n482_ = pi004 & ~pi078;
  assign new_n483_ = ~new_n443_ & ~new_n482_;
  assign new_n484_ = ~pi179 & new_n483_;
  assign new_n485_ = pi179 & ~new_n483_;
  assign new_n486_ = ~new_n484_ & ~new_n485_;
  assign new_n487_ = new_n481_ & new_n486_;
  assign new_n488_ = pi004 & ~pi076;
  assign new_n489_ = ~new_n443_ & ~new_n488_;
  assign new_n490_ = ~pi181 & new_n489_;
  assign new_n491_ = pi181 & ~new_n489_;
  assign new_n492_ = ~new_n490_ & ~new_n491_;
  assign new_n493_ = pi004 & ~pi075;
  assign new_n494_ = ~new_n443_ & ~new_n493_;
  assign new_n495_ = ~pi182 & new_n494_;
  assign new_n496_ = pi182 & ~new_n494_;
  assign new_n497_ = ~new_n495_ & ~new_n496_;
  assign new_n498_ = new_n492_ & new_n497_;
  assign new_n499_ = new_n487_ & new_n498_;
  assign new_n500_ = new_n476_ & new_n499_;
  assign new_n501_ = ~new_n442_ & new_n500_;
  assign new_n502_ = new_n466_ & new_n470_;
  assign new_n503_ = ~new_n458_ & ~new_n464_;
  assign new_n504_ = ~new_n502_ & new_n503_;
  assign new_n505_ = ~new_n459_ & ~new_n504_;
  assign new_n506_ = ~new_n453_ & new_n505_;
  assign new_n507_ = ~new_n452_ & ~new_n506_;
  assign new_n508_ = ~new_n447_ & ~new_n507_;
  assign new_n509_ = ~new_n446_ & ~new_n508_;
  assign new_n510_ = new_n499_ & ~new_n509_;
  assign new_n511_ = new_n481_ & new_n484_;
  assign new_n512_ = ~new_n479_ & ~new_n511_;
  assign new_n513_ = ~new_n490_ & new_n512_;
  assign new_n514_ = ~new_n491_ & ~new_n513_;
  assign new_n515_ = ~new_n496_ & new_n514_;
  assign new_n516_ = ~new_n495_ & ~new_n515_;
  assign new_n517_ = ~new_n510_ & new_n516_;
  assign new_n518_ = ~new_n501_ & new_n517_;
  assign new_n519_ = pi004 & ~pi138;
  assign new_n520_ = ~new_n443_ & ~new_n519_;
  assign new_n521_ = pi167 & ~new_n520_;
  assign new_n522_ = pi004 & ~pi131;
  assign new_n523_ = ~new_n443_ & ~new_n522_;
  assign new_n524_ = ~pi166 & new_n523_;
  assign new_n525_ = pi166 & ~new_n523_;
  assign new_n526_ = ~new_n524_ & ~new_n525_;
  assign new_n527_ = ~new_n521_ & new_n526_;
  assign new_n528_ = pi004 & ~pi137;
  assign new_n529_ = ~new_n443_ & ~new_n528_;
  assign new_n530_ = ~pi052 & new_n529_;
  assign new_n531_ = pi052 & ~new_n529_;
  assign new_n532_ = ~new_n530_ & ~new_n531_;
  assign new_n533_ = ~pi167 & new_n520_;
  assign new_n534_ = new_n532_ & ~new_n533_;
  assign new_n535_ = new_n527_ & new_n534_;
  assign new_n536_ = pi004 & ~pi135;
  assign new_n537_ = ~new_n443_ & ~new_n536_;
  assign new_n538_ = pi169 & ~new_n537_;
  assign new_n539_ = ~pi169 & new_n537_;
  assign new_n540_ = ~new_n538_ & ~new_n539_;
  assign new_n541_ = pi004 & ~pi136;
  assign new_n542_ = ~new_n443_ & ~new_n541_;
  assign new_n543_ = ~pi168 & new_n542_;
  assign new_n544_ = pi168 & ~new_n542_;
  assign new_n545_ = ~new_n543_ & ~new_n544_;
  assign new_n546_ = new_n540_ & new_n545_;
  assign new_n547_ = new_n535_ & new_n546_;
  assign new_n548_ = ~new_n518_ & new_n547_;
  assign new_n549_ = ~new_n521_ & ~new_n533_;
  assign new_n550_ = new_n524_ & new_n549_;
  assign new_n551_ = new_n532_ & new_n550_;
  assign new_n552_ = ~new_n530_ & ~new_n551_;
  assign new_n553_ = new_n546_ & ~new_n552_;
  assign new_n554_ = new_n532_ & new_n533_;
  assign new_n555_ = new_n546_ & new_n554_;
  assign new_n556_ = ~new_n538_ & new_n543_;
  assign new_n557_ = ~new_n539_ & ~new_n556_;
  assign new_n558_ = ~new_n555_ & new_n557_;
  assign new_n559_ = ~new_n553_ & new_n558_;
  assign new_n560_ = ~new_n548_ & new_n559_;
  assign new_n561_ = pi170 & pi204;
  assign new_n562_ = pi010 & ~new_n561_;
  assign new_n563_ = ~pi010 & new_n561_;
  assign new_n564_ = ~new_n562_ & ~new_n563_;
  assign new_n565_ = pi010 & new_n286_;
  assign new_n566_ = ~pi010 & ~new_n286_;
  assign new_n567_ = ~new_n565_ & ~new_n566_;
  assign new_n568_ = new_n564_ & ~new_n567_;
  assign new_n569_ = ~new_n560_ & new_n568_;
  assign po09 = new_n288_ | new_n569_;
  assign new_n571_ = pi004 & pi127;
  assign new_n572_ = ~new_n294_ & ~new_n571_;
  assign new_n573_ = ~pi004 & ~pi033;
  assign new_n574_ = pi004 & pi187;
  assign new_n575_ = ~new_n573_ & ~new_n574_;
  assign new_n576_ = ~new_n572_ & new_n575_;
  assign new_n577_ = pi004 & pi128;
  assign new_n578_ = ~new_n299_ & ~new_n577_;
  assign new_n579_ = ~pi004 & ~pi034;
  assign new_n580_ = pi004 & pi186;
  assign new_n581_ = ~new_n579_ & ~new_n580_;
  assign new_n582_ = new_n578_ & ~new_n581_;
  assign new_n583_ = pi004 & pi129;
  assign new_n584_ = ~new_n303_ & ~new_n583_;
  assign new_n585_ = ~pi004 & ~pi032;
  assign new_n586_ = pi004 & pi185;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign new_n588_ = new_n584_ & ~new_n587_;
  assign new_n589_ = ~pi004 & ~pi030;
  assign new_n590_ = new_n276_ & ~new_n589_;
  assign new_n591_ = ~new_n588_ & new_n590_;
  assign new_n592_ = ~new_n584_ & new_n587_;
  assign new_n593_ = ~new_n578_ & new_n581_;
  assign new_n594_ = ~new_n592_ & ~new_n593_;
  assign new_n595_ = ~new_n591_ & new_n594_;
  assign new_n596_ = ~new_n582_ & ~new_n595_;
  assign new_n597_ = ~new_n576_ & ~new_n596_;
  assign new_n598_ = pi004 & pi126;
  assign new_n599_ = ~new_n290_ & ~new_n598_;
  assign new_n600_ = ~pi004 & ~pi031;
  assign new_n601_ = pi004 & pi188;
  assign new_n602_ = ~new_n600_ & ~new_n601_;
  assign new_n603_ = new_n599_ & ~new_n602_;
  assign new_n604_ = new_n572_ & ~new_n575_;
  assign new_n605_ = ~new_n603_ & ~new_n604_;
  assign new_n606_ = ~new_n597_ & new_n605_;
  assign new_n607_ = ~new_n599_ & new_n602_;
  assign new_n608_ = ~new_n588_ & ~new_n603_;
  assign new_n609_ = ~new_n604_ & ~new_n607_;
  assign new_n610_ = new_n608_ & new_n609_;
  assign new_n611_ = ~new_n276_ & new_n589_;
  assign new_n612_ = pi047 & ~new_n590_;
  assign new_n613_ = ~new_n611_ & new_n612_;
  assign new_n614_ = ~new_n576_ & ~new_n582_;
  assign new_n615_ = new_n594_ & new_n614_;
  assign new_n616_ = new_n613_ & new_n615_;
  assign new_n617_ = new_n610_ & new_n616_;
  assign new_n618_ = ~new_n607_ & ~new_n617_;
  assign new_n619_ = ~new_n606_ & new_n618_;
  assign new_n620_ = pi004 & pi122;
  assign new_n621_ = ~new_n346_ & ~new_n620_;
  assign new_n622_ = ~pi004 & ~pi018;
  assign new_n623_ = pi004 & pi192;
  assign new_n624_ = ~new_n622_ & ~new_n623_;
  assign new_n625_ = ~new_n621_ & new_n624_;
  assign new_n626_ = pi004 & pi123;
  assign new_n627_ = ~new_n340_ & ~new_n626_;
  assign new_n628_ = ~pi004 & ~pi017;
  assign new_n629_ = pi004 & pi191;
  assign new_n630_ = ~new_n628_ & ~new_n629_;
  assign new_n631_ = ~new_n627_ & new_n630_;
  assign new_n632_ = ~new_n625_ & ~new_n631_;
  assign new_n633_ = new_n621_ & ~new_n624_;
  assign new_n634_ = new_n627_ & ~new_n630_;
  assign new_n635_ = ~new_n633_ & ~new_n634_;
  assign new_n636_ = new_n632_ & new_n635_;
  assign new_n637_ = pi004 & pi124;
  assign new_n638_ = ~new_n327_ & ~new_n637_;
  assign new_n639_ = ~pi004 & ~pi016;
  assign new_n640_ = pi004 & pi190;
  assign new_n641_ = ~new_n639_ & ~new_n640_;
  assign new_n642_ = ~new_n638_ & new_n641_;
  assign new_n643_ = pi004 & pi125;
  assign new_n644_ = ~new_n333_ & ~new_n643_;
  assign new_n645_ = ~pi004 & ~pi015;
  assign new_n646_ = pi004 & pi189;
  assign new_n647_ = ~new_n645_ & ~new_n646_;
  assign new_n648_ = ~new_n644_ & new_n647_;
  assign new_n649_ = ~new_n642_ & ~new_n648_;
  assign new_n650_ = new_n638_ & ~new_n641_;
  assign new_n651_ = new_n644_ & ~new_n647_;
  assign new_n652_ = ~new_n650_ & ~new_n651_;
  assign new_n653_ = new_n649_ & new_n652_;
  assign new_n654_ = new_n636_ & new_n653_;
  assign new_n655_ = ~new_n619_ & new_n654_;
  assign new_n656_ = ~new_n632_ & ~new_n633_;
  assign new_n657_ = ~new_n649_ & ~new_n650_;
  assign new_n658_ = new_n636_ & new_n657_;
  assign new_n659_ = ~new_n656_ & ~new_n658_;
  assign new_n660_ = ~new_n655_ & new_n659_;
  assign new_n661_ = pi004 & pi112;
  assign new_n662_ = ~new_n428_ & ~new_n661_;
  assign new_n663_ = ~pi004 & ~pi023;
  assign new_n664_ = pi004 & pi201;
  assign new_n665_ = ~new_n663_ & ~new_n664_;
  assign new_n666_ = ~new_n662_ & new_n665_;
  assign new_n667_ = pi004 & pi113;
  assign new_n668_ = ~new_n409_ & ~new_n667_;
  assign new_n669_ = ~pi004 & ~pi022;
  assign new_n670_ = pi004 & pi200;
  assign new_n671_ = ~new_n669_ & ~new_n670_;
  assign new_n672_ = ~new_n668_ & new_n671_;
  assign new_n673_ = ~new_n666_ & ~new_n672_;
  assign new_n674_ = new_n662_ & ~new_n665_;
  assign new_n675_ = new_n668_ & ~new_n671_;
  assign new_n676_ = ~new_n674_ & ~new_n675_;
  assign new_n677_ = new_n673_ & new_n676_;
  assign new_n678_ = pi004 & pi111;
  assign new_n679_ = ~new_n422_ & ~new_n678_;
  assign new_n680_ = ~pi004 & ~pi024;
  assign new_n681_ = pi004 & pi202;
  assign new_n682_ = ~new_n680_ & ~new_n681_;
  assign new_n683_ = ~new_n679_ & new_n682_;
  assign new_n684_ = new_n679_ & ~new_n682_;
  assign new_n685_ = ~new_n683_ & ~new_n684_;
  assign new_n686_ = pi004 & pi114;
  assign new_n687_ = ~new_n415_ & ~new_n686_;
  assign new_n688_ = ~pi004 & ~pi037;
  assign new_n689_ = pi004 & pi199;
  assign new_n690_ = ~new_n688_ & ~new_n689_;
  assign new_n691_ = ~new_n687_ & new_n690_;
  assign new_n692_ = new_n687_ & ~new_n690_;
  assign new_n693_ = ~new_n691_ & ~new_n692_;
  assign new_n694_ = new_n685_ & new_n693_;
  assign new_n695_ = new_n677_ & new_n694_;
  assign new_n696_ = pi004 & pi115;
  assign new_n697_ = ~new_n382_ & ~new_n696_;
  assign new_n698_ = ~pi004 & ~pi038;
  assign new_n699_ = pi004 & pi198;
  assign new_n700_ = ~new_n698_ & ~new_n699_;
  assign new_n701_ = ~new_n697_ & new_n700_;
  assign new_n702_ = pi004 & pi118;
  assign new_n703_ = ~new_n362_ & ~new_n702_;
  assign new_n704_ = ~pi004 & ~pi036;
  assign new_n705_ = pi004 & pi195;
  assign new_n706_ = ~new_n704_ & ~new_n705_;
  assign new_n707_ = new_n703_ & ~new_n706_;
  assign new_n708_ = ~new_n701_ & ~new_n707_;
  assign new_n709_ = pi004 & pi117;
  assign new_n710_ = ~new_n373_ & ~new_n709_;
  assign new_n711_ = ~pi004 & ~pi021;
  assign new_n712_ = pi004 & pi196;
  assign new_n713_ = ~new_n711_ & ~new_n712_;
  assign new_n714_ = new_n710_ & ~new_n713_;
  assign new_n715_ = pi004 & pi109;
  assign new_n716_ = ~new_n366_ & ~new_n715_;
  assign new_n717_ = ~pi004 & ~pi035;
  assign new_n718_ = pi004 & pi194;
  assign new_n719_ = ~new_n717_ & ~new_n718_;
  assign new_n720_ = new_n716_ & ~new_n719_;
  assign new_n721_ = ~new_n714_ & ~new_n720_;
  assign new_n722_ = new_n708_ & new_n721_;
  assign new_n723_ = ~new_n716_ & new_n719_;
  assign new_n724_ = ~new_n703_ & new_n706_;
  assign new_n725_ = ~new_n723_ & ~new_n724_;
  assign new_n726_ = new_n697_ & ~new_n700_;
  assign new_n727_ = pi004 & pi116;
  assign new_n728_ = ~new_n388_ & ~new_n727_;
  assign new_n729_ = ~pi004 & ~pi039;
  assign new_n730_ = pi004 & pi197;
  assign new_n731_ = ~new_n729_ & ~new_n730_;
  assign new_n732_ = new_n728_ & ~new_n731_;
  assign new_n733_ = ~new_n726_ & ~new_n732_;
  assign new_n734_ = ~new_n728_ & new_n731_;
  assign new_n735_ = ~new_n710_ & new_n713_;
  assign new_n736_ = ~new_n734_ & ~new_n735_;
  assign new_n737_ = new_n733_ & new_n736_;
  assign new_n738_ = new_n725_ & new_n737_;
  assign new_n739_ = new_n722_ & new_n738_;
  assign new_n740_ = new_n695_ & new_n739_;
  assign new_n741_ = ~new_n660_ & new_n740_;
  assign new_n742_ = ~new_n707_ & ~new_n725_;
  assign new_n743_ = ~new_n735_ & ~new_n742_;
  assign new_n744_ = ~new_n714_ & ~new_n743_;
  assign new_n745_ = ~new_n734_ & ~new_n744_;
  assign new_n746_ = new_n733_ & ~new_n745_;
  assign new_n747_ = ~new_n701_ & ~new_n746_;
  assign new_n748_ = new_n695_ & ~new_n747_;
  assign new_n749_ = new_n685_ & new_n691_;
  assign new_n750_ = new_n677_ & new_n749_;
  assign new_n751_ = ~new_n674_ & ~new_n684_;
  assign new_n752_ = ~new_n673_ & new_n751_;
  assign new_n753_ = ~new_n683_ & ~new_n752_;
  assign new_n754_ = ~new_n750_ & new_n753_;
  assign new_n755_ = ~new_n748_ & new_n754_;
  assign new_n756_ = ~new_n741_ & new_n755_;
  assign new_n757_ = pi004 & ~pi099;
  assign new_n758_ = ~new_n443_ & ~new_n757_;
  assign new_n759_ = pi004 & pi178;
  assign new_n760_ = ~pi004 & ~pi026;
  assign new_n761_ = ~new_n759_ & ~new_n760_;
  assign new_n762_ = ~new_n758_ & ~new_n761_;
  assign new_n763_ = pi004 & pi100;
  assign new_n764_ = ~new_n449_ & ~new_n763_;
  assign new_n765_ = pi004 & pi177;
  assign new_n766_ = ~pi004 & ~pi043;
  assign new_n767_ = ~new_n765_ & ~new_n766_;
  assign new_n768_ = ~new_n764_ & new_n767_;
  assign new_n769_ = ~new_n762_ & ~new_n768_;
  assign new_n770_ = new_n758_ & new_n761_;
  assign new_n771_ = pi004 & pi101;
  assign new_n772_ = ~new_n455_ & ~new_n771_;
  assign new_n773_ = pi004 & pi176;
  assign new_n774_ = ~pi004 & ~pi042;
  assign new_n775_ = ~new_n773_ & ~new_n774_;
  assign new_n776_ = new_n772_ & ~new_n775_;
  assign new_n777_ = ~new_n770_ & ~new_n776_;
  assign new_n778_ = new_n764_ & ~new_n767_;
  assign new_n779_ = ~new_n772_ & new_n775_;
  assign new_n780_ = ~new_n778_ & ~new_n779_;
  assign new_n781_ = new_n777_ & new_n780_;
  assign new_n782_ = new_n769_ & new_n781_;
  assign new_n783_ = pi004 & ~pi095;
  assign new_n784_ = ~new_n443_ & ~new_n783_;
  assign new_n785_ = pi004 & pi182;
  assign new_n786_ = ~pi004 & ~pi054;
  assign new_n787_ = ~new_n785_ & ~new_n786_;
  assign new_n788_ = ~new_n784_ & ~new_n787_;
  assign new_n789_ = new_n784_ & new_n787_;
  assign new_n790_ = ~new_n788_ & ~new_n789_;
  assign new_n791_ = pi004 & ~pi098;
  assign new_n792_ = ~new_n443_ & ~new_n791_;
  assign new_n793_ = pi004 & pi179;
  assign new_n794_ = ~pi004 & ~pi025;
  assign new_n795_ = ~new_n793_ & ~new_n794_;
  assign new_n796_ = new_n792_ & new_n795_;
  assign new_n797_ = ~new_n792_ & ~new_n795_;
  assign new_n798_ = ~new_n796_ & ~new_n797_;
  assign new_n799_ = new_n790_ & new_n798_;
  assign new_n800_ = pi004 & ~pi096;
  assign new_n801_ = ~new_n443_ & ~new_n800_;
  assign new_n802_ = pi004 & pi181;
  assign new_n803_ = ~pi004 & ~pi053;
  assign new_n804_ = ~new_n802_ & ~new_n803_;
  assign new_n805_ = new_n801_ & new_n804_;
  assign new_n806_ = pi004 & ~pi097;
  assign new_n807_ = ~new_n443_ & ~new_n806_;
  assign new_n808_ = pi004 & pi180;
  assign new_n809_ = ~pi004 & ~pi044;
  assign new_n810_ = ~new_n808_ & ~new_n809_;
  assign new_n811_ = new_n807_ & new_n810_;
  assign new_n812_ = ~new_n805_ & ~new_n811_;
  assign new_n813_ = ~new_n801_ & ~new_n804_;
  assign new_n814_ = ~new_n807_ & ~new_n810_;
  assign new_n815_ = ~new_n813_ & ~new_n814_;
  assign new_n816_ = new_n812_ & new_n815_;
  assign new_n817_ = pi004 & pi102;
  assign new_n818_ = ~new_n461_ & ~new_n817_;
  assign new_n819_ = pi004 & pi175;
  assign new_n820_ = ~pi004 & ~pi041;
  assign new_n821_ = ~new_n819_ & ~new_n820_;
  assign new_n822_ = ~new_n818_ & new_n821_;
  assign new_n823_ = new_n818_ & ~new_n821_;
  assign new_n824_ = ~new_n822_ & ~new_n823_;
  assign new_n825_ = pi004 & pi093;
  assign new_n826_ = ~new_n467_ & ~new_n825_;
  assign new_n827_ = pi004 & pi174;
  assign new_n828_ = ~pi004 & ~pi027;
  assign new_n829_ = ~new_n827_ & ~new_n828_;
  assign new_n830_ = ~new_n826_ & new_n829_;
  assign new_n831_ = new_n826_ & ~new_n829_;
  assign new_n832_ = ~new_n830_ & ~new_n831_;
  assign new_n833_ = new_n824_ & new_n832_;
  assign new_n834_ = new_n816_ & new_n833_;
  assign new_n835_ = new_n799_ & new_n834_;
  assign new_n836_ = new_n782_ & new_n835_;
  assign new_n837_ = ~new_n756_ & new_n836_;
  assign new_n838_ = new_n790_ & new_n796_;
  assign new_n839_ = ~new_n823_ & new_n830_;
  assign new_n840_ = ~new_n779_ & ~new_n822_;
  assign new_n841_ = ~new_n839_ & new_n840_;
  assign new_n842_ = ~new_n776_ & ~new_n778_;
  assign new_n843_ = ~new_n841_ & new_n842_;
  assign new_n844_ = ~new_n768_ & ~new_n770_;
  assign new_n845_ = ~new_n843_ & new_n844_;
  assign new_n846_ = ~new_n762_ & new_n799_;
  assign new_n847_ = ~new_n845_ & new_n846_;
  assign new_n848_ = ~new_n838_ & ~new_n847_;
  assign new_n849_ = new_n816_ & ~new_n848_;
  assign new_n850_ = ~new_n788_ & ~new_n813_;
  assign new_n851_ = ~new_n812_ & new_n850_;
  assign new_n852_ = ~new_n789_ & ~new_n851_;
  assign new_n853_ = ~new_n849_ & new_n852_;
  assign new_n854_ = ~new_n837_ & new_n853_;
  assign new_n855_ = pi004 & ~pi089;
  assign new_n856_ = ~new_n443_ & ~new_n855_;
  assign new_n857_ = pi004 & pi168;
  assign new_n858_ = ~pi004 & ~pi056;
  assign new_n859_ = ~new_n857_ & ~new_n858_;
  assign new_n860_ = new_n856_ & new_n859_;
  assign new_n861_ = pi004 & ~pi090;
  assign new_n862_ = ~new_n443_ & ~new_n861_;
  assign new_n863_ = pi004 & pi052;
  assign new_n864_ = ~pi004 & ~pi045;
  assign new_n865_ = ~new_n863_ & ~new_n864_;
  assign new_n866_ = new_n862_ & new_n865_;
  assign new_n867_ = ~new_n860_ & ~new_n866_;
  assign new_n868_ = pi004 & ~pi091;
  assign new_n869_ = ~new_n443_ & ~new_n868_;
  assign new_n870_ = pi004 & pi167;
  assign new_n871_ = ~pi004 & ~pi055;
  assign new_n872_ = ~new_n870_ & ~new_n871_;
  assign new_n873_ = ~new_n869_ & ~new_n872_;
  assign new_n874_ = new_n869_ & new_n872_;
  assign new_n875_ = ~new_n873_ & ~new_n874_;
  assign new_n876_ = ~new_n856_ & ~new_n859_;
  assign new_n877_ = ~new_n862_ & ~new_n865_;
  assign new_n878_ = ~new_n876_ & ~new_n877_;
  assign new_n879_ = new_n875_ & new_n878_;
  assign new_n880_ = new_n867_ & new_n879_;
  assign new_n881_ = pi004 & pi166;
  assign new_n882_ = ~pi004 & ~pi057;
  assign new_n883_ = ~new_n881_ & ~new_n882_;
  assign new_n884_ = ~new_n443_ & new_n883_;
  assign new_n885_ = pi004 & ~pi088;
  assign new_n886_ = ~new_n443_ & ~new_n885_;
  assign new_n887_ = pi004 & pi169;
  assign new_n888_ = ~pi004 & ~pi046;
  assign new_n889_ = ~new_n887_ & ~new_n888_;
  assign new_n890_ = ~new_n886_ & ~new_n889_;
  assign new_n891_ = ~new_n884_ & ~new_n890_;
  assign new_n892_ = new_n886_ & new_n889_;
  assign new_n893_ = new_n443_ & ~new_n883_;
  assign new_n894_ = ~new_n892_ & ~new_n893_;
  assign new_n895_ = new_n891_ & new_n894_;
  assign new_n896_ = new_n880_ & new_n895_;
  assign new_n897_ = ~new_n854_ & new_n896_;
  assign new_n898_ = new_n880_ & new_n884_;
  assign new_n899_ = new_n874_ & ~new_n877_;
  assign new_n900_ = new_n867_ & ~new_n899_;
  assign new_n901_ = ~new_n876_ & ~new_n900_;
  assign new_n902_ = ~new_n898_ & ~new_n901_;
  assign new_n903_ = ~new_n890_ & ~new_n902_;
  assign new_n904_ = ~pi164 & ~pi172;
  assign new_n905_ = pi204 & new_n904_;
  assign new_n906_ = pi010 & ~new_n905_;
  assign new_n907_ = ~new_n892_ & ~new_n906_;
  assign new_n908_ = ~new_n903_ & new_n907_;
  assign new_n909_ = ~new_n897_ & new_n908_;
  assign new_n910_ = pi164 & pi172;
  assign new_n911_ = ~pi010 & pi204;
  assign new_n912_ = ~new_n910_ & new_n911_;
  assign po10 = ~new_n909_ & ~new_n912_;
  assign new_n914_ = ~new_n292_ & ~new_n316_;
  assign new_n915_ = new_n318_ & new_n319_;
  assign new_n916_ = new_n320_ & new_n915_;
  assign new_n917_ = ~new_n314_ & ~new_n916_;
  assign new_n918_ = new_n914_ & ~new_n917_;
  assign new_n919_ = ~new_n914_ & new_n917_;
  assign po11 = ~new_n918_ & ~new_n919_;
  assign new_n921_ = ~new_n312_ & ~new_n915_;
  assign new_n922_ = new_n320_ & ~new_n921_;
  assign new_n923_ = ~new_n320_ & new_n921_;
  assign po12 = ~new_n922_ & ~new_n923_;
  assign new_n925_ = ~new_n305_ & ~new_n308_;
  assign new_n926_ = ~new_n318_ & new_n925_;
  assign new_n927_ = new_n319_ & ~new_n926_;
  assign new_n928_ = ~new_n319_ & new_n926_;
  assign po13 = ~new_n927_ & ~new_n928_;
  assign new_n930_ = ~new_n277_ & ~new_n283_;
  assign new_n931_ = new_n307_ & ~new_n930_;
  assign new_n932_ = ~new_n307_ & new_n930_;
  assign po14 = ~new_n931_ & ~new_n932_;
  assign new_n934_ = ~new_n325_ & new_n338_;
  assign new_n935_ = new_n355_ & ~new_n934_;
  assign new_n936_ = ~new_n343_ & ~new_n935_;
  assign new_n937_ = ~new_n342_ & ~new_n936_;
  assign new_n938_ = new_n350_ & ~new_n937_;
  assign new_n939_ = ~new_n350_ & new_n937_;
  assign po15 = ~new_n938_ & ~new_n939_;
  assign new_n941_ = new_n344_ & ~new_n935_;
  assign new_n942_ = ~new_n344_ & new_n935_;
  assign po16 = ~new_n941_ & ~new_n942_;
  assign new_n944_ = ~new_n325_ & ~new_n336_;
  assign new_n945_ = ~new_n335_ & ~new_n944_;
  assign new_n946_ = new_n331_ & ~new_n945_;
  assign new_n947_ = ~new_n331_ & new_n945_;
  assign po17 = ~new_n946_ & ~new_n947_;
  assign new_n949_ = ~new_n325_ & new_n337_;
  assign new_n950_ = new_n325_ & ~new_n337_;
  assign po18 = ~new_n949_ & ~new_n950_;
  assign new_n952_ = new_n451_ & ~new_n457_;
  assign new_n953_ = ~new_n451_ & new_n457_;
  assign new_n954_ = ~new_n952_ & ~new_n953_;
  assign new_n955_ = ~pi004 & pi069;
  assign new_n956_ = pi004 & pi083;
  assign new_n957_ = ~new_n955_ & ~new_n956_;
  assign new_n958_ = new_n445_ & ~new_n469_;
  assign new_n959_ = ~new_n445_ & new_n469_;
  assign new_n960_ = ~new_n958_ & ~new_n959_;
  assign new_n961_ = new_n957_ & new_n960_;
  assign new_n962_ = ~new_n957_ & ~new_n960_;
  assign new_n963_ = ~new_n961_ & ~new_n962_;
  assign new_n964_ = new_n477_ & new_n483_;
  assign new_n965_ = new_n478_ & new_n482_;
  assign new_n966_ = ~new_n964_ & ~new_n965_;
  assign new_n967_ = new_n489_ & new_n493_;
  assign new_n968_ = new_n488_ & new_n494_;
  assign new_n969_ = ~new_n967_ & ~new_n968_;
  assign new_n970_ = ~new_n966_ & new_n969_;
  assign new_n971_ = new_n966_ & ~new_n969_;
  assign new_n972_ = ~new_n970_ & ~new_n971_;
  assign new_n973_ = new_n463_ & ~new_n972_;
  assign new_n974_ = ~new_n463_ & new_n972_;
  assign new_n975_ = ~new_n973_ & ~new_n974_;
  assign new_n976_ = ~new_n963_ & new_n975_;
  assign new_n977_ = new_n963_ & ~new_n975_;
  assign new_n978_ = ~new_n976_ & ~new_n977_;
  assign new_n979_ = new_n954_ & ~new_n978_;
  assign new_n980_ = ~new_n954_ & new_n978_;
  assign new_n981_ = ~new_n979_ & ~new_n980_;
  assign new_n982_ = pi004 & ~new_n443_;
  assign new_n983_ = pi133 & pi134;
  assign new_n984_ = ~pi133 & ~pi134;
  assign new_n985_ = ~new_n983_ & ~new_n984_;
  assign new_n986_ = new_n982_ & new_n985_;
  assign new_n987_ = ~new_n443_ & new_n522_;
  assign new_n988_ = new_n536_ & new_n542_;
  assign new_n989_ = new_n537_ & new_n541_;
  assign new_n990_ = ~new_n988_ & ~new_n989_;
  assign new_n991_ = new_n520_ & new_n528_;
  assign new_n992_ = new_n519_ & new_n529_;
  assign new_n993_ = ~new_n991_ & ~new_n992_;
  assign new_n994_ = new_n990_ & ~new_n993_;
  assign new_n995_ = ~new_n990_ & new_n993_;
  assign new_n996_ = ~new_n994_ & ~new_n995_;
  assign new_n997_ = new_n987_ & ~new_n996_;
  assign new_n998_ = ~new_n987_ & new_n996_;
  assign new_n999_ = ~new_n997_ & ~new_n998_;
  assign new_n1000_ = new_n986_ & new_n999_;
  assign new_n1001_ = ~new_n986_ & ~new_n999_;
  assign new_n1002_ = ~new_n1000_ & ~new_n1001_;
  assign new_n1003_ = ~new_n410_ & new_n423_;
  assign new_n1004_ = new_n410_ & ~new_n423_;
  assign new_n1005_ = ~new_n1003_ & ~new_n1004_;
  assign new_n1006_ = new_n416_ & ~new_n429_;
  assign new_n1007_ = ~new_n416_ & new_n429_;
  assign new_n1008_ = ~new_n1006_ & ~new_n1007_;
  assign new_n1009_ = new_n1005_ & new_n1008_;
  assign new_n1010_ = ~new_n1005_ & ~new_n1008_;
  assign new_n1011_ = ~new_n1009_ & ~new_n1010_;
  assign new_n1012_ = new_n363_ & ~new_n1011_;
  assign new_n1013_ = ~new_n363_ & new_n1011_;
  assign new_n1014_ = ~new_n1012_ & ~new_n1013_;
  assign new_n1015_ = ~new_n367_ & new_n383_;
  assign new_n1016_ = new_n367_ & ~new_n383_;
  assign new_n1017_ = ~new_n1015_ & ~new_n1016_;
  assign new_n1018_ = new_n389_ & new_n1017_;
  assign new_n1019_ = ~new_n389_ & ~new_n1017_;
  assign new_n1020_ = ~new_n1018_ & ~new_n1019_;
  assign new_n1021_ = pi004 & pi149;
  assign new_n1022_ = ~pi004 & pi059;
  assign new_n1023_ = ~new_n1021_ & ~new_n1022_;
  assign new_n1024_ = new_n374_ & ~new_n1023_;
  assign new_n1025_ = ~new_n374_ & new_n1023_;
  assign new_n1026_ = ~new_n1024_ & ~new_n1025_;
  assign new_n1027_ = new_n1020_ & ~new_n1026_;
  assign new_n1028_ = ~new_n1020_ & new_n1026_;
  assign new_n1029_ = ~new_n1027_ & ~new_n1028_;
  assign new_n1030_ = new_n1014_ & new_n1029_;
  assign new_n1031_ = ~new_n1014_ & ~new_n1029_;
  assign new_n1032_ = ~new_n1030_ & ~new_n1031_;
  assign new_n1033_ = new_n328_ & ~new_n347_;
  assign new_n1034_ = ~new_n328_ & new_n347_;
  assign new_n1035_ = ~new_n1033_ & ~new_n1034_;
  assign new_n1036_ = new_n334_ & ~new_n341_;
  assign new_n1037_ = ~new_n334_ & new_n341_;
  assign new_n1038_ = ~new_n1036_ & ~new_n1037_;
  assign new_n1039_ = new_n1035_ & new_n1038_;
  assign new_n1040_ = ~new_n1035_ & ~new_n1038_;
  assign new_n1041_ = ~new_n1039_ & ~new_n1040_;
  assign new_n1042_ = new_n295_ & ~new_n1041_;
  assign new_n1043_ = ~new_n295_ & new_n1041_;
  assign new_n1044_ = ~new_n1042_ & ~new_n1043_;
  assign new_n1045_ = pi004 & pi161;
  assign new_n1046_ = ~pi004 & pi012;
  assign new_n1047_ = ~new_n1045_ & ~new_n1046_;
  assign new_n1048_ = new_n300_ & ~new_n1047_;
  assign new_n1049_ = ~new_n300_ & new_n1047_;
  assign new_n1050_ = ~new_n1048_ & ~new_n1049_;
  assign new_n1051_ = new_n304_ & new_n1050_;
  assign new_n1052_ = ~new_n304_ & ~new_n1050_;
  assign new_n1053_ = ~new_n1051_ & ~new_n1052_;
  assign new_n1054_ = new_n279_ & ~new_n291_;
  assign new_n1055_ = ~new_n279_ & new_n291_;
  assign new_n1056_ = ~new_n1054_ & ~new_n1055_;
  assign new_n1057_ = new_n1053_ & ~new_n1056_;
  assign new_n1058_ = ~new_n1053_ & new_n1056_;
  assign new_n1059_ = ~new_n1057_ & ~new_n1058_;
  assign new_n1060_ = new_n1044_ & new_n1059_;
  assign new_n1061_ = ~new_n1044_ & ~new_n1059_;
  assign new_n1062_ = ~new_n1060_ & ~new_n1061_;
  assign new_n1063_ = new_n1032_ & new_n1062_;
  assign new_n1064_ = ~new_n1002_ & new_n1063_;
  assign po19 = new_n981_ | ~new_n1064_;
  assign new_n1066_ = ~pi004 & pi030;
  assign new_n1067_ = pi004 & ~pi184;
  assign new_n1068_ = ~new_n1066_ & ~new_n1067_;
  assign new_n1069_ = new_n581_ & ~new_n587_;
  assign new_n1070_ = ~new_n581_ & new_n587_;
  assign new_n1071_ = ~new_n1069_ & ~new_n1070_;
  assign new_n1072_ = new_n1068_ & new_n1071_;
  assign new_n1073_ = ~new_n1068_ & ~new_n1071_;
  assign new_n1074_ = ~new_n1072_ & ~new_n1073_;
  assign new_n1075_ = pi004 & ~pi183;
  assign new_n1076_ = ~pi004 & pi029;
  assign new_n1077_ = ~new_n1075_ & ~new_n1076_;
  assign new_n1078_ = ~new_n575_ & ~new_n602_;
  assign new_n1079_ = new_n575_ & new_n602_;
  assign new_n1080_ = ~new_n1078_ & ~new_n1079_;
  assign new_n1081_ = ~new_n624_ & new_n641_;
  assign new_n1082_ = new_n624_ & ~new_n641_;
  assign new_n1083_ = ~new_n1081_ & ~new_n1082_;
  assign new_n1084_ = ~new_n630_ & new_n647_;
  assign new_n1085_ = new_n630_ & ~new_n647_;
  assign new_n1086_ = ~new_n1084_ & ~new_n1085_;
  assign new_n1087_ = new_n1083_ & new_n1086_;
  assign new_n1088_ = ~new_n1083_ & ~new_n1086_;
  assign new_n1089_ = ~new_n1087_ & ~new_n1088_;
  assign new_n1090_ = new_n1080_ & ~new_n1089_;
  assign new_n1091_ = ~new_n1080_ & new_n1089_;
  assign new_n1092_ = ~new_n1090_ & ~new_n1091_;
  assign new_n1093_ = new_n1077_ & new_n1092_;
  assign new_n1094_ = ~new_n1077_ & ~new_n1092_;
  assign new_n1095_ = ~new_n1093_ & ~new_n1094_;
  assign new_n1096_ = ~new_n1074_ & ~new_n1095_;
  assign new_n1097_ = ~new_n883_ & new_n889_;
  assign new_n1098_ = new_n883_ & ~new_n889_;
  assign new_n1099_ = ~new_n1097_ & ~new_n1098_;
  assign new_n1100_ = new_n859_ & new_n1099_;
  assign new_n1101_ = ~new_n859_ & ~new_n1099_;
  assign new_n1102_ = ~new_n1100_ & ~new_n1101_;
  assign new_n1103_ = ~new_n865_ & ~new_n872_;
  assign new_n1104_ = new_n865_ & new_n872_;
  assign new_n1105_ = ~new_n1103_ & ~new_n1104_;
  assign new_n1106_ = pi004 & ~pi165;
  assign new_n1107_ = ~pi004 & pi058;
  assign new_n1108_ = ~new_n1106_ & ~new_n1107_;
  assign new_n1109_ = new_n1105_ & ~new_n1108_;
  assign new_n1110_ = ~new_n1105_ & new_n1108_;
  assign new_n1111_ = ~new_n1109_ & ~new_n1110_;
  assign new_n1112_ = ~pi170 & ~pi171;
  assign new_n1113_ = pi170 & pi171;
  assign new_n1114_ = ~new_n1112_ & ~new_n1113_;
  assign new_n1115_ = pi004 & ~new_n1114_;
  assign new_n1116_ = ~new_n904_ & ~new_n910_;
  assign new_n1117_ = ~pi004 & ~new_n1116_;
  assign new_n1118_ = ~new_n1115_ & ~new_n1117_;
  assign new_n1119_ = ~new_n1111_ & new_n1118_;
  assign new_n1120_ = new_n1111_ & ~new_n1118_;
  assign new_n1121_ = ~new_n1119_ & ~new_n1120_;
  assign new_n1122_ = ~new_n1102_ & new_n1121_;
  assign new_n1123_ = new_n1102_ & ~new_n1121_;
  assign new_n1124_ = ~new_n1122_ & ~new_n1123_;
  assign new_n1125_ = ~new_n775_ & ~new_n821_;
  assign new_n1126_ = new_n775_ & new_n821_;
  assign new_n1127_ = ~new_n1125_ & ~new_n1126_;
  assign new_n1128_ = new_n804_ & ~new_n810_;
  assign new_n1129_ = ~new_n804_ & new_n810_;
  assign new_n1130_ = ~new_n1128_ & ~new_n1129_;
  assign new_n1131_ = new_n787_ & ~new_n795_;
  assign new_n1132_ = ~new_n787_ & new_n795_;
  assign new_n1133_ = ~new_n1131_ & ~new_n1132_;
  assign new_n1134_ = new_n1130_ & new_n1133_;
  assign new_n1135_ = ~new_n1130_ & ~new_n1133_;
  assign new_n1136_ = ~new_n1134_ & ~new_n1135_;
  assign new_n1137_ = new_n1127_ & ~new_n1136_;
  assign new_n1138_ = ~new_n1127_ & new_n1136_;
  assign new_n1139_ = ~new_n1137_ & ~new_n1138_;
  assign new_n1140_ = new_n761_ & ~new_n829_;
  assign new_n1141_ = ~new_n761_ & new_n829_;
  assign new_n1142_ = ~new_n1140_ & ~new_n1141_;
  assign new_n1143_ = new_n767_ & new_n1142_;
  assign new_n1144_ = ~new_n767_ & ~new_n1142_;
  assign new_n1145_ = ~new_n1143_ & ~new_n1144_;
  assign new_n1146_ = pi004 & ~pi173;
  assign new_n1147_ = ~pi004 & pi040;
  assign new_n1148_ = ~new_n1146_ & ~new_n1147_;
  assign new_n1149_ = new_n1145_ & ~new_n1148_;
  assign new_n1150_ = ~new_n1145_ & new_n1148_;
  assign new_n1151_ = ~new_n1149_ & ~new_n1150_;
  assign new_n1152_ = new_n1139_ & new_n1151_;
  assign new_n1153_ = ~new_n1139_ & ~new_n1151_;
  assign new_n1154_ = ~new_n1152_ & ~new_n1153_;
  assign new_n1155_ = ~new_n1124_ & new_n1154_;
  assign new_n1156_ = ~new_n1096_ & new_n1155_;
  assign new_n1157_ = new_n1074_ & new_n1095_;
  assign new_n1158_ = new_n700_ & ~new_n719_;
  assign new_n1159_ = ~new_n700_ & new_n719_;
  assign new_n1160_ = ~new_n1158_ & ~new_n1159_;
  assign new_n1161_ = new_n731_ & new_n1160_;
  assign new_n1162_ = ~new_n731_ & ~new_n1160_;
  assign new_n1163_ = ~new_n1161_ & ~new_n1162_;
  assign new_n1164_ = pi004 & ~pi193;
  assign new_n1165_ = ~pi004 & pi020;
  assign new_n1166_ = ~new_n1164_ & ~new_n1165_;
  assign new_n1167_ = ~new_n706_ & ~new_n713_;
  assign new_n1168_ = new_n706_ & new_n713_;
  assign new_n1169_ = ~new_n1167_ & ~new_n1168_;
  assign new_n1170_ = new_n665_ & ~new_n671_;
  assign new_n1171_ = ~new_n665_ & new_n671_;
  assign new_n1172_ = ~new_n1170_ & ~new_n1171_;
  assign new_n1173_ = new_n682_ & ~new_n690_;
  assign new_n1174_ = ~new_n682_ & new_n690_;
  assign new_n1175_ = ~new_n1173_ & ~new_n1174_;
  assign new_n1176_ = new_n1172_ & new_n1175_;
  assign new_n1177_ = ~new_n1172_ & ~new_n1175_;
  assign new_n1178_ = ~new_n1176_ & ~new_n1177_;
  assign new_n1179_ = new_n1169_ & ~new_n1178_;
  assign new_n1180_ = ~new_n1169_ & new_n1178_;
  assign new_n1181_ = ~new_n1179_ & ~new_n1180_;
  assign new_n1182_ = new_n1166_ & new_n1181_;
  assign new_n1183_ = ~new_n1166_ & ~new_n1181_;
  assign new_n1184_ = ~new_n1182_ & ~new_n1183_;
  assign new_n1185_ = ~new_n1163_ & new_n1184_;
  assign new_n1186_ = new_n1163_ & ~new_n1184_;
  assign new_n1187_ = ~new_n1185_ & ~new_n1186_;
  assign new_n1188_ = ~new_n1157_ & new_n1187_;
  assign po20 = ~new_n1156_ | ~new_n1188_;
  assign new_n1190_ = pi004 & ~pi092;
  assign new_n1191_ = ~new_n885_ & ~new_n1190_;
  assign new_n1192_ = new_n885_ & new_n1190_;
  assign new_n1193_ = ~new_n1191_ & ~new_n1192_;
  assign new_n1194_ = ~new_n855_ & ~new_n1193_;
  assign new_n1195_ = new_n855_ & new_n1193_;
  assign new_n1196_ = ~new_n443_ & ~new_n1195_;
  assign new_n1197_ = ~new_n1194_ & new_n1196_;
  assign new_n1198_ = new_n861_ & new_n869_;
  assign new_n1199_ = new_n862_ & new_n868_;
  assign new_n1200_ = ~new_n1198_ & ~new_n1199_;
  assign new_n1201_ = pi086 & pi087;
  assign new_n1202_ = ~pi086 & ~pi087;
  assign new_n1203_ = ~new_n1201_ & ~new_n1202_;
  assign new_n1204_ = new_n982_ & new_n1203_;
  assign new_n1205_ = ~new_n1200_ & ~new_n1204_;
  assign new_n1206_ = new_n1200_ & new_n1204_;
  assign new_n1207_ = ~new_n1205_ & ~new_n1206_;
  assign new_n1208_ = new_n1197_ & ~new_n1207_;
  assign new_n1209_ = ~new_n1197_ & new_n1207_;
  assign new_n1210_ = ~new_n1208_ & ~new_n1209_;
  assign new_n1211_ = new_n662_ & ~new_n668_;
  assign new_n1212_ = ~new_n662_ & new_n668_;
  assign new_n1213_ = ~new_n1211_ & ~new_n1212_;
  assign new_n1214_ = new_n679_ & ~new_n687_;
  assign new_n1215_ = ~new_n679_ & new_n687_;
  assign new_n1216_ = ~new_n1214_ & ~new_n1215_;
  assign new_n1217_ = new_n1213_ & new_n1216_;
  assign new_n1218_ = ~new_n1213_ & ~new_n1216_;
  assign new_n1219_ = ~new_n1217_ & ~new_n1218_;
  assign new_n1220_ = new_n703_ & ~new_n1219_;
  assign new_n1221_ = ~new_n703_ & new_n1219_;
  assign new_n1222_ = ~new_n1220_ & ~new_n1221_;
  assign new_n1223_ = new_n697_ & ~new_n716_;
  assign new_n1224_ = ~new_n697_ & new_n716_;
  assign new_n1225_ = ~new_n1223_ & ~new_n1224_;
  assign new_n1226_ = new_n728_ & new_n1225_;
  assign new_n1227_ = ~new_n728_ & ~new_n1225_;
  assign new_n1228_ = ~new_n1226_ & ~new_n1227_;
  assign new_n1229_ = pi004 & pi119;
  assign new_n1230_ = ~new_n1022_ & ~new_n1229_;
  assign new_n1231_ = new_n710_ & ~new_n1230_;
  assign new_n1232_ = ~new_n710_ & new_n1230_;
  assign new_n1233_ = ~new_n1231_ & ~new_n1232_;
  assign new_n1234_ = new_n1228_ & ~new_n1233_;
  assign new_n1235_ = ~new_n1228_ & new_n1233_;
  assign new_n1236_ = ~new_n1234_ & ~new_n1235_;
  assign new_n1237_ = new_n1222_ & new_n1236_;
  assign new_n1238_ = ~new_n1210_ & ~new_n1237_;
  assign new_n1239_ = ~new_n621_ & new_n638_;
  assign new_n1240_ = new_n621_ & ~new_n638_;
  assign new_n1241_ = ~new_n1239_ & ~new_n1240_;
  assign new_n1242_ = ~new_n627_ & new_n644_;
  assign new_n1243_ = new_n627_ & ~new_n644_;
  assign new_n1244_ = ~new_n1242_ & ~new_n1243_;
  assign new_n1245_ = new_n1241_ & new_n1244_;
  assign new_n1246_ = ~new_n1241_ & ~new_n1244_;
  assign new_n1247_ = ~new_n1245_ & ~new_n1246_;
  assign new_n1248_ = new_n572_ & ~new_n1247_;
  assign new_n1249_ = ~new_n572_ & new_n1247_;
  assign new_n1250_ = ~new_n1248_ & ~new_n1249_;
  assign new_n1251_ = pi004 & pi130;
  assign new_n1252_ = ~new_n1046_ & ~new_n1251_;
  assign new_n1253_ = new_n578_ & ~new_n1252_;
  assign new_n1254_ = ~new_n578_ & new_n1252_;
  assign new_n1255_ = ~new_n1253_ & ~new_n1254_;
  assign new_n1256_ = new_n584_ & new_n1255_;
  assign new_n1257_ = ~new_n584_ & ~new_n1255_;
  assign new_n1258_ = ~new_n1256_ & ~new_n1257_;
  assign new_n1259_ = pi004 & pi120;
  assign new_n1260_ = ~new_n276_ & ~new_n1259_;
  assign new_n1261_ = new_n599_ & ~new_n1260_;
  assign new_n1262_ = ~new_n599_ & new_n1260_;
  assign new_n1263_ = ~new_n1261_ & ~new_n1262_;
  assign new_n1264_ = new_n1258_ & ~new_n1263_;
  assign new_n1265_ = ~new_n1258_ & new_n1263_;
  assign new_n1266_ = ~new_n1264_ & ~new_n1265_;
  assign new_n1267_ = ~new_n1250_ & ~new_n1266_;
  assign new_n1268_ = ~new_n1222_ & ~new_n1236_;
  assign new_n1269_ = new_n1250_ & new_n1266_;
  assign new_n1270_ = ~new_n1268_ & ~new_n1269_;
  assign new_n1271_ = ~new_n1267_ & new_n1270_;
  assign new_n1272_ = new_n1238_ & new_n1271_;
  assign new_n1273_ = pi004 & pi103;
  assign new_n1274_ = ~new_n955_ & ~new_n1273_;
  assign new_n1275_ = new_n764_ & ~new_n826_;
  assign new_n1276_ = ~new_n764_ & new_n826_;
  assign new_n1277_ = ~new_n1275_ & ~new_n1276_;
  assign new_n1278_ = new_n1274_ & new_n1277_;
  assign new_n1279_ = ~new_n1274_ & ~new_n1277_;
  assign new_n1280_ = ~new_n1278_ & ~new_n1279_;
  assign new_n1281_ = new_n758_ & ~new_n772_;
  assign new_n1282_ = ~new_n758_ & new_n772_;
  assign new_n1283_ = ~new_n1281_ & ~new_n1282_;
  assign new_n1284_ = new_n792_ & new_n806_;
  assign new_n1285_ = new_n791_ & new_n807_;
  assign new_n1286_ = ~new_n1284_ & ~new_n1285_;
  assign new_n1287_ = new_n783_ & new_n801_;
  assign new_n1288_ = new_n784_ & new_n800_;
  assign new_n1289_ = ~new_n1287_ & ~new_n1288_;
  assign new_n1290_ = ~new_n1286_ & new_n1289_;
  assign new_n1291_ = new_n1286_ & ~new_n1289_;
  assign new_n1292_ = ~new_n1290_ & ~new_n1291_;
  assign new_n1293_ = new_n818_ & ~new_n1292_;
  assign new_n1294_ = ~new_n818_ & new_n1292_;
  assign new_n1295_ = ~new_n1293_ & ~new_n1294_;
  assign new_n1296_ = new_n1283_ & new_n1295_;
  assign new_n1297_ = ~new_n1283_ & ~new_n1295_;
  assign new_n1298_ = ~new_n1296_ & ~new_n1297_;
  assign new_n1299_ = new_n1280_ & ~new_n1298_;
  assign new_n1300_ = ~new_n1280_ & new_n1298_;
  assign new_n1301_ = ~new_n1299_ & ~new_n1300_;
  assign po21 = ~new_n1272_ | ~new_n1301_;
  assign new_n1303_ = ~new_n442_ & new_n472_;
  assign new_n1304_ = new_n442_ & ~new_n472_;
  assign po22 = ~new_n1303_ & ~new_n1304_;
  assign new_n1306_ = ~new_n518_ & new_n526_;
  assign new_n1307_ = new_n518_ & ~new_n526_;
  assign po23 = ~new_n1306_ & ~new_n1307_;
  assign new_n1309_ = ~new_n660_ & new_n739_;
  assign new_n1310_ = new_n747_ & ~new_n1309_;
  assign new_n1311_ = new_n695_ & ~new_n1310_;
  assign po24 = ~new_n754_ | new_n1311_;
  assign new_n1313_ = ~new_n475_ & new_n507_;
  assign new_n1314_ = new_n442_ & new_n507_;
  assign new_n1315_ = ~new_n1313_ & ~new_n1314_;
  assign new_n1316_ = new_n448_ & ~new_n1315_;
  assign new_n1317_ = ~new_n448_ & new_n1315_;
  assign po25 = new_n1316_ | new_n1317_;
  assign new_n1319_ = ~new_n442_ & new_n473_;
  assign new_n1320_ = new_n460_ & new_n1319_;
  assign new_n1321_ = ~new_n505_ & ~new_n1320_;
  assign new_n1322_ = new_n454_ & ~new_n1321_;
  assign new_n1323_ = ~new_n454_ & new_n1321_;
  assign po26 = ~new_n1322_ & ~new_n1323_;
  assign new_n1325_ = ~new_n464_ & ~new_n502_;
  assign new_n1326_ = ~new_n1319_ & new_n1325_;
  assign new_n1327_ = new_n460_ & ~new_n1326_;
  assign new_n1328_ = ~new_n460_ & new_n1326_;
  assign po27 = ~new_n1327_ & ~new_n1328_;
  assign new_n1330_ = ~new_n470_ & ~new_n1303_;
  assign new_n1331_ = new_n466_ & ~new_n1330_;
  assign new_n1332_ = ~new_n466_ & new_n1330_;
  assign po28 = ~new_n1331_ & ~new_n1332_;
  assign new_n1334_ = new_n552_ & ~new_n554_;
  assign new_n1335_ = ~new_n544_ & ~new_n1334_;
  assign new_n1336_ = ~new_n543_ & ~new_n1335_;
  assign new_n1337_ = ~new_n518_ & new_n535_;
  assign new_n1338_ = new_n545_ & new_n1337_;
  assign new_n1339_ = new_n1336_ & ~new_n1338_;
  assign new_n1340_ = new_n540_ & new_n1339_;
  assign new_n1341_ = ~new_n540_ & ~new_n1339_;
  assign po29 = new_n1340_ | new_n1341_;
  assign new_n1343_ = new_n1334_ & ~new_n1337_;
  assign new_n1344_ = new_n545_ & new_n1343_;
  assign new_n1345_ = ~new_n545_ & ~new_n1343_;
  assign po30 = new_n1344_ | new_n1345_;
  assign new_n1347_ = ~new_n524_ & ~new_n1306_;
  assign new_n1348_ = new_n549_ & ~new_n1347_;
  assign new_n1349_ = ~new_n533_ & ~new_n1348_;
  assign new_n1350_ = new_n532_ & new_n1349_;
  assign new_n1351_ = ~new_n532_ & ~new_n1349_;
  assign po31 = new_n1350_ | new_n1351_;
  assign new_n1353_ = ~new_n549_ & new_n1347_;
  assign po32 = ~new_n1348_ & ~new_n1353_;
  assign new_n1355_ = ~po01 & ~po02;
  assign new_n1356_ = ~po03 & ~po04;
  assign new_n1357_ = new_n1355_ & new_n1356_;
  assign new_n1358_ = ~po19 & new_n1357_;
  assign new_n1359_ = ~po21 & new_n1358_;
  assign po33 = po20 | ~new_n1359_;
  assign new_n1361_ = ~new_n442_ & new_n476_;
  assign new_n1362_ = new_n509_ & ~new_n1361_;
  assign new_n1363_ = new_n487_ & ~new_n1362_;
  assign new_n1364_ = ~new_n491_ & new_n1363_;
  assign new_n1365_ = ~new_n514_ & ~new_n1364_;
  assign new_n1366_ = new_n497_ & ~new_n1365_;
  assign new_n1367_ = ~new_n497_ & new_n1365_;
  assign po34 = ~new_n1366_ & ~new_n1367_;
  assign new_n1369_ = new_n512_ & ~new_n1363_;
  assign new_n1370_ = new_n492_ & ~new_n1369_;
  assign new_n1371_ = ~new_n492_ & new_n1369_;
  assign po35 = ~new_n1370_ & ~new_n1371_;
  assign new_n1373_ = ~new_n485_ & ~new_n1362_;
  assign new_n1374_ = ~new_n484_ & ~new_n1373_;
  assign new_n1375_ = new_n481_ & ~new_n1374_;
  assign new_n1376_ = ~new_n481_ & new_n1374_;
  assign po36 = ~new_n1375_ & ~new_n1376_;
  assign new_n1378_ = new_n486_ & ~new_n1362_;
  assign new_n1379_ = ~new_n486_ & new_n1362_;
  assign po37 = ~new_n1378_ & ~new_n1379_;
  assign new_n1381_ = ~new_n360_ & new_n370_;
  assign new_n1382_ = new_n360_ & ~new_n370_;
  assign po38 = ~new_n1381_ & ~new_n1382_;
  assign new_n1384_ = new_n560_ & ~new_n562_;
  assign new_n1385_ = ~new_n563_ & ~new_n1384_;
  assign new_n1386_ = ~new_n567_ & ~new_n1385_;
  assign new_n1387_ = new_n567_ & new_n1385_;
  assign po39 = new_n1386_ | new_n1387_;
  assign new_n1389_ = ~new_n560_ & ~new_n564_;
  assign new_n1390_ = new_n560_ & new_n564_;
  assign po40 = new_n1389_ | new_n1390_;
  assign new_n1392_ = new_n399_ & ~new_n401_;
  assign new_n1393_ = ~new_n391_ & ~new_n1392_;
  assign new_n1394_ = ~new_n390_ & ~new_n1393_;
  assign new_n1395_ = ~new_n360_ & new_n380_;
  assign new_n1396_ = new_n392_ & new_n1395_;
  assign new_n1397_ = new_n1394_ & ~new_n1396_;
  assign new_n1398_ = new_n386_ & ~new_n1397_;
  assign new_n1399_ = ~new_n386_ & new_n1397_;
  assign po41 = ~new_n1398_ & ~new_n1399_;
  assign new_n1401_ = new_n1392_ & ~new_n1395_;
  assign new_n1402_ = new_n392_ & ~new_n1401_;
  assign new_n1403_ = ~new_n392_ & new_n1401_;
  assign po42 = ~new_n1402_ & ~new_n1403_;
  assign new_n1405_ = ~new_n368_ & ~new_n1381_;
  assign new_n1406_ = new_n396_ & ~new_n1405_;
  assign new_n1407_ = ~new_n378_ & ~new_n1406_;
  assign new_n1408_ = new_n377_ & ~new_n1407_;
  assign new_n1409_ = ~new_n377_ & new_n1407_;
  assign po43 = ~new_n1408_ & ~new_n1409_;
  assign new_n1411_ = ~new_n396_ & new_n1405_;
  assign po44 = ~new_n1406_ & ~new_n1411_;
  assign new_n1413_ = ~new_n407_ & new_n420_;
  assign new_n1414_ = ~new_n430_ & new_n1413_;
  assign new_n1415_ = new_n439_ & ~new_n1414_;
  assign new_n1416_ = new_n426_ & ~new_n1415_;
  assign new_n1417_ = ~new_n426_ & new_n1415_;
  assign po45 = ~new_n1416_ & ~new_n1417_;
  assign new_n1419_ = new_n437_ & ~new_n1413_;
  assign new_n1420_ = new_n432_ & ~new_n1419_;
  assign new_n1421_ = ~new_n432_ & new_n1419_;
  assign po46 = ~new_n1420_ & ~new_n1421_;
  assign new_n1423_ = ~new_n407_ & ~new_n418_;
  assign new_n1424_ = ~new_n417_ & ~new_n1423_;
  assign new_n1425_ = new_n413_ & ~new_n1424_;
  assign new_n1426_ = ~new_n413_ & new_n1424_;
  assign po47 = ~new_n1425_ & ~new_n1426_;
  assign new_n1428_ = ~new_n407_ & new_n419_;
  assign new_n1429_ = new_n407_ & ~new_n419_;
  assign po48 = ~new_n1428_ & ~new_n1429_;
  assign new_n1431_ = ~new_n465_ & ~new_n470_;
  assign new_n1432_ = ~new_n464_ & ~new_n1431_;
  assign new_n1433_ = new_n507_ & ~new_n1432_;
  assign new_n1434_ = ~new_n507_ & new_n1432_;
  assign new_n1435_ = ~new_n1433_ & ~new_n1434_;
  assign new_n1436_ = new_n448_ & ~new_n1435_;
  assign new_n1437_ = ~new_n448_ & new_n1435_;
  assign new_n1438_ = ~new_n1436_ & ~new_n1437_;
  assign new_n1439_ = new_n454_ & ~new_n460_;
  assign new_n1440_ = ~new_n454_ & new_n460_;
  assign new_n1441_ = ~new_n1439_ & ~new_n1440_;
  assign new_n1442_ = new_n470_ & ~new_n505_;
  assign new_n1443_ = ~new_n459_ & ~new_n470_;
  assign new_n1444_ = ~new_n503_ & new_n1443_;
  assign new_n1445_ = new_n472_ & ~new_n1444_;
  assign new_n1446_ = ~new_n472_ & new_n1444_;
  assign new_n1447_ = ~new_n1445_ & ~new_n1446_;
  assign new_n1448_ = ~new_n1442_ & new_n1447_;
  assign new_n1449_ = new_n1441_ & ~new_n1448_;
  assign new_n1450_ = ~new_n1441_ & new_n1448_;
  assign new_n1451_ = ~new_n1449_ & ~new_n1450_;
  assign new_n1452_ = ~new_n1438_ & ~new_n1451_;
  assign new_n1453_ = new_n1438_ & new_n1451_;
  assign new_n1454_ = ~new_n1452_ & ~new_n1453_;
  assign new_n1455_ = new_n442_ & ~new_n1454_;
  assign new_n1456_ = ~new_n474_ & ~new_n505_;
  assign new_n1457_ = ~new_n507_ & new_n1456_;
  assign new_n1458_ = new_n453_ & ~new_n1456_;
  assign new_n1459_ = ~new_n1457_ & ~new_n1458_;
  assign new_n1460_ = ~new_n473_ & new_n1325_;
  assign new_n1461_ = new_n448_ & ~new_n1460_;
  assign new_n1462_ = ~new_n448_ & new_n1460_;
  assign new_n1463_ = ~new_n1461_ & ~new_n1462_;
  assign new_n1464_ = new_n1459_ & new_n1463_;
  assign new_n1465_ = ~new_n1459_ & ~new_n1463_;
  assign new_n1466_ = ~new_n1464_ & ~new_n1465_;
  assign new_n1467_ = ~new_n466_ & ~new_n470_;
  assign new_n1468_ = ~new_n502_ & ~new_n1467_;
  assign new_n1469_ = new_n1441_ & new_n1468_;
  assign new_n1470_ = ~new_n1441_ & ~new_n1468_;
  assign new_n1471_ = ~new_n1469_ & ~new_n1470_;
  assign new_n1472_ = ~new_n1466_ & ~new_n1471_;
  assign new_n1473_ = new_n1466_ & new_n1471_;
  assign new_n1474_ = ~new_n1472_ & ~new_n1473_;
  assign new_n1475_ = ~new_n442_ & ~new_n1474_;
  assign new_n1476_ = ~new_n1455_ & ~new_n1475_;
  assign new_n1477_ = ~new_n491_ & ~new_n512_;
  assign new_n1478_ = ~new_n513_ & ~new_n1477_;
  assign new_n1479_ = new_n497_ & new_n1478_;
  assign new_n1480_ = ~new_n497_ & ~new_n1478_;
  assign new_n1481_ = ~new_n1479_ & ~new_n1480_;
  assign new_n1482_ = new_n481_ & ~new_n1481_;
  assign new_n1483_ = ~new_n481_ & new_n1481_;
  assign new_n1484_ = ~new_n1482_ & ~new_n1483_;
  assign new_n1485_ = new_n485_ & ~new_n1484_;
  assign new_n1486_ = ~new_n485_ & new_n1484_;
  assign new_n1487_ = ~new_n1485_ & ~new_n1486_;
  assign new_n1488_ = new_n1362_ & new_n1487_;
  assign new_n1489_ = ~new_n481_ & ~new_n484_;
  assign new_n1490_ = ~new_n511_ & ~new_n1489_;
  assign new_n1491_ = ~new_n487_ & new_n512_;
  assign new_n1492_ = ~new_n490_ & new_n1491_;
  assign new_n1493_ = ~new_n491_ & ~new_n1491_;
  assign new_n1494_ = ~new_n1492_ & ~new_n1493_;
  assign new_n1495_ = new_n497_ & ~new_n1494_;
  assign new_n1496_ = ~new_n497_ & new_n1494_;
  assign new_n1497_ = ~new_n1495_ & ~new_n1496_;
  assign new_n1498_ = new_n1490_ & ~new_n1497_;
  assign new_n1499_ = ~new_n1490_ & new_n1497_;
  assign new_n1500_ = ~new_n1498_ & ~new_n1499_;
  assign new_n1501_ = ~new_n1362_ & new_n1500_;
  assign new_n1502_ = ~new_n1488_ & ~new_n1501_;
  assign new_n1503_ = new_n492_ & ~new_n1502_;
  assign new_n1504_ = ~new_n492_ & new_n1502_;
  assign new_n1505_ = ~new_n1503_ & ~new_n1504_;
  assign new_n1506_ = new_n1476_ & new_n1505_;
  assign new_n1507_ = ~new_n1476_ & ~new_n1505_;
  assign po49 = new_n1506_ | new_n1507_;
  assign new_n1509_ = ~new_n524_ & ~new_n530_;
  assign new_n1510_ = ~new_n554_ & new_n1509_;
  assign new_n1511_ = ~new_n526_ & new_n1510_;
  assign new_n1512_ = new_n524_ & ~new_n1334_;
  assign new_n1513_ = ~new_n526_ & ~new_n1512_;
  assign new_n1514_ = ~new_n1510_ & ~new_n1513_;
  assign new_n1515_ = ~new_n1511_ & ~new_n1514_;
  assign new_n1516_ = new_n532_ & ~new_n545_;
  assign new_n1517_ = ~new_n532_ & new_n545_;
  assign new_n1518_ = ~new_n1516_ & ~new_n1517_;
  assign new_n1519_ = ~new_n521_ & ~new_n524_;
  assign new_n1520_ = ~new_n533_ & ~new_n1519_;
  assign new_n1521_ = new_n1336_ & ~new_n1520_;
  assign new_n1522_ = ~new_n1336_ & new_n1520_;
  assign new_n1523_ = ~new_n1521_ & ~new_n1522_;
  assign new_n1524_ = new_n540_ & ~new_n1523_;
  assign new_n1525_ = ~new_n540_ & new_n1523_;
  assign new_n1526_ = ~new_n1524_ & ~new_n1525_;
  assign new_n1527_ = ~new_n1518_ & new_n1526_;
  assign new_n1528_ = new_n1518_ & ~new_n1526_;
  assign new_n1529_ = ~new_n1527_ & ~new_n1528_;
  assign new_n1530_ = new_n1515_ & ~new_n1529_;
  assign new_n1531_ = ~new_n1515_ & new_n1529_;
  assign new_n1532_ = ~new_n1530_ & ~new_n1531_;
  assign new_n1533_ = new_n518_ & new_n1532_;
  assign new_n1534_ = ~new_n524_ & ~new_n549_;
  assign new_n1535_ = ~new_n550_ & ~new_n1534_;
  assign new_n1536_ = new_n532_ & new_n1535_;
  assign new_n1537_ = ~new_n532_ & ~new_n1535_;
  assign new_n1538_ = ~new_n1536_ & ~new_n1537_;
  assign new_n1539_ = ~new_n527_ & ~new_n533_;
  assign new_n1540_ = ~new_n550_ & new_n1539_;
  assign new_n1541_ = new_n540_ & ~new_n1540_;
  assign new_n1542_ = ~new_n540_ & new_n1540_;
  assign new_n1543_ = ~new_n1541_ & ~new_n1542_;
  assign new_n1544_ = ~new_n535_ & new_n1334_;
  assign new_n1545_ = ~new_n1336_ & new_n1544_;
  assign new_n1546_ = new_n544_ & ~new_n1544_;
  assign new_n1547_ = ~new_n1545_ & ~new_n1546_;
  assign new_n1548_ = new_n545_ & ~new_n1547_;
  assign new_n1549_ = ~new_n545_ & new_n1547_;
  assign new_n1550_ = ~new_n1548_ & ~new_n1549_;
  assign new_n1551_ = new_n1543_ & new_n1550_;
  assign new_n1552_ = ~new_n1543_ & ~new_n1550_;
  assign new_n1553_ = ~new_n1551_ & ~new_n1552_;
  assign new_n1554_ = ~new_n1538_ & ~new_n1553_;
  assign new_n1555_ = new_n1538_ & new_n1553_;
  assign new_n1556_ = ~new_n1554_ & ~new_n1555_;
  assign new_n1557_ = ~new_n518_ & new_n1556_;
  assign new_n1558_ = ~new_n1533_ & ~new_n1557_;
  assign new_n1559_ = ~new_n286_ & new_n1389_;
  assign new_n1560_ = ~new_n287_ & new_n567_;
  assign new_n1561_ = new_n561_ & new_n566_;
  assign new_n1562_ = ~new_n1560_ & ~new_n1561_;
  assign new_n1563_ = ~new_n1389_ & new_n1562_;
  assign new_n1564_ = ~new_n1559_ & ~new_n1563_;
  assign new_n1565_ = new_n1558_ & ~new_n1564_;
  assign new_n1566_ = ~new_n1558_ & new_n1564_;
  assign po50 = ~new_n1565_ & ~new_n1566_;
  assign new_n1568_ = new_n377_ & ~new_n392_;
  assign new_n1569_ = ~new_n377_ & new_n392_;
  assign new_n1570_ = ~new_n1568_ & ~new_n1569_;
  assign new_n1571_ = ~new_n368_ & ~new_n375_;
  assign new_n1572_ = ~new_n401_ & new_n1571_;
  assign new_n1573_ = ~new_n370_ & new_n1572_;
  assign new_n1574_ = new_n368_ & ~new_n1392_;
  assign new_n1575_ = ~new_n370_ & ~new_n1574_;
  assign new_n1576_ = ~new_n1572_ & ~new_n1575_;
  assign new_n1577_ = ~new_n1573_ & ~new_n1576_;
  assign new_n1578_ = ~new_n364_ & ~new_n368_;
  assign new_n1579_ = ~new_n378_ & ~new_n1578_;
  assign new_n1580_ = new_n1394_ & ~new_n1579_;
  assign new_n1581_ = ~new_n1394_ & new_n1579_;
  assign new_n1582_ = ~new_n1580_ & ~new_n1581_;
  assign new_n1583_ = new_n386_ & ~new_n1582_;
  assign new_n1584_ = ~new_n386_ & new_n1582_;
  assign new_n1585_ = ~new_n1583_ & ~new_n1584_;
  assign new_n1586_ = new_n1577_ & new_n1585_;
  assign new_n1587_ = ~new_n1577_ & ~new_n1585_;
  assign new_n1588_ = ~new_n1586_ & ~new_n1587_;
  assign new_n1589_ = ~new_n1570_ & new_n1588_;
  assign new_n1590_ = new_n1570_ & ~new_n1588_;
  assign new_n1591_ = ~new_n1589_ & ~new_n1590_;
  assign new_n1592_ = new_n360_ & ~new_n1591_;
  assign new_n1593_ = ~new_n380_ & new_n1392_;
  assign new_n1594_ = ~new_n1394_ & new_n1593_;
  assign new_n1595_ = new_n391_ & ~new_n1593_;
  assign new_n1596_ = ~new_n1594_ & ~new_n1595_;
  assign new_n1597_ = ~new_n371_ & ~new_n378_;
  assign new_n1598_ = ~new_n397_ & new_n1597_;
  assign new_n1599_ = new_n386_ & ~new_n1598_;
  assign new_n1600_ = ~new_n386_ & new_n1598_;
  assign new_n1601_ = ~new_n1599_ & ~new_n1600_;
  assign new_n1602_ = new_n1596_ & new_n1601_;
  assign new_n1603_ = ~new_n1596_ & ~new_n1601_;
  assign new_n1604_ = ~new_n1602_ & ~new_n1603_;
  assign new_n1605_ = ~new_n368_ & ~new_n396_;
  assign new_n1606_ = ~new_n397_ & ~new_n1605_;
  assign new_n1607_ = new_n1570_ & new_n1606_;
  assign new_n1608_ = ~new_n1570_ & ~new_n1606_;
  assign new_n1609_ = ~new_n1607_ & ~new_n1608_;
  assign new_n1610_ = new_n1604_ & new_n1609_;
  assign new_n1611_ = ~new_n1604_ & ~new_n1609_;
  assign new_n1612_ = ~new_n360_ & ~new_n1611_;
  assign new_n1613_ = ~new_n1610_ & new_n1612_;
  assign new_n1614_ = ~new_n1592_ & ~new_n1613_;
  assign new_n1615_ = ~new_n431_ & new_n437_;
  assign new_n1616_ = ~new_n438_ & ~new_n1615_;
  assign new_n1617_ = new_n426_ & ~new_n1616_;
  assign new_n1618_ = ~new_n426_ & new_n1616_;
  assign new_n1619_ = ~new_n1617_ & ~new_n1618_;
  assign new_n1620_ = ~new_n418_ & new_n1619_;
  assign new_n1621_ = new_n418_ & ~new_n1619_;
  assign new_n1622_ = ~new_n1620_ & ~new_n1621_;
  assign new_n1623_ = new_n413_ & new_n1622_;
  assign new_n1624_ = ~new_n413_ & ~new_n1622_;
  assign new_n1625_ = ~new_n1623_ & ~new_n1624_;
  assign new_n1626_ = new_n407_ & new_n1625_;
  assign new_n1627_ = ~new_n413_ & ~new_n417_;
  assign new_n1628_ = ~new_n436_ & ~new_n1627_;
  assign new_n1629_ = ~new_n420_ & new_n437_;
  assign new_n1630_ = ~new_n431_ & new_n1629_;
  assign new_n1631_ = ~new_n430_ & ~new_n1629_;
  assign new_n1632_ = ~new_n1630_ & ~new_n1631_;
  assign new_n1633_ = ~new_n426_ & ~new_n1632_;
  assign new_n1634_ = new_n426_ & new_n1632_;
  assign new_n1635_ = ~new_n1633_ & ~new_n1634_;
  assign new_n1636_ = new_n1628_ & new_n1635_;
  assign new_n1637_ = ~new_n1628_ & ~new_n1635_;
  assign new_n1638_ = ~new_n1636_ & ~new_n1637_;
  assign new_n1639_ = ~new_n407_ & new_n1638_;
  assign new_n1640_ = ~new_n1626_ & ~new_n1639_;
  assign new_n1641_ = new_n432_ & ~new_n1640_;
  assign new_n1642_ = ~new_n432_ & new_n1640_;
  assign new_n1643_ = ~new_n1641_ & ~new_n1642_;
  assign new_n1644_ = new_n1614_ & new_n1643_;
  assign new_n1645_ = ~new_n1614_ & ~new_n1643_;
  assign po51 = ~new_n1644_ & ~new_n1645_;
  assign new_n1647_ = new_n317_ & new_n319_;
  assign new_n1648_ = ~new_n296_ & new_n1647_;
  assign new_n1649_ = ~new_n314_ & ~new_n1648_;
  assign new_n1650_ = new_n914_ & ~new_n1649_;
  assign new_n1651_ = ~new_n914_ & new_n1649_;
  assign new_n1652_ = ~new_n1650_ & ~new_n1651_;
  assign new_n1653_ = ~new_n281_ & new_n1647_;
  assign new_n1654_ = ~new_n312_ & ~new_n1653_;
  assign new_n1655_ = new_n277_ & ~new_n281_;
  assign new_n1656_ = ~new_n1654_ & new_n1655_;
  assign new_n1657_ = new_n1654_ & ~new_n1655_;
  assign new_n1658_ = ~new_n1656_ & ~new_n1657_;
  assign new_n1659_ = new_n282_ & ~new_n306_;
  assign new_n1660_ = new_n925_ & ~new_n1659_;
  assign new_n1661_ = new_n307_ & ~new_n1660_;
  assign new_n1662_ = ~new_n307_ & new_n1660_;
  assign new_n1663_ = ~new_n1661_ & ~new_n1662_;
  assign new_n1664_ = new_n1658_ & ~new_n1663_;
  assign new_n1665_ = ~new_n1658_ & new_n1663_;
  assign new_n1666_ = ~new_n1664_ & ~new_n1665_;
  assign new_n1667_ = new_n1652_ & ~new_n1666_;
  assign new_n1668_ = ~new_n1652_ & new_n1666_;
  assign new_n1669_ = ~new_n1667_ & ~new_n1668_;
  assign new_n1670_ = pi203 & ~new_n1669_;
  assign new_n1671_ = new_n314_ & ~new_n914_;
  assign new_n1672_ = ~new_n314_ & new_n914_;
  assign new_n1673_ = ~new_n1671_ & ~new_n1672_;
  assign new_n1674_ = new_n277_ & ~new_n312_;
  assign new_n1675_ = ~new_n277_ & ~new_n301_;
  assign new_n1676_ = ~new_n310_ & new_n1675_;
  assign new_n1677_ = new_n282_ & ~new_n1676_;
  assign new_n1678_ = ~new_n282_ & new_n1676_;
  assign new_n1679_ = ~new_n1677_ & ~new_n1678_;
  assign new_n1680_ = ~new_n1674_ & new_n1679_;
  assign new_n1681_ = ~new_n277_ & ~new_n306_;
  assign new_n1682_ = ~new_n305_ & ~new_n1681_;
  assign new_n1683_ = new_n1680_ & ~new_n1682_;
  assign new_n1684_ = ~new_n1680_ & new_n1682_;
  assign new_n1685_ = ~new_n1683_ & ~new_n1684_;
  assign new_n1686_ = new_n1673_ & ~new_n1685_;
  assign new_n1687_ = ~new_n1673_ & new_n1685_;
  assign new_n1688_ = ~new_n1686_ & ~new_n1687_;
  assign new_n1689_ = ~pi203 & ~new_n1688_;
  assign new_n1690_ = ~new_n1670_ & ~new_n1689_;
  assign new_n1691_ = ~new_n319_ & ~new_n320_;
  assign new_n1692_ = ~new_n321_ & ~new_n1691_;
  assign new_n1693_ = new_n343_ & new_n355_;
  assign new_n1694_ = new_n342_ & ~new_n355_;
  assign new_n1695_ = ~new_n1693_ & ~new_n1694_;
  assign new_n1696_ = new_n350_ & ~new_n1695_;
  assign new_n1697_ = ~new_n350_ & new_n1695_;
  assign new_n1698_ = ~new_n1696_ & ~new_n1697_;
  assign new_n1699_ = ~new_n331_ & new_n336_;
  assign new_n1700_ = new_n331_ & ~new_n336_;
  assign new_n1701_ = ~new_n1699_ & ~new_n1700_;
  assign new_n1702_ = ~new_n1698_ & ~new_n1701_;
  assign new_n1703_ = new_n1698_ & new_n1701_;
  assign new_n1704_ = ~new_n1702_ & ~new_n1703_;
  assign new_n1705_ = new_n325_ & ~new_n1704_;
  assign new_n1706_ = ~new_n331_ & ~new_n335_;
  assign new_n1707_ = ~new_n354_ & ~new_n1706_;
  assign new_n1708_ = ~new_n344_ & ~new_n350_;
  assign new_n1709_ = ~new_n351_ & ~new_n1708_;
  assign new_n1710_ = new_n1707_ & ~new_n1709_;
  assign new_n1711_ = ~new_n1707_ & new_n1709_;
  assign new_n1712_ = ~new_n1710_ & ~new_n1711_;
  assign new_n1713_ = ~new_n329_ & ~new_n1700_;
  assign new_n1714_ = ~new_n342_ & new_n1713_;
  assign new_n1715_ = ~new_n343_ & ~new_n1713_;
  assign new_n1716_ = ~new_n1714_ & ~new_n1715_;
  assign new_n1717_ = ~new_n1712_ & ~new_n1716_;
  assign new_n1718_ = new_n1712_ & new_n1716_;
  assign new_n1719_ = ~new_n1717_ & ~new_n1718_;
  assign new_n1720_ = ~new_n325_ & new_n1719_;
  assign new_n1721_ = ~new_n1705_ & ~new_n1720_;
  assign new_n1722_ = new_n1692_ & ~new_n1721_;
  assign new_n1723_ = ~new_n1692_ & new_n1721_;
  assign new_n1724_ = ~new_n1722_ & ~new_n1723_;
  assign new_n1725_ = new_n1690_ & new_n1724_;
  assign new_n1726_ = ~new_n1690_ & ~new_n1724_;
  assign po52 = ~new_n1725_ & ~new_n1726_;
endmodule


