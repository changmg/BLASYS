// Benchmark "c5315" written by ABC on Sat Jul 16 14:36:05 2022

module c5315 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71,
    po72, po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83,
    po84, po85, po86, po87, po88, po89, po90  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70,
    po71, po72, po73, po74, po75, po76, po77, po78, po79, po80, po81, po82,
    po83, po84, po85, po86, po87, po88, po89, po90;
  wire new_n276_, new_n277_, new_n278_, new_n280_, new_n281_, new_n282_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1064_,
    new_n1065_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1170_, new_n1171_,
    new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1223_, new_n1224_, new_n1225_,
    new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_;
  assign po00 = pi150 & pi153;
  assign po01 = pi065 & pi066;
  assign po02 = pi000 & pi133;
  assign po03 = pi062 & ~pi162;
  assign po04 = ~pi010 | pi161;
  assign po05 = ~pi135 | ~pi151;
  assign po07 = ~pi010 | ~pi011;
  assign po06 = ~pi064 | po07;
  assign new_n276_ = ~pi033 & pi160;
  assign new_n277_ = ~pi032 & ~pi160;
  assign new_n278_ = ~po07 & ~new_n277_;
  assign po08 = new_n276_ | ~new_n278_;
  assign new_n280_ = ~pi012 & pi160;
  assign new_n281_ = ~pi034 & ~pi160;
  assign new_n282_ = ~po07 & ~new_n281_;
  assign po09 = new_n280_ | ~new_n282_;
  assign po10 = ~pi031 | po07;
  assign new_n285_ = pi008 & pi160;
  assign new_n286_ = pi007 & ~pi160;
  assign new_n287_ = ~po07 & ~new_n286_;
  assign new_n288_ = ~new_n285_ & new_n287_;
  assign po11 = pi065 & ~new_n288_;
  assign new_n290_ = pi029 & pi160;
  assign new_n291_ = pi009 & ~pi160;
  assign new_n292_ = ~po07 & ~new_n291_;
  assign new_n293_ = ~new_n290_ & new_n292_;
  assign po12 = pi065 & ~new_n293_;
  assign new_n295_ = pi006 & pi160;
  assign new_n296_ = pi027 & ~pi160;
  assign new_n297_ = ~po07 & ~new_n296_;
  assign new_n298_ = ~new_n295_ & new_n297_;
  assign po13 = pi065 & ~new_n298_;
  assign new_n300_ = pi028 & pi160;
  assign new_n301_ = pi030 & ~pi160;
  assign new_n302_ = ~po07 & ~new_n301_;
  assign new_n303_ = ~new_n300_ & new_n302_;
  assign po14 = pi065 & ~new_n303_;
  assign new_n305_ = pi099 & pi118;
  assign new_n306_ = pi100 & ~pi118;
  assign new_n307_ = pi145 & ~new_n306_;
  assign new_n308_ = ~new_n305_ & new_n307_;
  assign new_n309_ = ~pi097 & pi118;
  assign new_n310_ = ~pi101 & ~pi118;
  assign new_n311_ = ~pi145 & ~new_n310_;
  assign new_n312_ = ~new_n309_ & new_n311_;
  assign new_n313_ = ~new_n308_ & ~new_n312_;
  assign new_n314_ = pi099 & pi116;
  assign new_n315_ = pi100 & ~pi116;
  assign new_n316_ = pi144 & ~new_n315_;
  assign new_n317_ = ~new_n314_ & new_n316_;
  assign new_n318_ = ~pi097 & pi116;
  assign new_n319_ = ~pi101 & ~pi116;
  assign new_n320_ = ~pi144 & ~new_n319_;
  assign new_n321_ = ~new_n318_ & new_n320_;
  assign new_n322_ = ~new_n317_ & ~new_n321_;
  assign new_n323_ = new_n313_ & new_n322_;
  assign new_n324_ = pi120 & ~pi166;
  assign new_n325_ = ~pi120 & ~pi165;
  assign new_n326_ = pi146 & ~new_n325_;
  assign new_n327_ = ~new_n324_ & new_n326_;
  assign new_n328_ = pi120 & pi163;
  assign new_n329_ = ~pi120 & pi164;
  assign new_n330_ = ~pi146 & ~new_n329_;
  assign new_n331_ = ~new_n328_ & new_n330_;
  assign new_n332_ = ~new_n327_ & ~new_n331_;
  assign new_n333_ = ~pi100 & ~pi114;
  assign new_n334_ = ~pi099 & pi114;
  assign new_n335_ = ~new_n333_ & ~new_n334_;
  assign new_n336_ = ~pi101 & ~pi112;
  assign new_n337_ = ~pi097 & pi112;
  assign new_n338_ = ~new_n336_ & ~new_n337_;
  assign new_n339_ = new_n335_ & ~new_n338_;
  assign new_n340_ = ~pi100 & ~pi129;
  assign new_n341_ = ~pi099 & pi129;
  assign new_n342_ = ~new_n340_ & ~new_n341_;
  assign new_n343_ = ~pi147 & ~pi163;
  assign new_n344_ = pi147 & pi166;
  assign new_n345_ = ~new_n343_ & ~new_n344_;
  assign new_n346_ = new_n342_ & new_n345_;
  assign new_n347_ = new_n339_ & new_n346_;
  assign new_n348_ = new_n332_ & new_n347_;
  assign new_n349_ = pi127 & ~pi166;
  assign new_n350_ = ~pi127 & ~pi165;
  assign new_n351_ = pi149 & ~new_n350_;
  assign new_n352_ = ~new_n349_ & new_n351_;
  assign new_n353_ = pi127 & pi163;
  assign new_n354_ = ~pi127 & pi164;
  assign new_n355_ = ~pi149 & ~new_n354_;
  assign new_n356_ = ~new_n353_ & new_n355_;
  assign new_n357_ = ~new_n352_ & ~new_n356_;
  assign new_n358_ = pi125 & ~pi166;
  assign new_n359_ = ~pi125 & ~pi165;
  assign new_n360_ = pi148 & ~new_n359_;
  assign new_n361_ = ~new_n358_ & new_n360_;
  assign new_n362_ = pi125 & pi163;
  assign new_n363_ = ~pi125 & pi164;
  assign new_n364_ = ~pi148 & ~new_n363_;
  assign new_n365_ = ~new_n362_ & new_n364_;
  assign new_n366_ = ~new_n361_ & ~new_n365_;
  assign new_n367_ = new_n357_ & new_n366_;
  assign new_n368_ = new_n348_ & new_n367_;
  assign po15 = new_n323_ & new_n368_;
  assign new_n370_ = pi091 & ~pi163;
  assign new_n371_ = ~pi091 & ~pi164;
  assign new_n372_ = ~pi143 & ~new_n371_;
  assign new_n373_ = ~new_n370_ & new_n372_;
  assign new_n374_ = pi091 & pi143;
  assign new_n375_ = ~pi166 & new_n374_;
  assign new_n376_ = ~pi091 & pi143;
  assign new_n377_ = ~pi165 & new_n376_;
  assign new_n378_ = ~new_n375_ & ~new_n377_;
  assign new_n379_ = ~new_n373_ & new_n378_;
  assign new_n380_ = pi089 & ~pi163;
  assign new_n381_ = ~pi089 & ~pi164;
  assign new_n382_ = ~pi142 & ~new_n381_;
  assign new_n383_ = ~new_n380_ & new_n382_;
  assign new_n384_ = pi089 & pi142;
  assign new_n385_ = ~pi166 & new_n384_;
  assign new_n386_ = ~pi089 & pi142;
  assign new_n387_ = ~pi165 & new_n386_;
  assign new_n388_ = ~new_n385_ & ~new_n387_;
  assign new_n389_ = ~new_n383_ & new_n388_;
  assign new_n390_ = pi106 & ~pi166;
  assign new_n391_ = ~pi106 & ~pi165;
  assign new_n392_ = pi138 & ~new_n391_;
  assign new_n393_ = ~new_n390_ & new_n392_;
  assign new_n394_ = pi106 & pi163;
  assign new_n395_ = ~pi106 & pi164;
  assign new_n396_ = ~pi138 & ~new_n395_;
  assign new_n397_ = ~new_n394_ & new_n396_;
  assign new_n398_ = ~new_n393_ & ~new_n397_;
  assign new_n399_ = ~new_n389_ & new_n398_;
  assign new_n400_ = ~new_n379_ & new_n399_;
  assign new_n401_ = pi102 & ~pi166;
  assign new_n402_ = ~pi102 & ~pi165;
  assign new_n403_ = pi136 & ~new_n402_;
  assign new_n404_ = ~new_n401_ & new_n403_;
  assign new_n405_ = pi102 & pi163;
  assign new_n406_ = ~pi102 & pi164;
  assign new_n407_ = ~pi136 & ~new_n406_;
  assign new_n408_ = ~new_n405_ & new_n407_;
  assign new_n409_ = ~new_n404_ & ~new_n408_;
  assign new_n410_ = pi095 & ~pi163;
  assign new_n411_ = ~pi095 & ~pi164;
  assign new_n412_ = ~pi140 & ~new_n411_;
  assign new_n413_ = ~new_n410_ & new_n412_;
  assign new_n414_ = pi095 & pi140;
  assign new_n415_ = ~pi166 & new_n414_;
  assign new_n416_ = ~pi095 & pi140;
  assign new_n417_ = ~pi165 & new_n416_;
  assign new_n418_ = ~new_n415_ & ~new_n417_;
  assign new_n419_ = ~new_n413_ & new_n418_;
  assign new_n420_ = new_n409_ & ~new_n419_;
  assign new_n421_ = pi087 & pi099;
  assign new_n422_ = ~pi087 & pi100;
  assign new_n423_ = pi141 & ~new_n422_;
  assign new_n424_ = ~new_n421_ & new_n423_;
  assign new_n425_ = pi087 & ~pi097;
  assign new_n426_ = ~pi087 & ~pi101;
  assign new_n427_ = ~pi141 & ~new_n426_;
  assign new_n428_ = ~new_n425_ & new_n427_;
  assign new_n429_ = ~new_n424_ & ~new_n428_;
  assign new_n430_ = pi093 & ~pi163;
  assign new_n431_ = ~pi093 & ~pi164;
  assign new_n432_ = ~pi139 & ~new_n431_;
  assign new_n433_ = ~new_n430_ & new_n432_;
  assign new_n434_ = pi093 & pi139;
  assign new_n435_ = ~pi166 & new_n434_;
  assign new_n436_ = ~pi093 & pi139;
  assign new_n437_ = ~pi165 & new_n436_;
  assign new_n438_ = ~new_n435_ & ~new_n437_;
  assign new_n439_ = ~new_n433_ & new_n438_;
  assign new_n440_ = new_n429_ & ~new_n439_;
  assign new_n441_ = pi108 & ~pi166;
  assign new_n442_ = ~pi108 & ~pi165;
  assign new_n443_ = pi134 & ~new_n442_;
  assign new_n444_ = ~new_n441_ & new_n443_;
  assign new_n445_ = pi108 & pi163;
  assign new_n446_ = ~pi108 & pi164;
  assign new_n447_ = ~pi134 & ~new_n446_;
  assign new_n448_ = ~new_n445_ & new_n447_;
  assign new_n449_ = ~new_n444_ & ~new_n448_;
  assign new_n450_ = pi104 & ~pi166;
  assign new_n451_ = ~pi104 & ~pi165;
  assign new_n452_ = pi137 & ~new_n451_;
  assign new_n453_ = ~new_n450_ & new_n452_;
  assign new_n454_ = pi104 & pi163;
  assign new_n455_ = ~pi104 & pi164;
  assign new_n456_ = ~pi137 & ~new_n455_;
  assign new_n457_ = ~new_n454_ & new_n456_;
  assign new_n458_ = ~new_n453_ & ~new_n457_;
  assign new_n459_ = new_n449_ & new_n458_;
  assign new_n460_ = new_n440_ & new_n459_;
  assign new_n461_ = new_n420_ & new_n460_;
  assign po16 = new_n400_ & new_n461_;
  assign new_n463_ = ~pi090 & pi123;
  assign new_n464_ = ~pi089 & ~pi123;
  assign new_n465_ = ~new_n463_ & ~new_n464_;
  assign new_n466_ = pi142 & new_n465_;
  assign new_n467_ = ~pi142 & ~new_n465_;
  assign new_n468_ = ~new_n466_ & ~new_n467_;
  assign new_n469_ = ~pi094 & pi123;
  assign new_n470_ = ~pi093 & ~pi123;
  assign new_n471_ = ~new_n469_ & ~new_n470_;
  assign new_n472_ = pi139 & new_n471_;
  assign new_n473_ = ~pi139 & ~new_n471_;
  assign new_n474_ = ~new_n472_ & ~new_n473_;
  assign new_n475_ = ~pi092 & pi123;
  assign new_n476_ = ~pi091 & ~pi123;
  assign new_n477_ = ~new_n475_ & ~new_n476_;
  assign new_n478_ = pi143 & new_n477_;
  assign new_n479_ = ~pi143 & ~new_n477_;
  assign new_n480_ = ~new_n478_ & ~new_n479_;
  assign new_n481_ = new_n474_ & new_n480_;
  assign new_n482_ = new_n468_ & new_n481_;
  assign new_n483_ = ~pi088 & pi123;
  assign new_n484_ = ~pi087 & ~pi123;
  assign new_n485_ = ~new_n483_ & ~new_n484_;
  assign new_n486_ = pi141 & new_n485_;
  assign new_n487_ = ~pi141 & ~new_n485_;
  assign new_n488_ = ~new_n486_ & ~new_n487_;
  assign new_n489_ = new_n482_ & new_n488_;
  assign new_n490_ = ~pi096 & pi123;
  assign new_n491_ = ~pi095 & ~pi123;
  assign new_n492_ = ~new_n490_ & ~new_n491_;
  assign new_n493_ = pi140 & new_n492_;
  assign new_n494_ = ~pi140 & ~new_n492_;
  assign new_n495_ = ~new_n493_ & ~new_n494_;
  assign new_n496_ = ~pi109 & pi123;
  assign new_n497_ = ~pi108 & ~pi123;
  assign new_n498_ = ~new_n496_ & ~new_n497_;
  assign new_n499_ = pi134 & new_n498_;
  assign new_n500_ = ~pi134 & ~new_n498_;
  assign new_n501_ = ~new_n499_ & ~new_n500_;
  assign new_n502_ = ~pi107 & pi123;
  assign new_n503_ = ~pi106 & ~pi123;
  assign new_n504_ = ~new_n502_ & ~new_n503_;
  assign new_n505_ = pi138 & new_n504_;
  assign new_n506_ = ~pi138 & ~new_n504_;
  assign new_n507_ = ~new_n505_ & ~new_n506_;
  assign new_n508_ = new_n501_ & new_n507_;
  assign new_n509_ = ~pi103 & pi123;
  assign new_n510_ = ~pi102 & ~pi123;
  assign new_n511_ = ~new_n509_ & ~new_n510_;
  assign new_n512_ = pi136 & new_n511_;
  assign new_n513_ = ~pi136 & ~new_n511_;
  assign new_n514_ = ~new_n512_ & ~new_n513_;
  assign new_n515_ = ~pi105 & pi123;
  assign new_n516_ = ~pi104 & ~pi123;
  assign new_n517_ = ~new_n515_ & ~new_n516_;
  assign new_n518_ = pi137 & new_n517_;
  assign new_n519_ = ~pi137 & ~new_n517_;
  assign new_n520_ = ~new_n518_ & ~new_n519_;
  assign new_n521_ = new_n514_ & new_n520_;
  assign new_n522_ = new_n508_ & new_n521_;
  assign new_n523_ = new_n495_ & new_n522_;
  assign po17 = new_n489_ & new_n523_;
  assign new_n525_ = ~pi121 & pi122;
  assign new_n526_ = ~pi120 & ~pi122;
  assign new_n527_ = ~new_n525_ & ~new_n526_;
  assign new_n528_ = pi146 & new_n527_;
  assign new_n529_ = ~pi146 & ~new_n527_;
  assign new_n530_ = ~new_n528_ & ~new_n529_;
  assign new_n531_ = pi122 & ~pi128;
  assign new_n532_ = ~pi122 & ~pi127;
  assign new_n533_ = ~new_n531_ & ~new_n532_;
  assign new_n534_ = pi149 & new_n533_;
  assign new_n535_ = ~pi149 & ~new_n533_;
  assign new_n536_ = ~new_n534_ & ~new_n535_;
  assign new_n537_ = pi122 & ~pi130;
  assign new_n538_ = ~pi122 & ~pi129;
  assign new_n539_ = ~new_n537_ & ~new_n538_;
  assign new_n540_ = new_n536_ & ~new_n539_;
  assign new_n541_ = pi122 & ~pi124;
  assign new_n542_ = pi147 & ~new_n541_;
  assign new_n543_ = ~pi147 & new_n541_;
  assign new_n544_ = ~new_n542_ & ~new_n543_;
  assign new_n545_ = pi122 & ~pi126;
  assign new_n546_ = ~pi122 & ~pi125;
  assign new_n547_ = ~new_n545_ & ~new_n546_;
  assign new_n548_ = pi148 & new_n547_;
  assign new_n549_ = ~pi148 & ~new_n547_;
  assign new_n550_ = ~new_n548_ & ~new_n549_;
  assign new_n551_ = new_n544_ & new_n550_;
  assign new_n552_ = new_n540_ & new_n551_;
  assign new_n553_ = new_n530_ & new_n552_;
  assign new_n554_ = ~pi113 & pi122;
  assign new_n555_ = ~pi112 & ~pi122;
  assign new_n556_ = ~new_n554_ & ~new_n555_;
  assign new_n557_ = ~pi115 & pi122;
  assign new_n558_ = ~pi114 & ~pi122;
  assign new_n559_ = ~new_n557_ & ~new_n558_;
  assign new_n560_ = ~new_n556_ & ~new_n559_;
  assign new_n561_ = ~pi117 & pi122;
  assign new_n562_ = ~pi116 & ~pi122;
  assign new_n563_ = ~new_n561_ & ~new_n562_;
  assign new_n564_ = pi144 & new_n563_;
  assign new_n565_ = ~pi144 & ~new_n563_;
  assign new_n566_ = ~new_n564_ & ~new_n565_;
  assign new_n567_ = ~pi119 & pi122;
  assign new_n568_ = ~pi118 & ~pi122;
  assign new_n569_ = ~new_n567_ & ~new_n568_;
  assign new_n570_ = pi145 & new_n569_;
  assign new_n571_ = ~pi145 & ~new_n569_;
  assign new_n572_ = ~new_n570_ & ~new_n571_;
  assign new_n573_ = new_n566_ & new_n572_;
  assign new_n574_ = new_n560_ & new_n573_;
  assign po18 = new_n553_ & new_n574_;
  assign new_n576_ = ~pi116 & ~pi118;
  assign new_n577_ = pi116 & pi118;
  assign new_n578_ = ~new_n576_ & ~new_n577_;
  assign new_n579_ = ~pi129 & ~pi131;
  assign new_n580_ = pi129 & pi131;
  assign new_n581_ = ~new_n579_ & ~new_n580_;
  assign new_n582_ = new_n578_ & ~new_n581_;
  assign new_n583_ = ~new_n578_ & new_n581_;
  assign new_n584_ = ~new_n582_ & ~new_n583_;
  assign new_n585_ = ~pi125 & ~pi127;
  assign new_n586_ = pi125 & pi127;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign new_n588_ = pi120 & new_n587_;
  assign new_n589_ = ~pi120 & ~new_n587_;
  assign new_n590_ = ~new_n588_ & ~new_n589_;
  assign new_n591_ = pi112 & ~pi114;
  assign new_n592_ = ~pi112 & pi114;
  assign new_n593_ = ~new_n591_ & ~new_n592_;
  assign new_n594_ = new_n590_ & ~new_n593_;
  assign new_n595_ = ~new_n590_ & new_n593_;
  assign new_n596_ = ~new_n594_ & ~new_n595_;
  assign new_n597_ = new_n584_ & new_n596_;
  assign new_n598_ = ~new_n584_ & ~new_n596_;
  assign po19 = ~new_n597_ & ~new_n598_;
  assign new_n600_ = ~pi091 & ~pi093;
  assign new_n601_ = pi091 & pi093;
  assign new_n602_ = ~new_n600_ & ~new_n601_;
  assign new_n603_ = ~pi095 & ~pi102;
  assign new_n604_ = pi095 & pi102;
  assign new_n605_ = ~new_n603_ & ~new_n604_;
  assign new_n606_ = pi108 & new_n605_;
  assign new_n607_ = ~pi108 & ~new_n605_;
  assign new_n608_ = ~new_n606_ & ~new_n607_;
  assign new_n609_ = new_n602_ & ~new_n608_;
  assign new_n610_ = ~new_n602_ & new_n608_;
  assign new_n611_ = ~new_n609_ & ~new_n610_;
  assign new_n612_ = ~pi104 & ~pi106;
  assign new_n613_ = pi104 & pi106;
  assign new_n614_ = ~new_n612_ & ~new_n613_;
  assign new_n615_ = pi110 & new_n614_;
  assign new_n616_ = ~pi110 & ~new_n614_;
  assign new_n617_ = ~new_n615_ & ~new_n616_;
  assign new_n618_ = pi087 & ~pi089;
  assign new_n619_ = ~pi087 & pi089;
  assign new_n620_ = ~new_n618_ & ~new_n619_;
  assign new_n621_ = new_n617_ & ~new_n620_;
  assign new_n622_ = ~new_n617_ & new_n620_;
  assign new_n623_ = ~new_n621_ & ~new_n622_;
  assign new_n624_ = new_n611_ & new_n623_;
  assign new_n625_ = ~new_n611_ & ~new_n623_;
  assign po20 = new_n624_ | new_n625_;
  assign new_n627_ = new_n499_ & new_n507_;
  assign new_n628_ = ~new_n505_ & ~new_n518_;
  assign new_n629_ = ~new_n627_ & new_n628_;
  assign new_n630_ = ~new_n519_ & ~new_n629_;
  assign new_n631_ = ~new_n512_ & ~new_n630_;
  assign new_n632_ = ~new_n513_ & ~new_n631_;
  assign new_n633_ = ~new_n493_ & ~new_n632_;
  assign new_n634_ = ~new_n494_ & ~new_n633_;
  assign new_n635_ = new_n489_ & new_n634_;
  assign new_n636_ = new_n472_ & new_n480_;
  assign new_n637_ = ~new_n478_ & ~new_n636_;
  assign new_n638_ = ~new_n466_ & new_n637_;
  assign new_n639_ = ~new_n467_ & ~new_n638_;
  assign new_n640_ = ~new_n487_ & new_n639_;
  assign new_n641_ = ~new_n486_ & ~new_n640_;
  assign po21 = new_n635_ | ~new_n641_;
  assign new_n643_ = ~new_n534_ & ~new_n539_;
  assign new_n644_ = ~new_n535_ & ~new_n549_;
  assign new_n645_ = ~new_n643_ & new_n644_;
  assign new_n646_ = ~new_n548_ & ~new_n645_;
  assign new_n647_ = ~new_n543_ & ~new_n646_;
  assign new_n648_ = ~new_n542_ & ~new_n647_;
  assign new_n649_ = new_n530_ & ~new_n648_;
  assign new_n650_ = ~new_n528_ & ~new_n649_;
  assign new_n651_ = new_n573_ & ~new_n650_;
  assign new_n652_ = ~new_n564_ & ~new_n570_;
  assign new_n653_ = ~new_n565_ & ~new_n652_;
  assign new_n654_ = new_n560_ & ~new_n653_;
  assign po22 = new_n651_ | ~new_n654_;
  assign new_n656_ = ~pi020 & ~new_n539_;
  assign new_n657_ = pi020 & new_n539_;
  assign new_n658_ = ~new_n656_ & ~new_n657_;
  assign new_n659_ = pi173 & ~pi174;
  assign new_n660_ = ~new_n658_ & new_n659_;
  assign new_n661_ = ~pi173 & ~pi174;
  assign new_n662_ = ~new_n342_ & new_n661_;
  assign new_n663_ = ~pi173 & pi174;
  assign new_n664_ = pi059 & new_n663_;
  assign new_n665_ = ~new_n662_ & ~new_n664_;
  assign po23 = ~new_n660_ & new_n665_;
  assign new_n667_ = ~new_n536_ & new_n656_;
  assign new_n668_ = new_n536_ & ~new_n656_;
  assign new_n669_ = new_n659_ & ~new_n668_;
  assign new_n670_ = ~new_n667_ & new_n669_;
  assign new_n671_ = ~new_n357_ & new_n661_;
  assign new_n672_ = pi057 & new_n663_;
  assign new_n673_ = ~new_n671_ & ~new_n672_;
  assign po24 = ~new_n670_ & new_n673_;
  assign new_n675_ = pi001 & new_n501_;
  assign new_n676_ = ~pi001 & ~new_n501_;
  assign new_n677_ = ~new_n675_ & ~new_n676_;
  assign new_n678_ = new_n659_ & new_n677_;
  assign new_n679_ = ~new_n449_ & new_n661_;
  assign new_n680_ = pi047 & new_n663_;
  assign new_n681_ = ~new_n679_ & ~new_n680_;
  assign po25 = ~new_n678_ & new_n681_;
  assign new_n683_ = pi020 & new_n553_;
  assign new_n684_ = new_n650_ & ~new_n683_;
  assign new_n685_ = new_n573_ & ~new_n684_;
  assign new_n686_ = ~new_n653_ & ~new_n685_;
  assign new_n687_ = ~new_n556_ & ~new_n686_;
  assign new_n688_ = new_n556_ & new_n559_;
  assign new_n689_ = ~new_n560_ & ~new_n688_;
  assign new_n690_ = new_n686_ & new_n689_;
  assign po26 = new_n687_ | new_n690_;
  assign new_n692_ = ~pi169 & pi170;
  assign new_n693_ = ~po25 & new_n692_;
  assign new_n694_ = ~pi169 & ~pi170;
  assign new_n695_ = ~po23 & new_n694_;
  assign new_n696_ = ~pi021 & pi170;
  assign new_n697_ = ~pi002 & ~pi170;
  assign new_n698_ = pi169 & ~new_n697_;
  assign new_n699_ = ~new_n696_ & new_n698_;
  assign new_n700_ = ~new_n695_ & ~new_n699_;
  assign po27 = new_n693_ | ~new_n700_;
  assign new_n702_ = ~new_n552_ & new_n648_;
  assign new_n703_ = ~pi020 & new_n648_;
  assign new_n704_ = ~new_n702_ & ~new_n703_;
  assign new_n705_ = new_n530_ & ~new_n704_;
  assign new_n706_ = ~new_n530_ & new_n704_;
  assign new_n707_ = ~new_n705_ & ~new_n706_;
  assign new_n708_ = new_n659_ & ~new_n707_;
  assign new_n709_ = ~new_n332_ & new_n661_;
  assign new_n710_ = pi018 & new_n663_;
  assign new_n711_ = ~new_n709_ & ~new_n710_;
  assign po28 = ~new_n708_ & new_n711_;
  assign new_n713_ = ~pi020 & new_n646_;
  assign new_n714_ = new_n540_ & ~new_n549_;
  assign new_n715_ = new_n646_ & ~new_n714_;
  assign new_n716_ = ~new_n713_ & ~new_n715_;
  assign new_n717_ = new_n544_ & ~new_n716_;
  assign new_n718_ = ~new_n544_ & new_n716_;
  assign new_n719_ = ~new_n717_ & ~new_n718_;
  assign new_n720_ = new_n659_ & ~new_n719_;
  assign new_n721_ = ~new_n345_ & new_n661_;
  assign new_n722_ = pi058 & new_n663_;
  assign new_n723_ = ~new_n721_ & ~new_n722_;
  assign po29 = ~new_n720_ & new_n723_;
  assign new_n725_ = ~new_n534_ & new_n656_;
  assign new_n726_ = ~new_n535_ & ~new_n725_;
  assign new_n727_ = new_n550_ & ~new_n726_;
  assign new_n728_ = ~new_n550_ & new_n726_;
  assign new_n729_ = ~new_n727_ & ~new_n728_;
  assign new_n730_ = new_n659_ & ~new_n729_;
  assign new_n731_ = ~new_n366_ & new_n661_;
  assign new_n732_ = pi049 & new_n663_;
  assign new_n733_ = ~new_n731_ & ~new_n732_;
  assign po30 = ~new_n730_ & new_n733_;
  assign new_n735_ = pi171 & ~pi172;
  assign new_n736_ = ~po25 & new_n735_;
  assign new_n737_ = ~pi171 & ~pi172;
  assign new_n738_ = ~po23 & new_n737_;
  assign new_n739_ = ~pi021 & pi171;
  assign new_n740_ = ~pi002 & ~pi171;
  assign new_n741_ = pi172 & ~new_n740_;
  assign new_n742_ = ~new_n739_ & new_n741_;
  assign new_n743_ = ~new_n738_ & ~new_n742_;
  assign po31 = new_n736_ | ~new_n743_;
  assign new_n745_ = new_n508_ & new_n520_;
  assign new_n746_ = ~new_n630_ & ~new_n745_;
  assign new_n747_ = ~pi001 & ~new_n630_;
  assign new_n748_ = ~new_n746_ & ~new_n747_;
  assign new_n749_ = ~new_n512_ & ~new_n748_;
  assign new_n750_ = ~new_n513_ & ~new_n749_;
  assign new_n751_ = new_n495_ & ~new_n750_;
  assign new_n752_ = ~new_n495_ & new_n750_;
  assign new_n753_ = ~new_n751_ & ~new_n752_;
  assign new_n754_ = new_n659_ & ~new_n753_;
  assign new_n755_ = new_n419_ & new_n661_;
  assign new_n756_ = pi052 & new_n663_;
  assign new_n757_ = ~new_n755_ & ~new_n756_;
  assign po32 = ~new_n754_ & new_n757_;
  assign new_n759_ = ~new_n514_ & new_n748_;
  assign new_n760_ = new_n514_ & ~new_n748_;
  assign new_n761_ = ~new_n759_ & ~new_n760_;
  assign new_n762_ = new_n659_ & ~new_n761_;
  assign new_n763_ = ~new_n409_ & new_n661_;
  assign new_n764_ = pi056 & new_n663_;
  assign new_n765_ = ~new_n763_ & ~new_n764_;
  assign po33 = ~new_n762_ & new_n765_;
  assign new_n767_ = ~new_n499_ & ~new_n675_;
  assign new_n768_ = new_n507_ & ~new_n767_;
  assign new_n769_ = ~new_n505_ & ~new_n768_;
  assign new_n770_ = new_n520_ & ~new_n769_;
  assign new_n771_ = ~new_n520_ & new_n769_;
  assign new_n772_ = ~new_n770_ & ~new_n771_;
  assign new_n773_ = new_n659_ & new_n772_;
  assign new_n774_ = ~new_n458_ & new_n661_;
  assign new_n775_ = pi055 & new_n663_;
  assign new_n776_ = ~new_n774_ & ~new_n775_;
  assign po34 = ~new_n773_ & new_n776_;
  assign new_n778_ = ~new_n499_ & ~new_n507_;
  assign new_n779_ = ~new_n675_ & new_n778_;
  assign new_n780_ = ~new_n768_ & ~new_n779_;
  assign new_n781_ = new_n659_ & new_n780_;
  assign new_n782_ = ~new_n398_ & new_n661_;
  assign new_n783_ = pi054 & new_n663_;
  assign new_n784_ = ~new_n782_ & ~new_n783_;
  assign po35 = ~new_n781_ & new_n784_;
  assign new_n786_ = new_n563_ & ~new_n569_;
  assign new_n787_ = ~new_n563_ & new_n569_;
  assign new_n788_ = ~new_n786_ & ~new_n787_;
  assign new_n789_ = new_n689_ & ~new_n788_;
  assign new_n790_ = ~new_n689_ & new_n788_;
  assign new_n791_ = ~new_n789_ & ~new_n790_;
  assign new_n792_ = pi122 & ~pi132;
  assign new_n793_ = ~pi122 & ~pi131;
  assign new_n794_ = ~new_n792_ & ~new_n793_;
  assign new_n795_ = new_n539_ & ~new_n794_;
  assign new_n796_ = ~new_n539_ & new_n794_;
  assign new_n797_ = ~new_n795_ & ~new_n796_;
  assign new_n798_ = new_n533_ & ~new_n797_;
  assign new_n799_ = ~new_n533_ & new_n797_;
  assign new_n800_ = ~new_n798_ & ~new_n799_;
  assign new_n801_ = new_n547_ & new_n800_;
  assign new_n802_ = ~new_n547_ & ~new_n800_;
  assign new_n803_ = ~new_n801_ & ~new_n802_;
  assign new_n804_ = new_n527_ & ~new_n541_;
  assign new_n805_ = ~pi121 & new_n541_;
  assign new_n806_ = ~new_n804_ & ~new_n805_;
  assign new_n807_ = new_n803_ & ~new_n806_;
  assign new_n808_ = ~new_n803_ & new_n806_;
  assign new_n809_ = ~new_n807_ & ~new_n808_;
  assign new_n810_ = new_n791_ & new_n809_;
  assign new_n811_ = ~new_n791_ & ~new_n809_;
  assign po36 = new_n810_ | new_n811_;
  assign new_n813_ = ~new_n498_ & new_n511_;
  assign new_n814_ = new_n498_ & ~new_n511_;
  assign new_n815_ = ~new_n813_ & ~new_n814_;
  assign new_n816_ = ~new_n504_ & new_n517_;
  assign new_n817_ = new_n504_ & ~new_n517_;
  assign new_n818_ = ~new_n816_ & ~new_n817_;
  assign new_n819_ = new_n815_ & new_n818_;
  assign new_n820_ = ~new_n815_ & ~new_n818_;
  assign new_n821_ = ~new_n819_ & ~new_n820_;
  assign new_n822_ = new_n492_ & ~new_n821_;
  assign new_n823_ = ~new_n492_ & new_n821_;
  assign new_n824_ = ~new_n822_ & ~new_n823_;
  assign new_n825_ = pi110 & ~pi123;
  assign new_n826_ = pi111 & pi123;
  assign new_n827_ = ~new_n825_ & ~new_n826_;
  assign new_n828_ = new_n477_ & ~new_n827_;
  assign new_n829_ = ~new_n477_ & new_n827_;
  assign new_n830_ = ~new_n828_ & ~new_n829_;
  assign new_n831_ = new_n465_ & new_n830_;
  assign new_n832_ = ~new_n465_ & ~new_n830_;
  assign new_n833_ = ~new_n831_ & ~new_n832_;
  assign new_n834_ = new_n471_ & ~new_n485_;
  assign new_n835_ = ~new_n471_ & new_n485_;
  assign new_n836_ = ~new_n834_ & ~new_n835_;
  assign new_n837_ = new_n833_ & ~new_n836_;
  assign new_n838_ = ~new_n833_ & new_n836_;
  assign new_n839_ = ~new_n837_ & ~new_n838_;
  assign new_n840_ = new_n824_ & new_n839_;
  assign new_n841_ = ~new_n824_ & ~new_n839_;
  assign po37 = new_n840_ | new_n841_;
  assign new_n843_ = pi001 & new_n523_;
  assign new_n844_ = ~new_n634_ & ~new_n843_;
  assign new_n845_ = ~new_n472_ & new_n844_;
  assign new_n846_ = ~new_n473_ & ~new_n845_;
  assign new_n847_ = new_n480_ & ~new_n846_;
  assign new_n848_ = ~new_n480_ & new_n846_;
  assign new_n849_ = ~new_n847_ & ~new_n848_;
  assign new_n850_ = new_n474_ & ~new_n844_;
  assign new_n851_ = ~new_n474_ & new_n844_;
  assign new_n852_ = ~new_n850_ & ~new_n851_;
  assign new_n853_ = ~new_n677_ & ~new_n780_;
  assign new_n854_ = ~new_n772_ & new_n853_;
  assign new_n855_ = new_n761_ & new_n854_;
  assign new_n856_ = new_n753_ & new_n855_;
  assign new_n857_ = ~new_n852_ & new_n856_;
  assign new_n858_ = new_n849_ & new_n857_;
  assign new_n859_ = new_n482_ & ~new_n844_;
  assign new_n860_ = ~new_n639_ & ~new_n859_;
  assign new_n861_ = new_n488_ & ~new_n860_;
  assign new_n862_ = ~new_n488_ & new_n860_;
  assign new_n863_ = ~new_n861_ & ~new_n862_;
  assign new_n864_ = new_n637_ & new_n844_;
  assign new_n865_ = ~new_n473_ & new_n480_;
  assign new_n866_ = ~new_n478_ & ~new_n865_;
  assign new_n867_ = ~new_n864_ & ~new_n866_;
  assign new_n868_ = new_n468_ & ~new_n867_;
  assign new_n869_ = ~new_n468_ & new_n867_;
  assign new_n870_ = ~new_n868_ & ~new_n869_;
  assign new_n871_ = ~new_n863_ & new_n870_;
  assign po38 = new_n858_ & new_n871_;
  assign new_n873_ = new_n572_ & ~new_n684_;
  assign new_n874_ = ~new_n572_ & new_n684_;
  assign new_n875_ = ~new_n873_ & ~new_n874_;
  assign new_n876_ = ~new_n657_ & new_n668_;
  assign new_n877_ = new_n729_ & new_n876_;
  assign new_n878_ = new_n719_ & new_n877_;
  assign new_n879_ = new_n707_ & new_n878_;
  assign new_n880_ = ~new_n875_ & new_n879_;
  assign new_n881_ = po26 & new_n880_;
  assign new_n882_ = ~new_n570_ & new_n684_;
  assign new_n883_ = ~new_n571_ & ~new_n882_;
  assign new_n884_ = new_n566_ & ~new_n883_;
  assign new_n885_ = ~new_n566_ & new_n883_;
  assign new_n886_ = ~new_n884_ & ~new_n885_;
  assign new_n887_ = ~new_n559_ & new_n686_;
  assign new_n888_ = new_n559_ & ~new_n686_;
  assign new_n889_ = ~new_n887_ & ~new_n888_;
  assign new_n890_ = new_n886_ & new_n889_;
  assign po39 = new_n881_ & new_n890_;
  assign new_n892_ = pi155 & ~pi156;
  assign new_n893_ = ~po25 & new_n892_;
  assign new_n894_ = ~pi155 & ~pi156;
  assign new_n895_ = ~po23 & new_n894_;
  assign new_n896_ = ~pi080 & pi155;
  assign new_n897_ = ~pi079 & ~pi155;
  assign new_n898_ = pi156 & ~new_n897_;
  assign new_n899_ = ~new_n896_ & new_n898_;
  assign new_n900_ = ~new_n895_ & ~new_n899_;
  assign new_n901_ = ~new_n893_ & new_n900_;
  assign po40 = pi063 & ~new_n901_;
  assign new_n903_ = pi157 & ~pi158;
  assign new_n904_ = ~po25 & new_n903_;
  assign new_n905_ = ~pi157 & ~pi158;
  assign new_n906_ = ~po23 & new_n905_;
  assign new_n907_ = ~pi080 & pi157;
  assign new_n908_ = ~pi079 & ~pi157;
  assign new_n909_ = pi158 & ~new_n908_;
  assign new_n910_ = ~new_n907_ & new_n909_;
  assign new_n911_ = ~new_n906_ & ~new_n910_;
  assign new_n912_ = ~new_n904_ & new_n911_;
  assign po41 = pi063 & ~new_n912_;
  assign new_n914_ = new_n692_ & ~po32;
  assign new_n915_ = new_n694_ & ~po28;
  assign new_n916_ = ~pi013 & pi170;
  assign new_n917_ = ~pi015 & ~pi170;
  assign new_n918_ = pi169 & ~new_n917_;
  assign new_n919_ = ~new_n916_ & new_n918_;
  assign new_n920_ = ~new_n915_ & ~new_n919_;
  assign po42 = new_n914_ | ~new_n920_;
  assign new_n922_ = new_n692_ & ~po33;
  assign new_n923_ = new_n694_ & ~po29;
  assign new_n924_ = ~pi005 & pi170;
  assign new_n925_ = ~pi026 & ~pi170;
  assign new_n926_ = pi169 & ~new_n925_;
  assign new_n927_ = ~new_n924_ & new_n926_;
  assign new_n928_ = ~new_n923_ & ~new_n927_;
  assign po43 = new_n922_ | ~new_n928_;
  assign new_n930_ = new_n692_ & ~po34;
  assign new_n931_ = new_n694_ & ~po30;
  assign new_n932_ = ~pi004 & pi170;
  assign new_n933_ = ~pi025 & ~pi170;
  assign new_n934_ = pi169 & ~new_n933_;
  assign new_n935_ = ~new_n932_ & new_n934_;
  assign new_n936_ = ~new_n931_ & ~new_n935_;
  assign po44 = new_n930_ | ~new_n936_;
  assign new_n938_ = new_n692_ & ~po35;
  assign new_n939_ = ~po24 & new_n694_;
  assign new_n940_ = ~pi024 & pi170;
  assign new_n941_ = ~pi023 & ~pi170;
  assign new_n942_ = pi169 & ~new_n941_;
  assign new_n943_ = ~new_n940_ & new_n942_;
  assign new_n944_ = ~new_n939_ & ~new_n943_;
  assign po45 = new_n938_ | ~new_n944_;
  assign new_n946_ = new_n735_ & ~po32;
  assign new_n947_ = ~po28 & new_n737_;
  assign new_n948_ = ~pi013 & pi171;
  assign new_n949_ = ~pi015 & ~pi171;
  assign new_n950_ = pi172 & ~new_n949_;
  assign new_n951_ = ~new_n948_ & new_n950_;
  assign new_n952_ = ~new_n947_ & ~new_n951_;
  assign po46 = new_n946_ | ~new_n952_;
  assign new_n954_ = new_n735_ & ~po33;
  assign new_n955_ = ~po29 & new_n737_;
  assign new_n956_ = ~pi005 & pi171;
  assign new_n957_ = ~pi026 & ~pi171;
  assign new_n958_ = pi172 & ~new_n957_;
  assign new_n959_ = ~new_n956_ & new_n958_;
  assign new_n960_ = ~new_n955_ & ~new_n959_;
  assign po47 = new_n954_ | ~new_n960_;
  assign new_n962_ = new_n735_ & ~po34;
  assign new_n963_ = ~po30 & new_n737_;
  assign new_n964_ = ~pi004 & pi171;
  assign new_n965_ = ~pi025 & ~pi171;
  assign new_n966_ = pi172 & ~new_n965_;
  assign new_n967_ = ~new_n964_ & new_n966_;
  assign new_n968_ = ~new_n963_ & ~new_n967_;
  assign po48 = new_n962_ | ~new_n968_;
  assign new_n970_ = new_n735_ & ~po35;
  assign new_n971_ = ~po24 & new_n737_;
  assign new_n972_ = ~pi024 & pi171;
  assign new_n973_ = ~pi023 & ~pi171;
  assign new_n974_ = pi172 & ~new_n973_;
  assign new_n975_ = ~new_n972_ & new_n974_;
  assign new_n976_ = ~new_n971_ & ~new_n975_;
  assign po49 = new_n970_ | ~new_n976_;
  assign new_n978_ = ~po32 & new_n892_;
  assign new_n979_ = ~po28 & new_n894_;
  assign new_n980_ = ~pi075 & pi155;
  assign new_n981_ = ~pi085 & ~pi155;
  assign new_n982_ = pi156 & ~new_n981_;
  assign new_n983_ = ~new_n980_ & new_n982_;
  assign new_n984_ = ~new_n979_ & ~new_n983_;
  assign new_n985_ = ~new_n978_ & new_n984_;
  assign po50 = pi063 & ~new_n985_;
  assign new_n987_ = ~po35 & new_n892_;
  assign new_n988_ = ~po24 & new_n894_;
  assign new_n989_ = ~pi071 & pi155;
  assign new_n990_ = ~pi081 & ~pi155;
  assign new_n991_ = pi156 & ~new_n990_;
  assign new_n992_ = ~new_n989_ & new_n991_;
  assign new_n993_ = ~new_n988_ & ~new_n992_;
  assign new_n994_ = ~new_n987_ & new_n993_;
  assign po51 = pi063 & ~new_n994_;
  assign new_n996_ = ~po34 & new_n892_;
  assign new_n997_ = ~po30 & new_n894_;
  assign new_n998_ = ~pi069 & pi155;
  assign new_n999_ = ~pi070 & ~pi155;
  assign new_n1000_ = pi156 & ~new_n999_;
  assign new_n1001_ = ~new_n998_ & new_n1000_;
  assign new_n1002_ = ~new_n997_ & ~new_n1001_;
  assign new_n1003_ = ~new_n996_ & new_n1002_;
  assign po52 = pi063 & ~new_n1003_;
  assign new_n1005_ = ~po33 & new_n892_;
  assign new_n1006_ = ~po29 & new_n894_;
  assign new_n1007_ = ~pi067 & pi155;
  assign new_n1008_ = ~pi068 & ~pi155;
  assign new_n1009_ = pi156 & ~new_n1008_;
  assign new_n1010_ = ~new_n1007_ & new_n1009_;
  assign new_n1011_ = ~new_n1006_ & ~new_n1010_;
  assign new_n1012_ = ~new_n1005_ & new_n1011_;
  assign po53 = pi063 & ~new_n1012_;
  assign new_n1014_ = ~po32 & new_n903_;
  assign new_n1015_ = ~po28 & new_n905_;
  assign new_n1016_ = ~pi075 & pi157;
  assign new_n1017_ = ~pi085 & ~pi157;
  assign new_n1018_ = pi158 & ~new_n1017_;
  assign new_n1019_ = ~new_n1016_ & new_n1018_;
  assign new_n1020_ = ~new_n1015_ & ~new_n1019_;
  assign new_n1021_ = ~new_n1014_ & new_n1020_;
  assign po54 = pi063 & ~new_n1021_;
  assign new_n1023_ = ~po35 & new_n903_;
  assign new_n1024_ = ~po24 & new_n905_;
  assign new_n1025_ = ~pi071 & pi157;
  assign new_n1026_ = ~pi081 & ~pi157;
  assign new_n1027_ = pi158 & ~new_n1026_;
  assign new_n1028_ = ~new_n1025_ & new_n1027_;
  assign new_n1029_ = ~new_n1024_ & ~new_n1028_;
  assign new_n1030_ = ~new_n1023_ & new_n1029_;
  assign po55 = pi063 & ~new_n1030_;
  assign new_n1032_ = ~po34 & new_n903_;
  assign new_n1033_ = ~po30 & new_n905_;
  assign new_n1034_ = ~pi069 & pi157;
  assign new_n1035_ = ~pi070 & ~pi157;
  assign new_n1036_ = pi158 & ~new_n1035_;
  assign new_n1037_ = ~new_n1034_ & new_n1036_;
  assign new_n1038_ = ~new_n1033_ & ~new_n1037_;
  assign new_n1039_ = ~new_n1032_ & new_n1038_;
  assign po56 = pi063 & ~new_n1039_;
  assign new_n1041_ = ~po33 & new_n903_;
  assign new_n1042_ = ~po29 & new_n905_;
  assign new_n1043_ = ~pi067 & pi157;
  assign new_n1044_ = ~pi068 & ~pi157;
  assign new_n1045_ = pi158 & ~new_n1044_;
  assign new_n1046_ = ~new_n1043_ & new_n1045_;
  assign new_n1047_ = ~new_n1042_ & ~new_n1046_;
  assign new_n1048_ = ~new_n1041_ & new_n1047_;
  assign po57 = pi063 & ~new_n1048_;
  assign new_n1050_ = pi167 & ~po26;
  assign new_n1051_ = ~pi060 & ~new_n556_;
  assign new_n1052_ = pi060 & new_n556_;
  assign new_n1053_ = ~new_n1051_ & ~new_n1052_;
  assign new_n1054_ = ~pi167 & ~new_n1053_;
  assign new_n1055_ = pi168 & ~new_n1054_;
  assign new_n1056_ = ~new_n1050_ & new_n1055_;
  assign new_n1057_ = pi061 & pi175;
  assign new_n1058_ = ~pi167 & new_n338_;
  assign new_n1059_ = pi053 & pi167;
  assign new_n1060_ = ~pi168 & ~new_n1059_;
  assign new_n1061_ = ~new_n1058_ & new_n1060_;
  assign new_n1062_ = ~new_n1057_ & ~new_n1061_;
  assign po58 = ~new_n1056_ & new_n1062_;
  assign new_n1064_ = ~pi060 & ~new_n887_;
  assign new_n1065_ = pi060 & new_n887_;
  assign po59 = new_n1064_ | new_n1065_;
  assign new_n1067_ = new_n659_ & ~po26;
  assign new_n1068_ = new_n338_ & new_n661_;
  assign new_n1069_ = pi053 & new_n663_;
  assign new_n1070_ = ~new_n1068_ & ~new_n1069_;
  assign po60 = ~new_n1067_ & new_n1070_;
  assign new_n1072_ = new_n659_ & ~new_n889_;
  assign new_n1073_ = ~new_n335_ & new_n661_;
  assign new_n1074_ = pi051 & new_n663_;
  assign new_n1075_ = ~new_n1073_ & ~new_n1074_;
  assign po61 = ~new_n1072_ & new_n1075_;
  assign new_n1077_ = new_n659_ & ~new_n886_;
  assign new_n1078_ = ~new_n322_ & new_n661_;
  assign new_n1079_ = pi046 & new_n663_;
  assign new_n1080_ = ~new_n1078_ & ~new_n1079_;
  assign po62 = ~new_n1077_ & new_n1080_;
  assign new_n1082_ = new_n659_ & new_n875_;
  assign new_n1083_ = ~new_n313_ & new_n661_;
  assign new_n1084_ = pi042 & new_n663_;
  assign new_n1085_ = ~new_n1083_ & ~new_n1084_;
  assign po63 = ~new_n1082_ & new_n1085_;
  assign new_n1087_ = pi098 & pi152;
  assign new_n1088_ = po00 & new_n1087_;
  assign new_n1089_ = ~po05 & new_n1088_;
  assign new_n1090_ = ~po19 & new_n1089_;
  assign new_n1091_ = ~po20 & new_n1090_;
  assign new_n1092_ = ~po37 & new_n1091_;
  assign po64 = ~po36 & new_n1092_;
  assign new_n1094_ = new_n659_ & new_n863_;
  assign new_n1095_ = ~new_n429_ & new_n661_;
  assign new_n1096_ = pi045 & new_n663_;
  assign new_n1097_ = ~new_n1095_ & ~new_n1096_;
  assign po65 = ~new_n1094_ & new_n1097_;
  assign new_n1099_ = new_n659_ & ~new_n870_;
  assign new_n1100_ = new_n389_ & new_n661_;
  assign new_n1101_ = pi044 & new_n663_;
  assign new_n1102_ = ~new_n1100_ & ~new_n1101_;
  assign po66 = ~new_n1099_ & new_n1102_;
  assign new_n1104_ = new_n659_ & ~new_n849_;
  assign new_n1105_ = new_n379_ & new_n661_;
  assign new_n1106_ = pi019 & new_n663_;
  assign new_n1107_ = ~new_n1105_ & ~new_n1106_;
  assign po67 = ~new_n1104_ & new_n1107_;
  assign new_n1109_ = new_n659_ & new_n852_;
  assign new_n1110_ = new_n439_ & new_n661_;
  assign new_n1111_ = pi043 & new_n663_;
  assign new_n1112_ = ~new_n1110_ & ~new_n1111_;
  assign po68 = ~new_n1109_ & new_n1112_;
  assign new_n1114_ = new_n735_ & ~po65;
  assign new_n1115_ = new_n737_ & ~po60;
  assign new_n1116_ = ~pi040 & pi171;
  assign new_n1117_ = ~pi041 & ~pi171;
  assign new_n1118_ = pi172 & ~new_n1117_;
  assign new_n1119_ = ~new_n1116_ & new_n1118_;
  assign new_n1120_ = ~new_n1115_ & ~new_n1119_;
  assign po69 = new_n1114_ | ~new_n1120_;
  assign new_n1122_ = new_n692_ & ~po65;
  assign new_n1123_ = new_n694_ & ~po60;
  assign new_n1124_ = ~pi040 & pi170;
  assign new_n1125_ = ~pi041 & ~pi170;
  assign new_n1126_ = pi169 & ~new_n1125_;
  assign new_n1127_ = ~new_n1124_ & new_n1126_;
  assign new_n1128_ = ~new_n1123_ & ~new_n1127_;
  assign po70 = new_n1122_ | ~new_n1128_;
  assign new_n1130_ = new_n692_ & ~po66;
  assign new_n1131_ = new_n694_ & ~po61;
  assign new_n1132_ = ~pi017 & pi170;
  assign new_n1133_ = ~pi016 & ~pi170;
  assign new_n1134_ = pi169 & ~new_n1133_;
  assign new_n1135_ = ~new_n1132_ & new_n1134_;
  assign new_n1136_ = ~new_n1131_ & ~new_n1135_;
  assign po71 = new_n1130_ | ~new_n1136_;
  assign new_n1138_ = new_n692_ & ~po67;
  assign new_n1139_ = new_n694_ & ~po62;
  assign new_n1140_ = ~pi039 & pi170;
  assign new_n1141_ = ~pi038 & ~pi170;
  assign new_n1142_ = pi169 & ~new_n1141_;
  assign new_n1143_ = ~new_n1140_ & new_n1142_;
  assign new_n1144_ = ~new_n1139_ & ~new_n1143_;
  assign po72 = new_n1138_ | ~new_n1144_;
  assign new_n1146_ = new_n692_ & ~po68;
  assign new_n1147_ = new_n694_ & ~po63;
  assign new_n1148_ = ~pi014 & pi170;
  assign new_n1149_ = ~pi035 & ~pi170;
  assign new_n1150_ = pi169 & ~new_n1149_;
  assign new_n1151_ = ~new_n1148_ & new_n1150_;
  assign new_n1152_ = ~new_n1147_ & ~new_n1151_;
  assign po73 = new_n1146_ | ~new_n1152_;
  assign new_n1154_ = new_n735_ & ~po66;
  assign new_n1155_ = new_n737_ & ~po61;
  assign new_n1156_ = ~pi017 & pi171;
  assign new_n1157_ = ~pi016 & ~pi171;
  assign new_n1158_ = pi172 & ~new_n1157_;
  assign new_n1159_ = ~new_n1156_ & new_n1158_;
  assign new_n1160_ = ~new_n1155_ & ~new_n1159_;
  assign po74 = new_n1154_ | ~new_n1160_;
  assign new_n1162_ = new_n735_ & ~po67;
  assign new_n1163_ = new_n737_ & ~po62;
  assign new_n1164_ = ~pi039 & pi171;
  assign new_n1165_ = ~pi038 & ~pi171;
  assign new_n1166_ = pi172 & ~new_n1165_;
  assign new_n1167_ = ~new_n1164_ & new_n1166_;
  assign new_n1168_ = ~new_n1163_ & ~new_n1167_;
  assign po75 = new_n1162_ | ~new_n1168_;
  assign new_n1170_ = new_n735_ & ~po68;
  assign new_n1171_ = new_n737_ & ~po63;
  assign new_n1172_ = ~pi014 & pi171;
  assign new_n1173_ = ~pi035 & ~pi171;
  assign new_n1174_ = pi172 & ~new_n1173_;
  assign new_n1175_ = ~new_n1172_ & new_n1174_;
  assign new_n1176_ = ~new_n1171_ & ~new_n1175_;
  assign po76 = new_n1170_ | ~new_n1176_;
  assign new_n1178_ = new_n892_ & ~po68;
  assign new_n1179_ = new_n894_ & ~po63;
  assign new_n1180_ = ~pi076 & pi155;
  assign new_n1181_ = ~pi086 & ~pi155;
  assign new_n1182_ = pi156 & ~new_n1181_;
  assign new_n1183_ = ~new_n1180_ & new_n1182_;
  assign new_n1184_ = ~new_n1179_ & ~new_n1183_;
  assign new_n1185_ = ~new_n1178_ & new_n1184_;
  assign po77 = pi063 & ~new_n1185_;
  assign new_n1187_ = new_n892_ & ~po67;
  assign new_n1188_ = new_n894_ & ~po62;
  assign new_n1189_ = ~pi074 & pi155;
  assign new_n1190_ = ~pi084 & ~pi155;
  assign new_n1191_ = pi156 & ~new_n1190_;
  assign new_n1192_ = ~new_n1189_ & new_n1191_;
  assign new_n1193_ = ~new_n1188_ & ~new_n1192_;
  assign new_n1194_ = ~new_n1187_ & new_n1193_;
  assign po78 = pi063 & ~new_n1194_;
  assign new_n1196_ = new_n892_ & ~po66;
  assign new_n1197_ = new_n894_ & ~po61;
  assign new_n1198_ = ~pi073 & pi155;
  assign new_n1199_ = ~pi083 & ~pi155;
  assign new_n1200_ = pi156 & ~new_n1199_;
  assign new_n1201_ = ~new_n1198_ & new_n1200_;
  assign new_n1202_ = ~new_n1197_ & ~new_n1201_;
  assign new_n1203_ = ~new_n1196_ & new_n1202_;
  assign po79 = pi063 & ~new_n1203_;
  assign new_n1205_ = new_n892_ & ~po65;
  assign new_n1206_ = new_n894_ & ~po60;
  assign new_n1207_ = ~pi072 & pi155;
  assign new_n1208_ = ~pi082 & ~pi155;
  assign new_n1209_ = pi156 & ~new_n1208_;
  assign new_n1210_ = ~new_n1207_ & new_n1209_;
  assign new_n1211_ = ~new_n1206_ & ~new_n1210_;
  assign new_n1212_ = ~new_n1205_ & new_n1211_;
  assign po80 = pi063 & ~new_n1212_;
  assign new_n1214_ = new_n903_ & ~po68;
  assign new_n1215_ = new_n905_ & ~po63;
  assign new_n1216_ = ~pi076 & pi157;
  assign new_n1217_ = ~pi086 & ~pi157;
  assign new_n1218_ = pi158 & ~new_n1217_;
  assign new_n1219_ = ~new_n1216_ & new_n1218_;
  assign new_n1220_ = ~new_n1215_ & ~new_n1219_;
  assign new_n1221_ = ~new_n1214_ & new_n1220_;
  assign po81 = pi063 & ~new_n1221_;
  assign new_n1223_ = new_n903_ & ~po67;
  assign new_n1224_ = new_n905_ & ~po62;
  assign new_n1225_ = ~pi074 & pi157;
  assign new_n1226_ = ~pi084 & ~pi157;
  assign new_n1227_ = pi158 & ~new_n1226_;
  assign new_n1228_ = ~new_n1225_ & new_n1227_;
  assign new_n1229_ = ~new_n1224_ & ~new_n1228_;
  assign new_n1230_ = ~new_n1223_ & new_n1229_;
  assign po82 = pi063 & ~new_n1230_;
  assign new_n1232_ = new_n903_ & ~po66;
  assign new_n1233_ = new_n905_ & ~po61;
  assign new_n1234_ = ~pi073 & pi157;
  assign new_n1235_ = ~pi083 & ~pi157;
  assign new_n1236_ = pi158 & ~new_n1235_;
  assign new_n1237_ = ~new_n1234_ & new_n1236_;
  assign new_n1238_ = ~new_n1233_ & ~new_n1237_;
  assign new_n1239_ = ~new_n1232_ & new_n1238_;
  assign po83 = pi063 & ~new_n1239_;
  assign new_n1241_ = new_n903_ & ~po65;
  assign new_n1242_ = new_n905_ & ~po60;
  assign new_n1243_ = ~pi072 & pi157;
  assign new_n1244_ = ~pi082 & ~pi157;
  assign new_n1245_ = pi158 & ~new_n1244_;
  assign new_n1246_ = ~new_n1243_ & new_n1245_;
  assign new_n1247_ = ~new_n1242_ & ~new_n1246_;
  assign new_n1248_ = ~new_n1241_ & new_n1247_;
  assign po84 = pi063 & ~new_n1248_;
  assign new_n1250_ = ~pi050 & ~pi173;
  assign new_n1251_ = ~new_n335_ & new_n338_;
  assign new_n1252_ = ~new_n339_ & ~new_n1251_;
  assign new_n1253_ = pi099 & pi127;
  assign new_n1254_ = pi100 & ~pi127;
  assign new_n1255_ = pi149 & ~new_n1254_;
  assign new_n1256_ = ~new_n1253_ & new_n1255_;
  assign new_n1257_ = ~pi097 & pi127;
  assign new_n1258_ = ~pi101 & ~pi127;
  assign new_n1259_ = ~pi149 & ~new_n1258_;
  assign new_n1260_ = ~new_n1257_ & new_n1259_;
  assign new_n1261_ = ~new_n1256_ & ~new_n1260_;
  assign new_n1262_ = pi099 & pi125;
  assign new_n1263_ = pi100 & ~pi125;
  assign new_n1264_ = pi148 & ~new_n1263_;
  assign new_n1265_ = ~new_n1262_ & new_n1264_;
  assign new_n1266_ = ~pi097 & pi125;
  assign new_n1267_ = ~pi101 & ~pi125;
  assign new_n1268_ = ~pi148 & ~new_n1267_;
  assign new_n1269_ = ~new_n1266_ & new_n1268_;
  assign new_n1270_ = ~new_n1265_ & ~new_n1269_;
  assign new_n1271_ = ~new_n1261_ & new_n1270_;
  assign new_n1272_ = new_n1261_ & ~new_n1270_;
  assign new_n1273_ = ~new_n1271_ & ~new_n1272_;
  assign new_n1274_ = ~pi099 & pi147;
  assign new_n1275_ = pi097 & ~pi147;
  assign new_n1276_ = ~new_n1274_ & ~new_n1275_;
  assign new_n1277_ = new_n1273_ & ~new_n1276_;
  assign new_n1278_ = ~new_n1273_ & new_n1276_;
  assign new_n1279_ = ~new_n1277_ & ~new_n1278_;
  assign new_n1280_ = ~new_n313_ & ~new_n322_;
  assign new_n1281_ = ~new_n323_ & ~new_n1280_;
  assign new_n1282_ = pi099 & pi120;
  assign new_n1283_ = pi100 & ~pi120;
  assign new_n1284_ = pi146 & ~new_n1283_;
  assign new_n1285_ = ~new_n1282_ & new_n1284_;
  assign new_n1286_ = ~pi097 & pi120;
  assign new_n1287_ = ~pi101 & ~pi120;
  assign new_n1288_ = ~pi146 & ~new_n1287_;
  assign new_n1289_ = ~new_n1286_ & new_n1288_;
  assign new_n1290_ = ~new_n1285_ & ~new_n1289_;
  assign new_n1291_ = ~new_n342_ & new_n1290_;
  assign new_n1292_ = new_n342_ & ~new_n1290_;
  assign new_n1293_ = ~new_n1291_ & ~new_n1292_;
  assign new_n1294_ = new_n1281_ & ~new_n1293_;
  assign new_n1295_ = ~new_n1281_ & new_n1293_;
  assign new_n1296_ = ~new_n1294_ & ~new_n1295_;
  assign new_n1297_ = ~new_n1279_ & new_n1296_;
  assign new_n1298_ = new_n1279_ & ~new_n1296_;
  assign new_n1299_ = ~new_n1297_ & ~new_n1298_;
  assign new_n1300_ = ~new_n1252_ & ~new_n1299_;
  assign new_n1301_ = new_n1252_ & new_n1299_;
  assign new_n1302_ = ~pi173 & ~new_n1301_;
  assign new_n1303_ = ~new_n1300_ & new_n1302_;
  assign new_n1304_ = ~pi174 & ~new_n1303_;
  assign new_n1305_ = ~new_n1250_ & ~new_n1304_;
  assign new_n1306_ = pi174 & ~new_n1305_;
  assign new_n1307_ = pi159 & new_n553_;
  assign new_n1308_ = new_n650_ & ~new_n1307_;
  assign new_n1309_ = new_n559_ & new_n565_;
  assign new_n1310_ = new_n559_ & new_n652_;
  assign new_n1311_ = new_n566_ & ~new_n1310_;
  assign new_n1312_ = ~new_n1309_ & ~new_n1311_;
  assign new_n1313_ = new_n570_ & new_n1312_;
  assign new_n1314_ = ~new_n570_ & ~new_n1312_;
  assign new_n1315_ = ~new_n573_ & ~new_n1314_;
  assign new_n1316_ = ~new_n1313_ & new_n1315_;
  assign new_n1317_ = ~new_n1308_ & ~new_n1316_;
  assign new_n1318_ = new_n571_ & ~new_n1312_;
  assign new_n1319_ = ~new_n571_ & new_n1312_;
  assign new_n1320_ = ~new_n1318_ & ~new_n1319_;
  assign new_n1321_ = new_n1308_ & new_n1320_;
  assign new_n1322_ = ~new_n1317_ & ~new_n1321_;
  assign new_n1323_ = ~new_n544_ & ~new_n550_;
  assign new_n1324_ = ~new_n551_ & ~new_n1323_;
  assign new_n1325_ = new_n530_ & ~new_n715_;
  assign new_n1326_ = ~new_n530_ & new_n715_;
  assign new_n1327_ = ~new_n1325_ & ~new_n1326_;
  assign new_n1328_ = ~new_n534_ & new_n539_;
  assign new_n1329_ = new_n534_ & ~new_n539_;
  assign new_n1330_ = ~new_n1328_ & ~new_n1329_;
  assign new_n1331_ = new_n702_ & ~new_n1330_;
  assign new_n1332_ = ~new_n702_ & new_n1330_;
  assign new_n1333_ = ~new_n1331_ & ~new_n1332_;
  assign new_n1334_ = ~new_n1327_ & new_n1333_;
  assign new_n1335_ = new_n1327_ & ~new_n1333_;
  assign new_n1336_ = pi159 & ~new_n1335_;
  assign new_n1337_ = ~new_n1334_ & new_n1336_;
  assign new_n1338_ = ~new_n530_ & new_n648_;
  assign new_n1339_ = ~new_n649_ & ~new_n1338_;
  assign new_n1340_ = ~new_n535_ & ~new_n1328_;
  assign new_n1341_ = new_n646_ & ~new_n1340_;
  assign new_n1342_ = ~new_n646_ & new_n1340_;
  assign new_n1343_ = ~new_n1341_ & ~new_n1342_;
  assign new_n1344_ = ~new_n1339_ & ~new_n1343_;
  assign new_n1345_ = new_n1339_ & new_n1343_;
  assign new_n1346_ = ~pi159 & ~new_n1345_;
  assign new_n1347_ = ~new_n1344_ & new_n1346_;
  assign new_n1348_ = ~new_n1337_ & ~new_n1347_;
  assign new_n1349_ = new_n689_ & ~new_n1348_;
  assign new_n1350_ = ~new_n689_ & new_n1348_;
  assign new_n1351_ = ~new_n1349_ & ~new_n1350_;
  assign new_n1352_ = ~new_n1324_ & new_n1351_;
  assign new_n1353_ = new_n1324_ & ~new_n1351_;
  assign new_n1354_ = ~new_n1352_ & ~new_n1353_;
  assign new_n1355_ = ~new_n1322_ & ~new_n1354_;
  assign new_n1356_ = new_n1322_ & new_n1354_;
  assign new_n1357_ = pi173 & ~new_n1356_;
  assign new_n1358_ = ~new_n1355_ & new_n1357_;
  assign new_n1359_ = new_n1304_ & ~new_n1358_;
  assign po85 = ~new_n1306_ & ~new_n1359_;
  assign new_n1361_ = ~pi048 & ~pi173;
  assign new_n1362_ = pi099 & pi102;
  assign new_n1363_ = pi100 & ~pi102;
  assign new_n1364_ = pi136 & ~new_n1363_;
  assign new_n1365_ = ~new_n1362_ & new_n1364_;
  assign new_n1366_ = ~pi097 & pi102;
  assign new_n1367_ = ~pi101 & ~pi102;
  assign new_n1368_ = ~pi136 & ~new_n1367_;
  assign new_n1369_ = ~new_n1366_ & new_n1368_;
  assign new_n1370_ = ~new_n1365_ & ~new_n1369_;
  assign new_n1371_ = pi099 & pi108;
  assign new_n1372_ = pi100 & ~pi108;
  assign new_n1373_ = pi134 & ~new_n1372_;
  assign new_n1374_ = ~new_n1371_ & new_n1373_;
  assign new_n1375_ = ~pi097 & pi108;
  assign new_n1376_ = ~pi101 & ~pi108;
  assign new_n1377_ = ~pi134 & ~new_n1376_;
  assign new_n1378_ = ~new_n1375_ & new_n1377_;
  assign new_n1379_ = ~new_n1374_ & ~new_n1378_;
  assign new_n1380_ = ~new_n1370_ & new_n1379_;
  assign new_n1381_ = new_n1370_ & ~new_n1379_;
  assign new_n1382_ = ~new_n1380_ & ~new_n1381_;
  assign new_n1383_ = pi093 & pi097;
  assign new_n1384_ = ~pi093 & pi101;
  assign new_n1385_ = ~pi139 & ~new_n1384_;
  assign new_n1386_ = ~new_n1383_ & new_n1385_;
  assign new_n1387_ = pi099 & new_n434_;
  assign new_n1388_ = pi100 & new_n436_;
  assign new_n1389_ = ~new_n1387_ & ~new_n1388_;
  assign new_n1390_ = ~new_n1386_ & new_n1389_;
  assign new_n1391_ = new_n429_ & ~new_n1390_;
  assign new_n1392_ = ~new_n429_ & new_n1390_;
  assign new_n1393_ = ~new_n1391_ & ~new_n1392_;
  assign new_n1394_ = new_n1382_ & ~new_n1393_;
  assign new_n1395_ = ~new_n1382_ & new_n1393_;
  assign new_n1396_ = ~new_n1394_ & ~new_n1395_;
  assign new_n1397_ = pi099 & pi106;
  assign new_n1398_ = pi100 & ~pi106;
  assign new_n1399_ = pi138 & ~new_n1398_;
  assign new_n1400_ = ~new_n1397_ & new_n1399_;
  assign new_n1401_ = ~pi097 & pi106;
  assign new_n1402_ = ~pi101 & ~pi106;
  assign new_n1403_ = ~pi138 & ~new_n1402_;
  assign new_n1404_ = ~new_n1401_ & new_n1403_;
  assign new_n1405_ = ~new_n1400_ & ~new_n1404_;
  assign new_n1406_ = pi099 & pi104;
  assign new_n1407_ = pi100 & ~pi104;
  assign new_n1408_ = pi137 & ~new_n1407_;
  assign new_n1409_ = ~new_n1406_ & new_n1408_;
  assign new_n1410_ = ~pi097 & pi104;
  assign new_n1411_ = ~pi101 & ~pi104;
  assign new_n1412_ = ~pi137 & ~new_n1411_;
  assign new_n1413_ = ~new_n1410_ & new_n1412_;
  assign new_n1414_ = ~new_n1409_ & ~new_n1413_;
  assign new_n1415_ = ~new_n1405_ & new_n1414_;
  assign new_n1416_ = new_n1405_ & ~new_n1414_;
  assign new_n1417_ = ~new_n1415_ & ~new_n1416_;
  assign new_n1418_ = pi095 & pi097;
  assign new_n1419_ = ~pi095 & pi101;
  assign new_n1420_ = ~pi140 & ~new_n1419_;
  assign new_n1421_ = ~new_n1418_ & new_n1420_;
  assign new_n1422_ = pi099 & new_n414_;
  assign new_n1423_ = pi100 & new_n416_;
  assign new_n1424_ = ~new_n1422_ & ~new_n1423_;
  assign new_n1425_ = ~new_n1421_ & new_n1424_;
  assign new_n1426_ = new_n1417_ & new_n1425_;
  assign new_n1427_ = ~new_n1417_ & ~new_n1425_;
  assign new_n1428_ = ~new_n1426_ & ~new_n1427_;
  assign new_n1429_ = pi089 & pi097;
  assign new_n1430_ = ~pi089 & pi101;
  assign new_n1431_ = ~pi142 & ~new_n1430_;
  assign new_n1432_ = ~new_n1429_ & new_n1431_;
  assign new_n1433_ = pi099 & new_n384_;
  assign new_n1434_ = pi100 & new_n386_;
  assign new_n1435_ = ~new_n1433_ & ~new_n1434_;
  assign new_n1436_ = ~new_n1432_ & new_n1435_;
  assign new_n1437_ = pi091 & pi097;
  assign new_n1438_ = ~pi091 & pi101;
  assign new_n1439_ = ~pi143 & ~new_n1438_;
  assign new_n1440_ = ~new_n1437_ & new_n1439_;
  assign new_n1441_ = pi099 & new_n374_;
  assign new_n1442_ = pi100 & new_n376_;
  assign new_n1443_ = ~new_n1441_ & ~new_n1442_;
  assign new_n1444_ = ~new_n1440_ & new_n1443_;
  assign new_n1445_ = new_n1436_ & ~new_n1444_;
  assign new_n1446_ = ~new_n1436_ & new_n1444_;
  assign new_n1447_ = ~new_n1445_ & ~new_n1446_;
  assign new_n1448_ = new_n1428_ & ~new_n1447_;
  assign new_n1449_ = ~new_n1428_ & new_n1447_;
  assign new_n1450_ = ~new_n1448_ & ~new_n1449_;
  assign new_n1451_ = ~new_n1396_ & new_n1450_;
  assign new_n1452_ = new_n1396_ & ~new_n1450_;
  assign new_n1453_ = ~pi173 & ~new_n1452_;
  assign new_n1454_ = ~new_n1451_ & new_n1453_;
  assign new_n1455_ = ~pi174 & ~new_n1454_;
  assign new_n1456_ = ~new_n1361_ & ~new_n1455_;
  assign new_n1457_ = pi174 & ~new_n1456_;
  assign new_n1458_ = ~new_n514_ & ~new_n520_;
  assign new_n1459_ = ~new_n521_ & ~new_n1458_;
  assign new_n1460_ = new_n468_ & ~new_n1459_;
  assign new_n1461_ = ~new_n468_ & new_n1459_;
  assign new_n1462_ = ~new_n1460_ & ~new_n1461_;
  assign new_n1463_ = pi154 & new_n523_;
  assign new_n1464_ = ~new_n634_ & ~new_n1463_;
  assign new_n1465_ = ~new_n467_ & ~new_n637_;
  assign new_n1466_ = ~new_n638_ & ~new_n1465_;
  assign new_n1467_ = new_n488_ & ~new_n1466_;
  assign new_n1468_ = ~new_n488_ & new_n1466_;
  assign new_n1469_ = ~new_n1467_ & ~new_n1468_;
  assign new_n1470_ = new_n473_ & ~new_n480_;
  assign new_n1471_ = ~new_n865_ & ~new_n1470_;
  assign new_n1472_ = new_n1469_ & new_n1471_;
  assign new_n1473_ = ~new_n1469_ & ~new_n1471_;
  assign new_n1474_ = ~new_n1472_ & ~new_n1473_;
  assign new_n1475_ = new_n1464_ & new_n1474_;
  assign new_n1476_ = ~new_n472_ & ~new_n480_;
  assign new_n1477_ = ~new_n636_ & ~new_n1476_;
  assign new_n1478_ = ~new_n467_ & ~new_n866_;
  assign new_n1479_ = ~new_n639_ & new_n866_;
  assign new_n1480_ = ~new_n1478_ & ~new_n1479_;
  assign new_n1481_ = ~new_n488_ & ~new_n1480_;
  assign new_n1482_ = new_n488_ & new_n1480_;
  assign new_n1483_ = ~new_n1481_ & ~new_n1482_;
  assign new_n1484_ = ~new_n1477_ & ~new_n1483_;
  assign new_n1485_ = new_n1477_ & new_n1483_;
  assign new_n1486_ = ~new_n1464_ & ~new_n1485_;
  assign new_n1487_ = ~new_n1484_ & new_n1486_;
  assign new_n1488_ = ~new_n1475_ & ~new_n1487_;
  assign new_n1489_ = ~new_n505_ & ~new_n627_;
  assign new_n1490_ = ~new_n508_ & new_n1489_;
  assign new_n1491_ = new_n495_ & ~new_n1490_;
  assign new_n1492_ = ~new_n495_ & new_n1490_;
  assign new_n1493_ = ~new_n1491_ & ~new_n1492_;
  assign new_n1494_ = ~new_n627_ & ~new_n778_;
  assign new_n1495_ = ~new_n512_ & new_n746_;
  assign new_n1496_ = ~new_n522_ & ~new_n632_;
  assign new_n1497_ = ~new_n746_ & ~new_n1496_;
  assign new_n1498_ = ~new_n1495_ & ~new_n1497_;
  assign new_n1499_ = new_n1494_ & ~new_n1498_;
  assign new_n1500_ = ~new_n1494_ & new_n1498_;
  assign new_n1501_ = ~new_n1499_ & ~new_n1500_;
  assign new_n1502_ = new_n1493_ & ~new_n1501_;
  assign new_n1503_ = ~new_n1493_ & new_n1501_;
  assign new_n1504_ = ~new_n1502_ & ~new_n1503_;
  assign new_n1505_ = pi154 & ~new_n1504_;
  assign new_n1506_ = new_n507_ & ~new_n632_;
  assign new_n1507_ = ~new_n507_ & new_n632_;
  assign new_n1508_ = ~new_n1506_ & ~new_n1507_;
  assign new_n1509_ = new_n499_ & ~new_n630_;
  assign new_n1510_ = ~new_n499_ & ~new_n519_;
  assign new_n1511_ = ~new_n628_ & new_n1510_;
  assign new_n1512_ = new_n501_ & ~new_n1511_;
  assign new_n1513_ = ~new_n501_ & new_n1511_;
  assign new_n1514_ = ~new_n1512_ & ~new_n1513_;
  assign new_n1515_ = ~new_n1509_ & new_n1514_;
  assign new_n1516_ = new_n495_ & ~new_n1489_;
  assign new_n1517_ = ~new_n495_ & new_n1489_;
  assign new_n1518_ = ~new_n1516_ & ~new_n1517_;
  assign new_n1519_ = ~new_n1515_ & new_n1518_;
  assign new_n1520_ = new_n1515_ & ~new_n1518_;
  assign new_n1521_ = ~new_n1519_ & ~new_n1520_;
  assign new_n1522_ = new_n1508_ & new_n1521_;
  assign new_n1523_ = ~new_n1508_ & ~new_n1521_;
  assign new_n1524_ = ~new_n1522_ & ~new_n1523_;
  assign new_n1525_ = ~pi154 & ~new_n1524_;
  assign new_n1526_ = ~new_n1505_ & ~new_n1525_;
  assign new_n1527_ = new_n1488_ & ~new_n1526_;
  assign new_n1528_ = ~new_n1488_ & new_n1526_;
  assign new_n1529_ = ~new_n1527_ & ~new_n1528_;
  assign new_n1530_ = ~new_n1462_ & new_n1529_;
  assign new_n1531_ = new_n1462_ & ~new_n1529_;
  assign new_n1532_ = pi173 & ~new_n1531_;
  assign new_n1533_ = ~new_n1530_ & new_n1532_;
  assign new_n1534_ = new_n1455_ & ~new_n1533_;
  assign po86 = ~new_n1457_ & ~new_n1534_;
  assign new_n1536_ = pi037 & pi174;
  assign new_n1537_ = ~new_n1534_ & ~new_n1536_;
  assign new_n1538_ = new_n692_ & ~new_n1537_;
  assign new_n1539_ = pi036 & pi174;
  assign new_n1540_ = ~new_n1359_ & ~new_n1539_;
  assign new_n1541_ = new_n694_ & ~new_n1540_;
  assign new_n1542_ = ~pi022 & pi170;
  assign new_n1543_ = ~pi003 & ~pi170;
  assign new_n1544_ = pi169 & ~new_n1543_;
  assign new_n1545_ = ~new_n1542_ & new_n1544_;
  assign new_n1546_ = ~new_n1541_ & ~new_n1545_;
  assign po87 = new_n1538_ | ~new_n1546_;
  assign new_n1548_ = new_n735_ & ~new_n1537_;
  assign new_n1549_ = new_n737_ & ~new_n1540_;
  assign new_n1550_ = ~pi022 & pi171;
  assign new_n1551_ = ~pi003 & ~pi171;
  assign new_n1552_ = pi172 & ~new_n1551_;
  assign new_n1553_ = ~new_n1550_ & new_n1552_;
  assign new_n1554_ = ~new_n1549_ & ~new_n1553_;
  assign po88 = new_n1548_ | ~new_n1554_;
  assign new_n1556_ = new_n892_ & ~new_n1537_;
  assign new_n1557_ = new_n894_ & ~new_n1540_;
  assign new_n1558_ = ~pi078 & pi155;
  assign new_n1559_ = ~pi077 & ~pi155;
  assign new_n1560_ = pi156 & ~new_n1559_;
  assign new_n1561_ = ~new_n1558_ & new_n1560_;
  assign new_n1562_ = ~new_n1557_ & ~new_n1561_;
  assign new_n1563_ = ~new_n1556_ & new_n1562_;
  assign po89 = ~pi063 | new_n1563_;
  assign new_n1565_ = new_n903_ & ~new_n1537_;
  assign new_n1566_ = new_n905_ & ~new_n1540_;
  assign new_n1567_ = ~pi078 & pi157;
  assign new_n1568_ = ~pi077 & ~pi157;
  assign new_n1569_ = pi158 & ~new_n1568_;
  assign new_n1570_ = ~new_n1567_ & new_n1569_;
  assign new_n1571_ = ~new_n1566_ & ~new_n1570_;
  assign new_n1572_ = ~new_n1565_ & new_n1571_;
  assign po90 = ~pi063 | new_n1572_;
endmodule


