// Benchmark "c7552" written by ABC on Thu Jul 14 21:14:45 2022

module c7552 ( 
    G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47,
    G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65,
    G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83,
    G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110,
    G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134,
    G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156,
    G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168,
    G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216,
    G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228,
    G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240,
    \IN-G339 , G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492,
    G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247,
    G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737,
    G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427,
    G4432, G4437, G4526, G4528,
    G339,           
               
               
     G279,    G402, G404, G406, G408, G410,  
    G284,   G292,    G278, G373, G246, G258, 
     G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416,
     G295, G324, G252,  G310, G313, G316, G319, G327, G330, G333,
    G336, G418,  G298, G301, G304, G307, G344, G422,  G419, 
    G359, G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399  );
  input  G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41,
    G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63,
    G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81,
    G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106,
    G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130,
    G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154,
    G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166,
    G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190,
    G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202,
    G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214,
    G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226,
    G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238,
    G239, G240, \IN-G339 , G1197, G1455, G1459, G1462, G1469, G1480, G1486,
    G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239,
    G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729,
    G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420,
    G4427, G4432, G4437, G4526, G4528;
  output G339,           
               
               
     G279,    G402, G404, G406, G408, G410,  
    G284,   G292,    G278, G373, G246, G258, 
     G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416,
     G295, G324, G252,  G310, G313, G316, G319, G327, G330, G333,
    G336, G418,  G298, G301, G304, G307, G344, G422,  G419, 
    G359, G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399;
  wire new_new_n317__, new_new_n318__, new_new_n320__, new_new_n321__,
    new_new_n323__, new_new_n324__, new_new_n326__, new_new_n327__,
    new_new_n330__, new_new_n333__, new_new_n334__, new_new_n335__,
    new_new_n336__, new_new_n337__, new_new_n338__, new_new_n339__,
    new_new_n340__, new_new_n341__, new_new_n343__, new_new_n344__,
    new_new_n345__, new_new_n346__, new_new_n347__, new_new_n348__,
    new_new_n349__, new_new_n350__, new_new_n351__, new_new_n352__,
    new_new_n353__, new_new_n354__, new_new_n355__, new_new_n356__,
    new_new_n357__, new_new_n358__, new_new_n359__, new_new_n360__,
    new_new_n361__, new_new_n362__, new_new_n363__, new_new_n364__,
    new_new_n365__, new_new_n366__, new_new_n367__, new_new_n368__,
    new_new_n369__, new_new_n370__, new_new_n371__, new_new_n372__,
    new_new_n373__, new_new_n374__, new_new_n375__, new_new_n376__,
    new_new_n377__, new_new_n378__, new_new_n379__, new_new_n380__,
    new_new_n381__, new_new_n382__, new_new_n383__, new_new_n384__,
    new_new_n385__, new_new_n386__, new_new_n387__, new_new_n388__,
    new_new_n389__, new_new_n390__, new_new_n391__, new_new_n392__,
    new_new_n393__, new_new_n394__, new_new_n395__, new_new_n396__,
    new_new_n397__, new_new_n398__, new_new_n399__, new_new_n400__,
    new_new_n401__, new_new_n402__, new_new_n403__, new_new_n404__,
    new_new_n405__, new_new_n406__, new_new_n407__, new_new_n408__,
    new_new_n409__, new_new_n410__, new_new_n411__, new_new_n412__,
    new_new_n413__, new_new_n414__, new_new_n415__, new_new_n416__,
    new_new_n417__, new_new_n418__, new_new_n419__, new_new_n420__,
    new_new_n421__, new_new_n422__, new_new_n423__, new_new_n424__,
    new_new_n425__, new_new_n426__, new_new_n427__, new_new_n428__,
    new_new_n429__, new_new_n430__, new_new_n431__, new_new_n432__,
    new_new_n433__, new_new_n434__, new_new_n435__, new_new_n436__,
    new_new_n437__, new_new_n438__, new_new_n439__, new_new_n440__,
    new_new_n441__, new_new_n442__, new_new_n443__, new_new_n444__,
    new_new_n445__, new_new_n446__, new_new_n447__, new_new_n448__,
    new_new_n449__, new_new_n450__, new_new_n451__, new_new_n452__,
    new_new_n453__, new_new_n454__, new_new_n455__, new_new_n456__,
    new_new_n457__, new_new_n458__, new_new_n459__, new_new_n460__,
    new_new_n461__, new_new_n462__, new_new_n463__, new_new_n464__,
    new_new_n465__, new_new_n466__, new_new_n467__, new_new_n468__,
    new_new_n469__, new_new_n470__, new_new_n471__, new_new_n472__,
    new_new_n473__, new_new_n474__, new_new_n475__, new_new_n476__,
    new_new_n477__, new_new_n478__, new_new_n479__, new_new_n480__,
    new_new_n481__, new_new_n482__, new_new_n483__, new_new_n484__,
    new_new_n485__, new_new_n486__, new_new_n487__, new_new_n488__,
    new_new_n489__, new_new_n490__, new_new_n491__, new_new_n492__,
    new_new_n493__, new_new_n494__, new_new_n495__, new_new_n496__,
    new_new_n497__, new_new_n498__, new_new_n499__, new_new_n500__,
    new_new_n501__, new_new_n502__, new_new_n503__, new_new_n504__,
    new_new_n505__, new_new_n506__, new_new_n507__, new_new_n508__,
    new_new_n509__, new_new_n510__, new_new_n511__, new_new_n512__,
    new_new_n513__, new_new_n514__, new_new_n515__, new_new_n516__,
    new_new_n517__, new_new_n518__, new_new_n519__, new_new_n520__,
    new_new_n521__, new_new_n522__, new_new_n523__, new_new_n524__,
    new_new_n525__, new_new_n526__, new_new_n527__, new_new_n528__,
    new_new_n529__, new_new_n530__, new_new_n531__, new_new_n532__,
    new_new_n533__, new_new_n534__, new_new_n535__, new_new_n536__,
    new_new_n537__, new_new_n538__, new_new_n539__, new_new_n540__,
    new_new_n541__, new_new_n542__, new_new_n543__, new_new_n544__,
    new_new_n545__, new_new_n546__, new_new_n547__, new_new_n548__,
    new_new_n549__, new_new_n550__, new_new_n551__, new_new_n552__,
    new_new_n553__, new_new_n554__, new_new_n555__, new_new_n556__,
    new_new_n557__, new_new_n558__, new_new_n559__, new_new_n560__,
    new_new_n561__, new_new_n562__, new_new_n563__, new_new_n564__,
    new_new_n565__, new_new_n566__, new_new_n567__, new_new_n568__,
    new_new_n569__, new_new_n570__, new_new_n571__, new_new_n572__,
    new_new_n573__, new_new_n574__, new_new_n575__, new_new_n576__,
    new_new_n577__, new_new_n578__, new_new_n579__, new_new_n580__,
    new_new_n581__, new_new_n582__, new_new_n583__, new_new_n584__,
    new_new_n585__, new_new_n586__, new_new_n587__, new_new_n588__,
    new_new_n589__, new_new_n590__, new_new_n591__, new_new_n592__,
    new_new_n593__, new_new_n594__, new_new_n595__, new_new_n596__,
    new_new_n597__, new_new_n598__, new_new_n599__, new_new_n600__,
    new_new_n601__, new_new_n602__, new_new_n603__, new_new_n604__,
    new_new_n605__, new_new_n606__, new_new_n607__, new_new_n608__,
    new_new_n609__, new_new_n610__, new_new_n611__, new_new_n612__,
    new_new_n613__, new_new_n614__, new_new_n615__, new_new_n616__,
    new_new_n617__, new_new_n618__, new_new_n619__, new_new_n620__,
    new_new_n621__, new_new_n622__, new_new_n623__, new_new_n624__,
    new_new_n625__, new_new_n626__, new_new_n628__, new_new_n629__,
    new_new_n630__, new_new_n631__, new_new_n632__, new_new_n633__,
    new_new_n634__, new_new_n635__, new_new_n636__, new_new_n637__,
    new_new_n638__, new_new_n639__, new_new_n640__, new_new_n641__,
    new_new_n642__, new_new_n643__, new_new_n644__, new_new_n645__,
    new_new_n646__, new_new_n647__, new_new_n648__, new_new_n649__,
    new_new_n650__, new_new_n651__, new_new_n652__, new_new_n653__,
    new_new_n654__, new_new_n655__, new_new_n656__, new_new_n657__,
    new_new_n658__, new_new_n659__, new_new_n660__, new_new_n661__,
    new_new_n662__, new_new_n663__, new_new_n664__, new_new_n665__,
    new_new_n666__, new_new_n667__, new_new_n668__, new_new_n669__,
    new_new_n670__, new_new_n671__, new_new_n672__, new_new_n673__,
    new_new_n674__, new_new_n675__, new_new_n676__, new_new_n677__,
    new_new_n678__, new_new_n679__, new_new_n680__, new_new_n681__,
    new_new_n682__, new_new_n683__, new_new_n684__, new_new_n685__,
    new_new_n686__, new_new_n687__, new_new_n688__, new_new_n689__,
    new_new_n690__, new_new_n691__, new_new_n692__, new_new_n693__,
    new_new_n694__, new_new_n695__, new_new_n696__, new_new_n697__,
    new_new_n698__, new_new_n699__, new_new_n700__, new_new_n701__,
    new_new_n702__, new_new_n703__, new_new_n704__, new_new_n705__,
    new_new_n706__, new_new_n707__, new_new_n708__, new_new_n709__,
    new_new_n710__, new_new_n711__, new_new_n712__, new_new_n713__,
    new_new_n714__, new_new_n715__, new_new_n716__, new_new_n717__,
    new_new_n718__, new_new_n719__, new_new_n720__, new_new_n721__,
    new_new_n722__, new_new_n723__, new_new_n724__, new_new_n725__,
    new_new_n726__, new_new_n727__, new_new_n728__, new_new_n729__,
    new_new_n730__, new_new_n731__, new_new_n732__, new_new_n733__,
    new_new_n734__, new_new_n735__, new_new_n736__, new_new_n737__,
    new_new_n738__, new_new_n739__, new_new_n740__, new_new_n741__,
    new_new_n742__, new_new_n743__, new_new_n744__, new_new_n745__,
    new_new_n746__, new_new_n747__, new_new_n748__, new_new_n749__,
    new_new_n750__, new_new_n751__, new_new_n752__, new_new_n753__,
    new_new_n754__, new_new_n755__, new_new_n756__, new_new_n757__,
    new_new_n758__, new_new_n759__, new_new_n760__, new_new_n761__,
    new_new_n762__, new_new_n763__, new_new_n764__, new_new_n765__,
    new_new_n766__, new_new_n767__, new_new_n768__, new_new_n769__,
    new_new_n770__, new_new_n771__, new_new_n772__, new_new_n773__,
    new_new_n774__, new_new_n775__, new_new_n776__, new_new_n777__,
    new_new_n778__, new_new_n779__, new_new_n780__, new_new_n781__,
    new_new_n782__, new_new_n783__, new_new_n784__, new_new_n785__,
    new_new_n786__, new_new_n787__, new_new_n788__, new_new_n789__,
    new_new_n790__, new_new_n791__, new_new_n792__, new_new_n793__,
    new_new_n794__, new_new_n795__, new_new_n796__, new_new_n797__,
    new_new_n798__, new_new_n799__, new_new_n800__, new_new_n801__,
    new_new_n802__, new_new_n803__, new_new_n804__, new_new_n805__,
    new_new_n806__, new_new_n807__, new_new_n808__, new_new_n809__,
    new_new_n810__, new_new_n811__, new_new_n812__, new_new_n813__,
    new_new_n814__, new_new_n815__, new_new_n816__, new_new_n817__,
    new_new_n818__, new_new_n819__, new_new_n820__, new_new_n821__,
    new_new_n822__, new_new_n823__, new_new_n824__, new_new_n825__,
    new_new_n826__, new_new_n827__, new_new_n828__, new_new_n829__,
    new_new_n830__, new_new_n831__, new_new_n832__, new_new_n833__,
    new_new_n834__, new_new_n835__, new_new_n836__, new_new_n837__,
    new_new_n838__, new_new_n839__, new_new_n840__, new_new_n841__,
    new_new_n842__, new_new_n843__, new_new_n844__, new_new_n845__,
    new_new_n846__, new_new_n847__, new_new_n848__, new_new_n849__,
    new_new_n850__, new_new_n851__, new_new_n852__, new_new_n853__,
    new_new_n854__, new_new_n855__, new_new_n856__, new_new_n857__,
    new_new_n858__, new_new_n859__, new_new_n860__, new_new_n861__,
    new_new_n862__, new_new_n863__, new_new_n864__, new_new_n865__,
    new_new_n866__, new_new_n867__, new_new_n868__, new_new_n869__,
    new_new_n870__, new_new_n871__, new_new_n872__, new_new_n873__,
    new_new_n874__, new_new_n875__, new_new_n876__, new_new_n877__,
    new_new_n878__, new_new_n879__, new_new_n880__, new_new_n881__,
    new_new_n882__, new_new_n883__, new_new_n884__, new_new_n885__,
    new_new_n886__, new_new_n887__, new_new_n888__, new_new_n889__,
    new_new_n890__, new_new_n891__, new_new_n892__, new_new_n893__,
    new_new_n894__, new_new_n895__, new_new_n896__, new_new_n897__,
    new_new_n898__, new_new_n899__, new_new_n900__, new_new_n901__,
    new_new_n902__, new_new_n903__, new_new_n904__, new_new_n905__,
    new_new_n906__, new_new_n907__, new_new_n908__, new_new_n909__,
    new_new_n910__, new_new_n911__, new_new_n912__, new_new_n913__,
    new_new_n914__, new_new_n915__, new_new_n916__, new_new_n917__,
    new_new_n918__, new_new_n919__, new_new_n920__, new_new_n921__,
    new_new_n922__, new_new_n923__, new_new_n924__, new_new_n925__,
    new_new_n926__, new_new_n927__, new_new_n928__, new_new_n929__,
    new_new_n930__, new_new_n931__, new_new_n932__, new_new_n933__,
    new_new_n934__, new_new_n935__, new_new_n936__, new_new_n937__,
    new_new_n938__, new_new_n939__, new_new_n940__, new_new_n941__,
    new_new_n942__, new_new_n943__, new_new_n944__, new_new_n945__,
    new_new_n946__, new_new_n947__, new_new_n948__, new_new_n949__,
    new_new_n950__, new_new_n951__, new_new_n952__, new_new_n953__,
    new_new_n954__, new_new_n955__, new_new_n956__, new_new_n957__,
    new_new_n958__, new_new_n959__, new_new_n960__, new_new_n961__,
    new_new_n962__, new_new_n963__, new_new_n964__, new_new_n965__,
    new_new_n966__, new_new_n967__, new_new_n968__, new_new_n969__,
    new_new_n971__, new_new_n972__, new_new_n973__, new_new_n974__,
    new_new_n975__, new_new_n976__, new_new_n978__, new_new_n979__,
    new_new_n980__, new_new_n982__, new_new_n983__, new_new_n984__,
    new_new_n985__, new_new_n987__, new_new_n988__, new_new_n989__,
    new_new_n991__, new_new_n992__, new_new_n993__, new_new_n994__,
    new_new_n995__, new_new_n996__, new_new_n998__, new_new_n999__,
    new_new_n1001__, new_new_n1002__, new_new_n1003__, new_new_n1004__,
    new_new_n1006__, new_new_n1007__, new_new_n1009__, new_new_n1010__,
    new_new_n1011__, new_new_n1012__, new_new_n1013__, new_new_n1014__,
    new_new_n1015__, new_new_n1016__, new_new_n1017__, new_new_n1018__,
    new_new_n1019__, new_new_n1020__, new_new_n1021__, new_new_n1022__,
    new_new_n1023__, new_new_n1024__, new_new_n1025__, new_new_n1026__,
    new_new_n1027__, new_new_n1028__, new_new_n1029__, new_new_n1030__,
    new_new_n1031__, new_new_n1032__, new_new_n1033__, new_new_n1034__,
    new_new_n1035__, new_new_n1036__, new_new_n1037__, new_new_n1038__,
    new_new_n1039__, new_new_n1040__, new_new_n1041__, new_new_n1042__,
    new_new_n1043__, new_new_n1044__, new_new_n1045__, new_new_n1046__,
    new_new_n1047__, new_new_n1048__, new_new_n1049__, new_new_n1050__,
    new_new_n1051__, new_new_n1052__, new_new_n1053__, new_new_n1054__,
    new_new_n1055__, new_new_n1056__, new_new_n1057__, new_new_n1058__,
    new_new_n1059__, new_new_n1060__, new_new_n1061__, new_new_n1062__,
    new_new_n1063__, new_new_n1064__, new_new_n1065__, new_new_n1066__,
    new_new_n1067__, new_new_n1068__, new_new_n1069__, new_new_n1070__,
    new_new_n1071__, new_new_n1072__, new_new_n1073__, new_new_n1074__,
    new_new_n1075__, new_new_n1076__, new_new_n1077__, new_new_n1078__,
    new_new_n1079__, new_new_n1080__, new_new_n1081__, new_new_n1082__,
    new_new_n1083__, new_new_n1084__, new_new_n1085__, new_new_n1086__,
    new_new_n1087__, new_new_n1088__, new_new_n1089__, new_new_n1090__,
    new_new_n1091__, new_new_n1092__, new_new_n1093__, new_new_n1094__,
    new_new_n1095__, new_new_n1096__, new_new_n1097__, new_new_n1098__,
    new_new_n1099__, new_new_n1100__, new_new_n1101__, new_new_n1102__,
    new_new_n1103__, new_new_n1104__, new_new_n1105__, new_new_n1106__,
    new_new_n1107__, new_new_n1108__, new_new_n1109__, new_new_n1110__,
    new_new_n1111__, new_new_n1112__, new_new_n1113__, new_new_n1114__,
    new_new_n1115__, new_new_n1116__, new_new_n1117__, new_new_n1118__,
    new_new_n1119__, new_new_n1120__, new_new_n1121__, new_new_n1123__,
    new_new_n1124__, new_new_n1125__, new_new_n1126__, new_new_n1127__,
    new_new_n1128__, new_new_n1129__, new_new_n1130__, new_new_n1131__,
    new_new_n1132__, new_new_n1133__, new_new_n1134__, new_new_n1135__,
    new_new_n1136__, new_new_n1137__, new_new_n1138__, new_new_n1139__,
    new_new_n1140__, new_new_n1141__, new_new_n1142__, new_new_n1143__,
    new_new_n1144__, new_new_n1145__, new_new_n1146__, new_new_n1147__,
    new_new_n1148__, new_new_n1149__, new_new_n1150__, new_new_n1151__,
    new_new_n1152__, new_new_n1153__, new_new_n1154__, new_new_n1155__,
    new_new_n1156__, new_new_n1157__, new_new_n1158__, new_new_n1159__,
    new_new_n1160__, new_new_n1161__, new_new_n1162__, new_new_n1163__,
    new_new_n1164__, new_new_n1165__, new_new_n1166__, new_new_n1167__,
    new_new_n1168__, new_new_n1169__, new_new_n1170__, new_new_n1171__,
    new_new_n1172__, new_new_n1173__, new_new_n1174__, new_new_n1175__,
    new_new_n1176__, new_new_n1177__, new_new_n1178__, new_new_n1179__,
    new_new_n1180__, new_new_n1181__, new_new_n1182__, new_new_n1183__,
    new_new_n1184__, new_new_n1185__, new_new_n1186__, new_new_n1187__,
    new_new_n1188__, new_new_n1189__, new_new_n1190__, new_new_n1191__,
    new_new_n1192__, new_new_n1193__, new_new_n1194__, new_new_n1195__,
    new_new_n1196__, new_new_n1197__, new_new_n1198__, new_new_n1199__,
    new_new_n1200__, new_new_n1201__, new_new_n1202__, new_new_n1203__,
    new_new_n1204__, new_new_n1205__, new_new_n1206__, new_new_n1207__,
    new_new_n1208__, new_new_n1209__, new_new_n1210__, new_new_n1211__,
    new_new_n1212__, new_new_n1213__, new_new_n1214__, new_new_n1215__,
    new_new_n1216__, new_new_n1217__, new_new_n1218__, new_new_n1219__,
    new_new_n1220__, new_new_n1221__, new_new_n1222__, new_new_n1223__,
    new_new_n1224__, new_new_n1225__, new_new_n1226__, new_new_n1227__,
    new_new_n1228__, new_new_n1229__, new_new_n1230__, new_new_n1231__,
    new_new_n1232__, new_new_n1233__, new_new_n1234__, new_new_n1235__,
    new_new_n1236__, new_new_n1237__, new_new_n1238__, new_new_n1239__,
    new_new_n1240__, new_new_n1241__, new_new_n1242__, new_new_n1243__,
    new_new_n1244__, new_new_n1245__, new_new_n1247__, new_new_n1248__,
    new_new_n1249__, new_new_n1250__, new_new_n1251__, new_new_n1252__,
    new_new_n1253__, new_new_n1254__, new_new_n1255__, new_new_n1256__,
    new_new_n1257__, new_new_n1258__, new_new_n1259__, new_new_n1260__,
    new_new_n1261__, new_new_n1262__, new_new_n1263__, new_new_n1264__,
    new_new_n1265__, new_new_n1266__, new_new_n1267__, new_new_n1268__,
    new_new_n1269__, new_new_n1270__, new_new_n1271__, new_new_n1272__,
    new_new_n1273__, new_new_n1274__, new_new_n1275__, new_new_n1276__,
    new_new_n1277__, new_new_n1278__, new_new_n1279__, new_new_n1280__,
    new_new_n1281__, new_new_n1282__, new_new_n1283__, new_new_n1284__,
    new_new_n1285__, new_new_n1286__, new_new_n1287__, new_new_n1288__,
    new_new_n1289__, new_new_n1290__, new_new_n1291__, new_new_n1292__,
    new_new_n1293__, new_new_n1294__, new_new_n1295__, new_new_n1296__,
    new_new_n1297__, new_new_n1298__, new_new_n1299__, new_new_n1300__,
    new_new_n1301__, new_new_n1302__, new_new_n1303__, new_new_n1304__,
    new_new_n1305__, new_new_n1306__, new_new_n1307__, new_new_n1308__,
    new_new_n1309__, new_new_n1310__, new_new_n1311__, new_new_n1312__,
    new_new_n1313__, new_new_n1314__, new_new_n1315__, new_new_n1316__,
    new_new_n1317__, new_new_n1318__, new_new_n1319__, new_new_n1320__,
    new_new_n1321__, new_new_n1322__, new_new_n1323__, new_new_n1324__,
    new_new_n1325__, new_new_n1326__, new_new_n1327__, new_new_n1328__,
    new_new_n1329__, new_new_n1330__, new_new_n1331__, new_new_n1332__,
    new_new_n1333__, new_new_n1334__, new_new_n1335__, new_new_n1336__,
    new_new_n1337__, new_new_n1338__, new_new_n1339__, new_new_n1340__,
    new_new_n1341__, new_new_n1342__, new_new_n1343__, new_new_n1344__,
    new_new_n1345__, new_new_n1346__, new_new_n1347__, new_new_n1348__,
    new_new_n1349__, new_new_n1350__, new_new_n1351__, new_new_n1352__,
    new_new_n1353__, new_new_n1354__, new_new_n1355__, new_new_n1356__,
    new_new_n1357__, new_new_n1358__, new_new_n1360__, new_new_n1361__,
    new_new_n1363__, new_new_n1364__, new_new_n1366__, new_new_n1367__,
    new_new_n1368__, new_new_n1370__, new_new_n1371__, new_new_n1372__,
    new_new_n1373__, new_new_n1374__, new_new_n1376__, new_new_n1377__,
    new_new_n1378__, new_new_n1379__, new_new_n1380__, new_new_n1382__,
    new_new_n1383__, new_new_n1384__, new_new_n1385__, new_new_n1387__,
    new_new_n1388__, new_new_n1389__, new_new_n1391__, new_new_n1392__,
    new_new_n1393__, new_new_n1394__, new_new_n1395__, new_new_n1396__,
    new_new_n1397__, new_new_n1398__, new_new_n1400__, new_new_n1401__,
    new_new_n1402__, new_new_n1404__, new_new_n1405__, new_new_n1406__,
    new_new_n1407__, new_new_n1408__, new_new_n1410__, new_new_n1412__,
    new_new_n1413__, new_new_n1414__, new_new_n1415__, new_new_n1416__,
    new_new_n1418__, new_new_n1419__, new_new_n1420__, new_new_n1421__,
    new_new_n1422__, new_new_n1423__, new_new_n1424__, new_new_n1426__,
    new_new_n1427__, new_new_n1428__, new_new_n1430__, new_new_n1431__,
    new_new_n1432__, new_new_n1433__, new_new_n1435__, new_new_n1436__,
    new_new_n1438__, new_new_n1439__, new_new_n1441__, new_new_n1442__,
    new_new_n1443__, new_new_n1444__, new_new_n1446__, new_new_n1447__,
    new_new_n1449__, new_new_n1450__, new_new_n1451__, new_new_n1452__,
    new_new_n1453__, new_new_n1454__, new_new_n1455__, new_new_n1456__,
    new_new_n1458__, new_new_n1459__, new_new_n1460__, new_new_n1462__,
    new_new_n1463__, new_new_n1464__, new_new_n1465__, new_new_n1466__,
    new_new_n1468__, new_new_n1470__, new_new_n1471__, new_new_n1472__,
    new_new_n1473__, new_new_n1474__, new_new_n1476__, new_new_n1477__,
    new_new_n1478__, new_new_n1480__, new_new_n1481__, new_new_n1482__,
    new_new_n1483__, new_new_n1485__, new_new_n1486__, new_new_n1488__,
    new_new_n1489__, new_new_n1490__, new_new_n1491__, new_new_n1492__,
    new_new_n1493__, new_new_n1494__, new_new_n1495__, new_new_n1496__,
    new_new_n1497__, new_new_n1498__, new_new_n1499__, new_new_n1500__,
    new_new_n1501__, new_new_n1502__, new_new_n1503__, new_new_n1504__,
    new_new_n1505__, new_new_n1506__, new_new_n1507__, new_new_n1508__,
    new_new_n1509__, new_new_n1510__, new_new_n1511__, new_new_n1512__,
    new_new_n1513__, new_new_n1514__, new_new_n1515__, new_new_n1516__,
    new_new_n1517__, new_new_n1518__, new_new_n1519__, new_new_n1520__,
    new_new_n1521__, new_new_n1522__, new_new_n1523__, new_new_n1524__,
    new_new_n1525__, new_new_n1526__, new_new_n1527__, new_new_n1528__,
    new_new_n1529__, new_new_n1530__, new_new_n1531__, new_new_n1532__,
    new_new_n1533__, new_new_n1534__, new_new_n1535__, new_new_n1536__,
    new_new_n1537__, new_new_n1538__, new_new_n1539__, new_new_n1540__,
    new_new_n1541__, new_new_n1542__, new_new_n1543__, new_new_n1544__,
    new_new_n1545__, new_new_n1546__, new_new_n1547__, new_new_n1548__,
    new_new_n1549__, new_new_n1550__, new_new_n1551__, new_new_n1552__,
    new_new_n1553__, new_new_n1554__, new_new_n1555__, new_new_n1556__,
    new_new_n1557__, new_new_n1558__, new_new_n1559__, new_new_n1560__,
    new_new_n1561__, new_new_n1562__, new_new_n1563__, new_new_n1564__,
    new_new_n1566__, new_new_n1567__, new_new_n1568__, new_new_n1569__,
    new_new_n1570__, new_new_n1571__, new_new_n1572__, new_new_n1573__,
    new_new_n1574__, new_new_n1575__, new_new_n1576__, new_new_n1577__,
    new_new_n1578__, new_new_n1579__, new_new_n1580__, new_new_n1581__,
    new_new_n1582__, new_new_n1583__, new_new_n1584__, new_new_n1585__,
    new_new_n1586__, new_new_n1587__, new_new_n1588__, new_new_n1589__,
    new_new_n1590__, new_new_n1591__, new_new_n1592__, new_new_n1593__,
    new_new_n1594__, new_new_n1595__, new_new_n1596__, new_new_n1597__,
    new_new_n1598__, new_new_n1599__, new_new_n1600__, new_new_n1601__,
    new_new_n1602__, new_new_n1603__, new_new_n1604__, new_new_n1605__,
    new_new_n1606__, new_new_n1607__, new_new_n1608__, new_new_n1609__,
    new_new_n1610__, new_new_n1611__, new_new_n1612__, new_new_n1613__,
    new_new_n1614__, new_new_n1615__, new_new_n1616__, new_new_n1617__,
    new_new_n1618__, new_new_n1619__, new_new_n1620__, new_new_n1621__,
    new_new_n1622__, new_new_n1623__, new_new_n1625__, new_new_n1626__,
    new_new_n1627__, new_new_n1628__, new_new_n1629__, new_new_n1630__,
    new_new_n1631__, new_new_n1632__, new_new_n1633__, new_new_n1634__,
    new_new_n1635__, new_new_n1636__, new_new_n1637__, new_new_n1638__,
    new_new_n1639__, new_new_n1640__, new_new_n1641__, new_new_n1642__,
    new_new_n1643__, new_new_n1644__, new_new_n1645__, new_new_n1646__,
    new_new_n1647__, new_new_n1648__, new_new_n1649__, new_new_n1650__,
    new_new_n1651__, new_new_n1652__, new_new_n1653__, new_new_n1654__,
    new_new_n1655__, new_new_n1656__, new_new_n1657__, new_new_n1658__,
    new_new_n1659__, new_new_n1660__, new_new_n1661__, new_new_n1662__,
    new_new_n1663__, new_new_n1664__, new_new_n1665__, new_new_n1666__,
    new_new_n1667__, new_new_n1668__, new_new_n1669__, new_new_n1670__,
    new_new_n1671__, new_new_n1672__, new_new_n1673__, new_new_n1674__,
    new_new_n1675__, new_new_n1676__, new_new_n1677__, new_new_n1678__,
    new_new_n1679__, new_new_n1680__, new_new_n1681__, new_new_n1682__,
    new_new_n1683__, new_new_n1684__, new_new_n1685__, new_new_n1686__,
    new_new_n1687__, new_new_n1688__, new_new_n1689__, new_new_n1690__,
    new_new_n1691__, new_new_n1692__, new_new_n1693__, new_new_n1694__,
    new_new_n1695__, new_new_n1696__, new_new_n1697__, new_new_n1698__,
    new_new_n1699__, new_new_n1700__, new_new_n1701__, new_new_n1702__,
    new_new_n1704__, new_new_n1705__, new_new_n1706__, new_new_n1707__,
    new_new_n1708__, new_new_n1709__, new_new_n1710__, new_new_n1711__,
    new_new_n1712__, new_new_n1713__, new_new_n1714__, new_new_n1715__,
    new_new_n1716__, new_new_n1717__, new_new_n1718__, new_new_n1719__,
    new_new_n1720__, new_new_n1721__, new_new_n1722__, new_new_n1723__,
    new_new_n1724__, new_new_n1725__, new_new_n1726__, new_new_n1727__,
    new_new_n1728__, new_new_n1729__, new_new_n1730__, new_new_n1731__,
    new_new_n1732__, new_new_n1733__, new_new_n1734__, new_new_n1735__,
    new_new_n1736__, new_new_n1737__, new_new_n1738__, new_new_n1739__,
    new_new_n1740__, new_new_n1741__, new_new_n1742__, new_new_n1743__,
    new_new_n1744__, new_new_n1745__, new_new_n1746__, new_new_n1747__,
    new_new_n1748__, new_new_n1749__, new_new_n1750__, new_new_n1751__,
    new_new_n1752__, new_new_n1753__, new_new_n1754__, new_new_n1755__,
    new_new_n1756__, new_new_n1757__, new_new_n1758__, new_new_n1759__,
    new_new_n1760__, new_new_n1761__, new_new_n1762__, new_new_n1763__,
    new_new_n1764__, new_new_n1765__, new_new_n1766__, new_new_n1767__,
    new_new_n1768__, new_new_n1769__, new_new_n1770__, new_new_n1771__,
    new_new_n1772__, new_new_n1773__, new_new_n1774__, new_new_n1775__,
    new_new_n1776__, new_new_n1777__, new_new_n1778__, new_new_n1779__,
    new_new_n1780__, new_new_n1781__, new_new_n1782__, new_new_n1783__;
  assign G402 = G5 | G57;
  assign new_new_n317__ = G150 & G184;
  assign new_new_n318__ = G228 & G240;
  assign G404 = ~new_new_n317__ | ~new_new_n318__;
  assign new_new_n320__ = G152 & G210;
  assign new_new_n321__ = G218 & G230;
  assign G406 = ~new_new_n320__ | ~new_new_n321__;
  assign new_new_n323__ = G182 & G183;
  assign new_new_n324__ = G185 & G186;
  assign G408 = ~new_new_n323__ | ~new_new_n324__;
  assign new_new_n326__ = G162 & G172;
  assign new_new_n327__ = G188 & G199;
  assign G410 = ~new_new_n326__ | ~new_new_n327__;
  assign G284 = G5 | ~G1197;
  assign new_new_n330__ = ~G5 & G133;
  assign G292 = ~G134 | ~new_new_n330__;
  assign G278 = G1 & G163;
  assign new_new_n333__ = ~G18 & G41;
  assign new_new_n334__ = ~G3701 & new_new_n333__;
  assign new_new_n335__ = G18 & G229;
  assign new_new_n336__ = ~new_new_n333__ & ~new_new_n335__;
  assign new_new_n337__ = ~G18 & G3701;
  assign new_new_n338__ = new_new_n336__ & new_new_n337__;
  assign new_new_n339__ = ~new_new_n334__ & ~new_new_n338__;
  assign new_new_n340__ = G4526 & new_new_n339__;
  assign new_new_n341__ = ~G4526 & ~new_new_n339__;
  assign G373 = ~new_new_n340__ & ~new_new_n341__;
  assign new_new_n343__ = G1496 & G4528;
  assign new_new_n344__ = G1492 & new_new_n343__;
  assign new_new_n345__ = G38 & ~new_new_n344__;
  assign new_new_n346__ = G1492 & G4528;
  assign new_new_n347__ = G38 & ~new_new_n346__;
  assign new_new_n348__ = ~G38 & new_new_n346__;
  assign new_new_n349__ = ~new_new_n347__ & ~new_new_n348__;
  assign new_new_n350__ = G9 & G12;
  assign new_new_n351__ = G18 & ~G157;
  assign new_new_n352__ = ~new_new_n350__ & ~new_new_n351__;
  assign new_new_n353__ = ~G2236 & new_new_n352__;
  assign new_new_n354__ = G2236 & ~new_new_n352__;
  assign new_new_n355__ = ~new_new_n353__ & ~new_new_n354__;
  assign new_new_n356__ = ~G18 & G135;
  assign new_new_n357__ = G18 & G158;
  assign new_new_n358__ = ~new_new_n356__ & ~new_new_n357__;
  assign new_new_n359__ = ~G2230 & ~new_new_n358__;
  assign new_new_n360__ = G2230 & new_new_n358__;
  assign new_new_n361__ = ~new_new_n359__ & ~new_new_n360__;
  assign new_new_n362__ = ~G18 & G144;
  assign new_new_n363__ = G18 & G159;
  assign new_new_n364__ = ~new_new_n362__ & ~new_new_n363__;
  assign new_new_n365__ = ~G2224 & ~new_new_n364__;
  assign new_new_n366__ = G2224 & new_new_n364__;
  assign new_new_n367__ = ~new_new_n365__ & ~new_new_n366__;
  assign new_new_n368__ = ~G18 & G138;
  assign new_new_n369__ = G18 & G160;
  assign new_new_n370__ = ~new_new_n368__ & ~new_new_n369__;
  assign new_new_n371__ = ~G2218 & ~new_new_n370__;
  assign new_new_n372__ = G2218 & new_new_n370__;
  assign new_new_n373__ = ~new_new_n371__ & ~new_new_n372__;
  assign new_new_n374__ = ~G18 & G147;
  assign new_new_n375__ = G18 & G151;
  assign new_new_n376__ = ~new_new_n374__ & ~new_new_n375__;
  assign new_new_n377__ = ~G2211 & ~new_new_n376__;
  assign new_new_n378__ = G2211 & new_new_n376__;
  assign new_new_n379__ = ~new_new_n377__ & ~new_new_n378__;
  assign new_new_n380__ = new_new_n373__ & new_new_n379__;
  assign new_new_n381__ = new_new_n367__ & new_new_n380__;
  assign new_new_n382__ = new_new_n361__ & new_new_n381__;
  assign new_new_n383__ = new_new_n355__ & new_new_n382__;
  assign new_new_n384__ = G18 & ~G154;
  assign new_new_n385__ = ~new_new_n350__ & ~new_new_n384__;
  assign new_new_n386__ = ~G2253 & new_new_n385__;
  assign new_new_n387__ = G2253 & ~new_new_n385__;
  assign new_new_n388__ = ~new_new_n386__ & ~new_new_n387__;
  assign new_new_n389__ = G18 & ~G155;
  assign new_new_n390__ = ~new_new_n350__ & ~new_new_n389__;
  assign new_new_n391__ = ~G2247 & new_new_n390__;
  assign new_new_n392__ = G2247 & ~new_new_n390__;
  assign new_new_n393__ = ~new_new_n391__ & ~new_new_n392__;
  assign new_new_n394__ = G18 & ~G156;
  assign new_new_n395__ = ~new_new_n350__ & ~new_new_n394__;
  assign new_new_n396__ = ~G2239 & new_new_n395__;
  assign new_new_n397__ = G2239 & ~new_new_n395__;
  assign new_new_n398__ = ~new_new_n396__ & ~new_new_n397__;
  assign new_new_n399__ = new_new_n393__ & new_new_n398__;
  assign new_new_n400__ = G18 & ~G153;
  assign new_new_n401__ = ~new_new_n350__ & ~new_new_n400__;
  assign new_new_n402__ = ~G2256 & new_new_n401__;
  assign new_new_n403__ = G2256 & ~new_new_n401__;
  assign new_new_n404__ = ~new_new_n402__ & ~new_new_n403__;
  assign new_new_n405__ = new_new_n388__ & new_new_n404__;
  assign new_new_n406__ = new_new_n399__ & new_new_n405__;
  assign new_new_n407__ = G18 & G235;
  assign new_new_n408__ = ~G18 & G103;
  assign new_new_n409__ = ~new_new_n407__ & ~new_new_n408__;
  assign new_new_n410__ = G3723 & new_new_n409__;
  assign new_new_n411__ = G18 & G236;
  assign new_new_n412__ = ~G18 & G23;
  assign new_new_n413__ = ~new_new_n411__ & ~new_new_n412__;
  assign new_new_n414__ = G3717 & new_new_n413__;
  assign new_new_n415__ = ~G3717 & ~new_new_n413__;
  assign new_new_n416__ = G18 & G237;
  assign new_new_n417__ = ~G18 & G26;
  assign new_new_n418__ = ~new_new_n416__ & ~new_new_n417__;
  assign new_new_n419__ = G3711 & new_new_n418__;
  assign new_new_n420__ = G18 & G238;
  assign new_new_n421__ = ~G18 & G29;
  assign new_new_n422__ = ~new_new_n420__ & ~new_new_n421__;
  assign new_new_n423__ = ~G3705 & ~new_new_n422__;
  assign new_new_n424__ = G3705 & new_new_n422__;
  assign new_new_n425__ = ~new_new_n423__ & ~new_new_n424__;
  assign new_new_n426__ = new_new_n334__ & new_new_n425__;
  assign new_new_n427__ = ~G3711 & ~new_new_n418__;
  assign new_new_n428__ = ~new_new_n423__ & ~new_new_n427__;
  assign new_new_n429__ = ~new_new_n426__ & new_new_n428__;
  assign new_new_n430__ = ~new_new_n419__ & ~new_new_n429__;
  assign new_new_n431__ = ~new_new_n415__ & ~new_new_n430__;
  assign new_new_n432__ = ~new_new_n414__ & ~new_new_n431__;
  assign new_new_n433__ = ~new_new_n410__ & new_new_n432__;
  assign new_new_n434__ = ~G3723 & ~new_new_n409__;
  assign new_new_n435__ = ~new_new_n419__ & ~new_new_n427__;
  assign new_new_n436__ = ~new_new_n414__ & ~new_new_n415__;
  assign new_new_n437__ = new_new_n435__ & new_new_n436__;
  assign new_new_n438__ = new_new_n339__ & new_new_n425__;
  assign new_new_n439__ = G4526 & new_new_n438__;
  assign new_new_n440__ = ~new_new_n410__ & new_new_n437__;
  assign new_new_n441__ = new_new_n439__ & new_new_n440__;
  assign new_new_n442__ = ~new_new_n434__ & ~new_new_n441__;
  assign new_new_n443__ = ~new_new_n433__ & new_new_n442__;
  assign new_new_n444__ = G18 & G233;
  assign new_new_n445__ = ~G18 & G127;
  assign new_new_n446__ = ~new_new_n444__ & ~new_new_n445__;
  assign new_new_n447__ = ~G3737 & ~new_new_n446__;
  assign new_new_n448__ = G3737 & new_new_n446__;
  assign new_new_n449__ = ~new_new_n447__ & ~new_new_n448__;
  assign new_new_n450__ = G18 & G234;
  assign new_new_n451__ = ~G18 & G130;
  assign new_new_n452__ = ~new_new_n450__ & ~new_new_n451__;
  assign new_new_n453__ = ~G3729 & ~new_new_n452__;
  assign new_new_n454__ = G3729 & new_new_n452__;
  assign new_new_n455__ = ~new_new_n453__ & ~new_new_n454__;
  assign new_new_n456__ = new_new_n449__ & new_new_n455__;
  assign new_new_n457__ = G18 & G232;
  assign new_new_n458__ = ~G18 & G124;
  assign new_new_n459__ = ~new_new_n457__ & ~new_new_n458__;
  assign new_new_n460__ = ~G3743 & ~new_new_n459__;
  assign new_new_n461__ = G3743 & new_new_n459__;
  assign new_new_n462__ = ~new_new_n460__ & ~new_new_n461__;
  assign new_new_n463__ = G18 & G231;
  assign new_new_n464__ = ~G18 & G100;
  assign new_new_n465__ = ~new_new_n463__ & ~new_new_n464__;
  assign new_new_n466__ = G3749 & new_new_n465__;
  assign new_new_n467__ = ~G3749 & ~new_new_n465__;
  assign new_new_n468__ = ~new_new_n466__ & ~new_new_n467__;
  assign new_new_n469__ = new_new_n462__ & new_new_n468__;
  assign new_new_n470__ = new_new_n456__ & new_new_n469__;
  assign new_new_n471__ = ~new_new_n443__ & new_new_n470__;
  assign new_new_n472__ = new_new_n449__ & new_new_n453__;
  assign new_new_n473__ = ~new_new_n447__ & ~new_new_n472__;
  assign new_new_n474__ = new_new_n469__ & ~new_new_n473__;
  assign new_new_n475__ = new_new_n460__ & ~new_new_n466__;
  assign new_new_n476__ = ~new_new_n467__ & ~new_new_n475__;
  assign new_new_n477__ = ~new_new_n474__ & new_new_n476__;
  assign new_new_n478__ = ~new_new_n471__ & new_new_n477__;
  assign new_new_n479__ = G18 & G223;
  assign new_new_n480__ = ~G18 & G47;
  assign new_new_n481__ = ~new_new_n479__ & ~new_new_n480__;
  assign new_new_n482__ = G4415 & new_new_n481__;
  assign new_new_n483__ = ~G4415 & ~new_new_n481__;
  assign new_new_n484__ = ~new_new_n482__ & ~new_new_n483__;
  assign new_new_n485__ = G18 & G224;
  assign new_new_n486__ = ~G18 & G121;
  assign new_new_n487__ = ~new_new_n485__ & ~new_new_n486__;
  assign new_new_n488__ = ~G4410 & ~new_new_n487__;
  assign new_new_n489__ = G4410 & new_new_n487__;
  assign new_new_n490__ = ~new_new_n488__ & ~new_new_n489__;
  assign new_new_n491__ = G18 & G226;
  assign new_new_n492__ = ~G18 & G97;
  assign new_new_n493__ = ~new_new_n491__ & ~new_new_n492__;
  assign new_new_n494__ = G4400 & new_new_n493__;
  assign new_new_n495__ = G18 & G217;
  assign new_new_n496__ = ~G18 & G118;
  assign new_new_n497__ = ~new_new_n495__ & ~new_new_n496__;
  assign new_new_n498__ = ~G4394 & ~new_new_n497__;
  assign new_new_n499__ = G4394 & new_new_n497__;
  assign new_new_n500__ = ~new_new_n498__ & ~new_new_n499__;
  assign new_new_n501__ = ~new_new_n494__ & new_new_n500__;
  assign new_new_n502__ = G18 & G225;
  assign new_new_n503__ = ~G18 & G94;
  assign new_new_n504__ = ~new_new_n502__ & ~new_new_n503__;
  assign new_new_n505__ = ~G4405 & ~new_new_n504__;
  assign new_new_n506__ = G4405 & new_new_n504__;
  assign new_new_n507__ = ~new_new_n505__ & ~new_new_n506__;
  assign new_new_n508__ = ~G4400 & ~new_new_n493__;
  assign new_new_n509__ = new_new_n507__ & ~new_new_n508__;
  assign new_new_n510__ = new_new_n501__ & new_new_n509__;
  assign new_new_n511__ = new_new_n484__ & new_new_n490__;
  assign new_new_n512__ = new_new_n510__ & new_new_n511__;
  assign new_new_n513__ = ~new_new_n478__ & new_new_n512__;
  assign new_new_n514__ = ~new_new_n482__ & new_new_n488__;
  assign new_new_n515__ = ~new_new_n494__ & ~new_new_n508__;
  assign new_new_n516__ = new_new_n498__ & new_new_n515__;
  assign new_new_n517__ = new_new_n507__ & new_new_n516__;
  assign new_new_n518__ = ~new_new_n505__ & ~new_new_n517__;
  assign new_new_n519__ = new_new_n511__ & ~new_new_n518__;
  assign new_new_n520__ = new_new_n507__ & new_new_n508__;
  assign new_new_n521__ = new_new_n511__ & new_new_n520__;
  assign new_new_n522__ = ~new_new_n483__ & ~new_new_n514__;
  assign new_new_n523__ = ~new_new_n521__ & new_new_n522__;
  assign new_new_n524__ = ~new_new_n519__ & new_new_n523__;
  assign new_new_n525__ = ~new_new_n513__ & new_new_n524__;
  assign new_new_n526__ = G18 & G221;
  assign new_new_n527__ = ~G18 & G32;
  assign new_new_n528__ = ~new_new_n526__ & ~new_new_n527__;
  assign new_new_n529__ = ~G4427 & ~new_new_n528__;
  assign new_new_n530__ = G4427 & new_new_n528__;
  assign new_new_n531__ = ~new_new_n529__ & ~new_new_n530__;
  assign new_new_n532__ = G18 & G222;
  assign new_new_n533__ = ~G18 & G35;
  assign new_new_n534__ = ~new_new_n532__ & ~new_new_n533__;
  assign new_new_n535__ = ~G4420 & ~new_new_n534__;
  assign new_new_n536__ = G4420 & new_new_n534__;
  assign new_new_n537__ = ~new_new_n535__ & ~new_new_n536__;
  assign new_new_n538__ = new_new_n531__ & new_new_n537__;
  assign new_new_n539__ = G18 & G219;
  assign new_new_n540__ = ~G18 & G66;
  assign new_new_n541__ = ~new_new_n539__ & ~new_new_n540__;
  assign new_new_n542__ = ~G4437 & ~new_new_n541__;
  assign new_new_n543__ = G4437 & new_new_n541__;
  assign new_new_n544__ = ~new_new_n542__ & ~new_new_n543__;
  assign new_new_n545__ = G18 & G220;
  assign new_new_n546__ = ~G18 & G50;
  assign new_new_n547__ = ~new_new_n545__ & ~new_new_n546__;
  assign new_new_n548__ = G4432 & new_new_n547__;
  assign new_new_n549__ = ~G4432 & ~new_new_n547__;
  assign new_new_n550__ = ~new_new_n548__ & ~new_new_n549__;
  assign new_new_n551__ = new_new_n544__ & new_new_n550__;
  assign new_new_n552__ = new_new_n538__ & new_new_n551__;
  assign new_new_n553__ = ~new_new_n525__ & new_new_n552__;
  assign new_new_n554__ = new_new_n531__ & new_new_n535__;
  assign new_new_n555__ = ~new_new_n529__ & ~new_new_n554__;
  assign new_new_n556__ = ~new_new_n548__ & ~new_new_n555__;
  assign new_new_n557__ = ~new_new_n549__ & ~new_new_n556__;
  assign new_new_n558__ = ~new_new_n542__ & new_new_n557__;
  assign new_new_n559__ = ~new_new_n543__ & ~new_new_n558__;
  assign new_new_n560__ = ~new_new_n553__ & ~new_new_n559__;
  assign new_new_n561__ = new_new_n383__ & new_new_n406__;
  assign new_new_n562__ = ~new_new_n560__ & new_new_n561__;
  assign new_new_n563__ = new_new_n393__ & new_new_n396__;
  assign new_new_n564__ = ~new_new_n391__ & ~new_new_n563__;
  assign new_new_n565__ = ~new_new_n386__ & new_new_n564__;
  assign new_new_n566__ = ~new_new_n387__ & ~new_new_n565__;
  assign new_new_n567__ = ~new_new_n403__ & new_new_n566__;
  assign new_new_n568__ = new_new_n373__ & new_new_n377__;
  assign new_new_n569__ = ~new_new_n365__ & ~new_new_n371__;
  assign new_new_n570__ = ~new_new_n568__ & new_new_n569__;
  assign new_new_n571__ = ~new_new_n366__ & ~new_new_n570__;
  assign new_new_n572__ = ~new_new_n360__ & new_new_n571__;
  assign new_new_n573__ = ~new_new_n359__ & ~new_new_n572__;
  assign new_new_n574__ = ~new_new_n354__ & ~new_new_n573__;
  assign new_new_n575__ = ~new_new_n353__ & ~new_new_n574__;
  assign new_new_n576__ = new_new_n406__ & ~new_new_n575__;
  assign new_new_n577__ = ~new_new_n402__ & ~new_new_n567__;
  assign new_new_n578__ = ~new_new_n576__ & new_new_n577__;
  assign new_new_n579__ = ~new_new_n562__ & new_new_n578__;
  assign new_new_n580__ = G18 & ~G213;
  assign new_new_n581__ = ~new_new_n350__ & ~new_new_n580__;
  assign new_new_n582__ = G1486 & ~new_new_n581__;
  assign new_new_n583__ = ~G1486 & new_new_n581__;
  assign new_new_n584__ = ~new_new_n582__ & ~new_new_n583__;
  assign new_new_n585__ = G18 & ~G214;
  assign new_new_n586__ = ~new_new_n350__ & ~new_new_n585__;
  assign new_new_n587__ = ~G1480 & new_new_n586__;
  assign new_new_n588__ = G1480 & ~new_new_n586__;
  assign new_new_n589__ = ~new_new_n587__ & ~new_new_n588__;
  assign new_new_n590__ = G18 & ~G216;
  assign new_new_n591__ = ~new_new_n350__ & ~new_new_n590__;
  assign new_new_n592__ = G1469 & ~new_new_n591__;
  assign new_new_n593__ = G18 & ~G209;
  assign new_new_n594__ = ~new_new_n350__ & ~new_new_n593__;
  assign new_new_n595__ = ~G1462 & new_new_n594__;
  assign new_new_n596__ = G1462 & ~new_new_n594__;
  assign new_new_n597__ = ~new_new_n595__ & ~new_new_n596__;
  assign new_new_n598__ = ~new_new_n592__ & new_new_n597__;
  assign new_new_n599__ = G18 & ~G215;
  assign new_new_n600__ = ~new_new_n350__ & ~new_new_n599__;
  assign new_new_n601__ = ~G106 & new_new_n600__;
  assign new_new_n602__ = G106 & ~new_new_n600__;
  assign new_new_n603__ = ~new_new_n601__ & ~new_new_n602__;
  assign new_new_n604__ = ~G1469 & new_new_n591__;
  assign new_new_n605__ = new_new_n603__ & ~new_new_n604__;
  assign new_new_n606__ = new_new_n598__ & new_new_n605__;
  assign new_new_n607__ = new_new_n584__ & new_new_n589__;
  assign new_new_n608__ = new_new_n606__ & new_new_n607__;
  assign new_new_n609__ = ~new_new_n579__ & new_new_n608__;
  assign new_new_n610__ = ~new_new_n582__ & new_new_n587__;
  assign new_new_n611__ = ~new_new_n592__ & ~new_new_n604__;
  assign new_new_n612__ = new_new_n595__ & new_new_n611__;
  assign new_new_n613__ = new_new_n603__ & new_new_n612__;
  assign new_new_n614__ = ~new_new_n601__ & ~new_new_n613__;
  assign new_new_n615__ = new_new_n607__ & ~new_new_n614__;
  assign new_new_n616__ = new_new_n603__ & new_new_n604__;
  assign new_new_n617__ = new_new_n607__ & new_new_n616__;
  assign new_new_n618__ = ~new_new_n583__ & ~new_new_n610__;
  assign new_new_n619__ = ~new_new_n617__ & new_new_n618__;
  assign new_new_n620__ = ~new_new_n615__ & new_new_n619__;
  assign new_new_n621__ = ~new_new_n609__ & new_new_n620__;
  assign new_new_n622__ = G38 & new_new_n343__;
  assign new_new_n623__ = ~G38 & ~new_new_n343__;
  assign new_new_n624__ = ~new_new_n622__ & ~new_new_n623__;
  assign new_new_n625__ = new_new_n349__ & ~new_new_n624__;
  assign new_new_n626__ = ~new_new_n621__ & new_new_n625__;
  assign G246 = new_new_n345__ | new_new_n626__;
  assign new_new_n628__ = G18 & G1462;
  assign new_new_n629__ = ~G18 & ~G113;
  assign new_new_n630__ = ~new_new_n628__ & ~new_new_n629__;
  assign new_new_n631__ = ~new_new_n350__ & new_new_n630__;
  assign new_new_n632__ = G18 & ~G169;
  assign new_new_n633__ = ~new_new_n350__ & ~new_new_n632__;
  assign new_new_n634__ = G18 & G1469;
  assign new_new_n635__ = ~G18 & ~G111;
  assign new_new_n636__ = ~new_new_n634__ & ~new_new_n635__;
  assign new_new_n637__ = ~new_new_n633__ & ~new_new_n636__;
  assign new_new_n638__ = new_new_n633__ & new_new_n636__;
  assign new_new_n639__ = G18 & ~G167;
  assign new_new_n640__ = ~new_new_n350__ & ~new_new_n639__;
  assign new_new_n641__ = G18 & G1480;
  assign new_new_n642__ = ~G18 & ~G112;
  assign new_new_n643__ = ~new_new_n641__ & ~new_new_n642__;
  assign new_new_n644__ = new_new_n640__ & new_new_n643__;
  assign new_new_n645__ = G18 & ~G168;
  assign new_new_n646__ = ~new_new_n350__ & ~new_new_n645__;
  assign new_new_n647__ = G18 & G106;
  assign new_new_n648__ = ~G18 & ~G87;
  assign new_new_n649__ = ~new_new_n647__ & ~new_new_n648__;
  assign new_new_n650__ = new_new_n646__ & new_new_n649__;
  assign new_new_n651__ = ~new_new_n644__ & ~new_new_n650__;
  assign new_new_n652__ = ~new_new_n640__ & ~new_new_n643__;
  assign new_new_n653__ = ~new_new_n646__ & ~new_new_n649__;
  assign new_new_n654__ = ~new_new_n637__ & ~new_new_n638__;
  assign new_new_n655__ = ~new_new_n652__ & ~new_new_n653__;
  assign new_new_n656__ = new_new_n654__ & new_new_n655__;
  assign new_new_n657__ = new_new_n651__ & new_new_n656__;
  assign new_new_n658__ = G18 & ~G166;
  assign new_new_n659__ = ~new_new_n350__ & ~new_new_n658__;
  assign new_new_n660__ = G18 & G1486;
  assign new_new_n661__ = ~G18 & ~G88;
  assign new_new_n662__ = ~new_new_n660__ & ~new_new_n661__;
  assign new_new_n663__ = ~new_new_n659__ & ~new_new_n662__;
  assign new_new_n664__ = new_new_n659__ & new_new_n662__;
  assign new_new_n665__ = new_new_n350__ & ~new_new_n630__;
  assign new_new_n666__ = G18 & ~G174;
  assign new_new_n667__ = ~new_new_n350__ & ~new_new_n666__;
  assign new_new_n668__ = G18 & G2253;
  assign new_new_n669__ = ~G18 & ~G109;
  assign new_new_n670__ = ~new_new_n668__ & ~new_new_n669__;
  assign new_new_n671__ = new_new_n667__ & new_new_n670__;
  assign new_new_n672__ = G18 & ~G175;
  assign new_new_n673__ = ~new_new_n350__ & ~new_new_n672__;
  assign new_new_n674__ = G18 & G2247;
  assign new_new_n675__ = ~G18 & ~G86;
  assign new_new_n676__ = ~new_new_n674__ & ~new_new_n675__;
  assign new_new_n677__ = new_new_n673__ & new_new_n676__;
  assign new_new_n678__ = ~new_new_n671__ & ~new_new_n677__;
  assign new_new_n679__ = ~new_new_n667__ & ~new_new_n670__;
  assign new_new_n680__ = ~new_new_n673__ & ~new_new_n676__;
  assign new_new_n681__ = ~new_new_n679__ & ~new_new_n680__;
  assign new_new_n682__ = new_new_n678__ & new_new_n681__;
  assign new_new_n683__ = G18 & ~G173;
  assign new_new_n684__ = ~new_new_n350__ & ~new_new_n683__;
  assign new_new_n685__ = G18 & G2256;
  assign new_new_n686__ = ~G18 & ~G110;
  assign new_new_n687__ = ~new_new_n685__ & ~new_new_n686__;
  assign new_new_n688__ = ~new_new_n684__ & ~new_new_n687__;
  assign new_new_n689__ = new_new_n684__ & new_new_n687__;
  assign new_new_n690__ = ~new_new_n688__ & ~new_new_n689__;
  assign new_new_n691__ = G18 & ~G176;
  assign new_new_n692__ = ~new_new_n350__ & ~new_new_n691__;
  assign new_new_n693__ = G18 & G2239;
  assign new_new_n694__ = ~G18 & ~G63;
  assign new_new_n695__ = ~new_new_n693__ & ~new_new_n694__;
  assign new_new_n696__ = new_new_n692__ & new_new_n695__;
  assign new_new_n697__ = new_new_n690__ & new_new_n696__;
  assign new_new_n698__ = ~new_new_n692__ & ~new_new_n695__;
  assign new_new_n699__ = ~new_new_n696__ & ~new_new_n698__;
  assign new_new_n700__ = new_new_n690__ & new_new_n699__;
  assign new_new_n701__ = G18 & ~G177;
  assign new_new_n702__ = ~new_new_n350__ & ~new_new_n701__;
  assign new_new_n703__ = G18 & G2236;
  assign new_new_n704__ = ~G18 & ~G64;
  assign new_new_n705__ = ~new_new_n703__ & ~new_new_n704__;
  assign new_new_n706__ = ~new_new_n702__ & ~new_new_n705__;
  assign new_new_n707__ = G18 & G178;
  assign new_new_n708__ = ~new_new_n356__ & ~new_new_n707__;
  assign new_new_n709__ = G18 & G2230;
  assign new_new_n710__ = ~G18 & ~G85;
  assign new_new_n711__ = ~new_new_n709__ & ~new_new_n710__;
  assign new_new_n712__ = ~new_new_n708__ & new_new_n711__;
  assign new_new_n713__ = new_new_n702__ & new_new_n705__;
  assign new_new_n714__ = G18 & G179;
  assign new_new_n715__ = ~new_new_n362__ & ~new_new_n714__;
  assign new_new_n716__ = G18 & G2224;
  assign new_new_n717__ = ~G18 & ~G84;
  assign new_new_n718__ = ~new_new_n716__ & ~new_new_n717__;
  assign new_new_n719__ = new_new_n715__ & ~new_new_n718__;
  assign new_new_n720__ = new_new_n708__ & ~new_new_n711__;
  assign new_new_n721__ = ~new_new_n715__ & new_new_n718__;
  assign new_new_n722__ = G18 & G180;
  assign new_new_n723__ = ~new_new_n368__ & ~new_new_n722__;
  assign new_new_n724__ = G18 & G2218;
  assign new_new_n725__ = ~G18 & ~G83;
  assign new_new_n726__ = ~new_new_n724__ & ~new_new_n725__;
  assign new_new_n727__ = ~new_new_n723__ & new_new_n726__;
  assign new_new_n728__ = new_new_n723__ & ~new_new_n726__;
  assign new_new_n729__ = G18 & G171;
  assign new_new_n730__ = ~new_new_n374__ & ~new_new_n729__;
  assign new_new_n731__ = G18 & G2211;
  assign new_new_n732__ = ~G18 & ~G65;
  assign new_new_n733__ = ~new_new_n731__ & ~new_new_n732__;
  assign new_new_n734__ = ~new_new_n730__ & new_new_n733__;
  assign new_new_n735__ = ~new_new_n728__ & new_new_n734__;
  assign new_new_n736__ = ~new_new_n721__ & ~new_new_n727__;
  assign new_new_n737__ = ~new_new_n735__ & new_new_n736__;
  assign new_new_n738__ = ~new_new_n719__ & ~new_new_n720__;
  assign new_new_n739__ = ~new_new_n737__ & new_new_n738__;
  assign new_new_n740__ = ~new_new_n712__ & ~new_new_n713__;
  assign new_new_n741__ = ~new_new_n739__ & new_new_n740__;
  assign new_new_n742__ = new_new_n700__ & ~new_new_n706__;
  assign new_new_n743__ = ~new_new_n741__ & new_new_n742__;
  assign new_new_n744__ = ~new_new_n697__ & ~new_new_n743__;
  assign new_new_n745__ = new_new_n682__ & ~new_new_n744__;
  assign new_new_n746__ = new_new_n730__ & ~new_new_n733__;
  assign new_new_n747__ = G18 & G189;
  assign new_new_n748__ = ~new_new_n540__ & ~new_new_n747__;
  assign new_new_n749__ = ~G18 & ~G62;
  assign new_new_n750__ = G18 & G4437;
  assign new_new_n751__ = ~new_new_n749__ & ~new_new_n750__;
  assign new_new_n752__ = ~new_new_n748__ & new_new_n751__;
  assign new_new_n753__ = new_new_n748__ & ~new_new_n751__;
  assign new_new_n754__ = ~new_new_n752__ & ~new_new_n753__;
  assign new_new_n755__ = G18 & G192;
  assign new_new_n756__ = ~new_new_n533__ & ~new_new_n755__;
  assign new_new_n757__ = ~G18 & ~G79;
  assign new_new_n758__ = G18 & G4420;
  assign new_new_n759__ = ~new_new_n757__ & ~new_new_n758__;
  assign new_new_n760__ = ~new_new_n756__ & new_new_n759__;
  assign new_new_n761__ = new_new_n756__ & ~new_new_n759__;
  assign new_new_n762__ = G18 & G190;
  assign new_new_n763__ = ~new_new_n546__ & ~new_new_n762__;
  assign new_new_n764__ = ~G18 & ~G61;
  assign new_new_n765__ = G18 & G4432;
  assign new_new_n766__ = ~new_new_n764__ & ~new_new_n765__;
  assign new_new_n767__ = ~new_new_n763__ & new_new_n766__;
  assign new_new_n768__ = G18 & G191;
  assign new_new_n769__ = ~new_new_n527__ & ~new_new_n768__;
  assign new_new_n770__ = ~G18 & ~G60;
  assign new_new_n771__ = G18 & G4427;
  assign new_new_n772__ = ~new_new_n770__ & ~new_new_n771__;
  assign new_new_n773__ = ~new_new_n769__ & new_new_n772__;
  assign new_new_n774__ = ~new_new_n767__ & ~new_new_n773__;
  assign new_new_n775__ = new_new_n763__ & ~new_new_n766__;
  assign new_new_n776__ = new_new_n769__ & ~new_new_n772__;
  assign new_new_n777__ = ~new_new_n775__ & ~new_new_n776__;
  assign new_new_n778__ = new_new_n774__ & new_new_n777__;
  assign new_new_n779__ = ~new_new_n760__ & ~new_new_n761__;
  assign new_new_n780__ = new_new_n754__ & new_new_n779__;
  assign new_new_n781__ = new_new_n778__ & new_new_n780__;
  assign new_new_n782__ = G18 & G193;
  assign new_new_n783__ = ~new_new_n480__ & ~new_new_n782__;
  assign new_new_n784__ = ~G18 & ~G80;
  assign new_new_n785__ = G18 & G4415;
  assign new_new_n786__ = ~new_new_n784__ & ~new_new_n785__;
  assign new_new_n787__ = new_new_n783__ & ~new_new_n786__;
  assign new_new_n788__ = G18 & G187;
  assign new_new_n789__ = ~new_new_n496__ & ~new_new_n788__;
  assign new_new_n790__ = ~G18 & ~G77;
  assign new_new_n791__ = G18 & G4394;
  assign new_new_n792__ = ~new_new_n790__ & ~new_new_n791__;
  assign new_new_n793__ = ~new_new_n789__ & new_new_n792__;
  assign new_new_n794__ = G18 & G196;
  assign new_new_n795__ = ~new_new_n492__ & ~new_new_n794__;
  assign new_new_n796__ = ~G18 & ~G78;
  assign new_new_n797__ = G18 & G4400;
  assign new_new_n798__ = ~new_new_n796__ & ~new_new_n797__;
  assign new_new_n799__ = ~new_new_n795__ & new_new_n798__;
  assign new_new_n800__ = ~new_new_n793__ & ~new_new_n799__;
  assign new_new_n801__ = G18 & G194;
  assign new_new_n802__ = ~new_new_n486__ & ~new_new_n801__;
  assign new_new_n803__ = ~G18 & ~G81;
  assign new_new_n804__ = G18 & G4410;
  assign new_new_n805__ = ~new_new_n803__ & ~new_new_n804__;
  assign new_new_n806__ = new_new_n802__ & ~new_new_n805__;
  assign new_new_n807__ = ~new_new_n802__ & new_new_n805__;
  assign new_new_n808__ = G18 & G195;
  assign new_new_n809__ = ~new_new_n503__ & ~new_new_n808__;
  assign new_new_n810__ = ~G18 & ~G59;
  assign new_new_n811__ = G18 & G4405;
  assign new_new_n812__ = ~new_new_n810__ & ~new_new_n811__;
  assign new_new_n813__ = ~new_new_n809__ & new_new_n812__;
  assign new_new_n814__ = ~new_new_n783__ & new_new_n786__;
  assign new_new_n815__ = new_new_n795__ & ~new_new_n798__;
  assign new_new_n816__ = new_new_n809__ & ~new_new_n812__;
  assign new_new_n817__ = new_new_n789__ & ~new_new_n792__;
  assign new_new_n818__ = ~new_new_n787__ & ~new_new_n806__;
  assign new_new_n819__ = ~new_new_n807__ & ~new_new_n813__;
  assign new_new_n820__ = ~new_new_n814__ & ~new_new_n815__;
  assign new_new_n821__ = ~new_new_n816__ & ~new_new_n817__;
  assign new_new_n822__ = new_new_n820__ & new_new_n821__;
  assign new_new_n823__ = new_new_n818__ & new_new_n819__;
  assign new_new_n824__ = new_new_n800__ & new_new_n823__;
  assign new_new_n825__ = new_new_n822__ & new_new_n824__;
  assign new_new_n826__ = G18 & G200;
  assign new_new_n827__ = ~new_new_n464__ & ~new_new_n826__;
  assign new_new_n828__ = ~G18 & ~G56;
  assign new_new_n829__ = G18 & G3749;
  assign new_new_n830__ = ~new_new_n828__ & ~new_new_n829__;
  assign new_new_n831__ = new_new_n827__ & ~new_new_n830__;
  assign new_new_n832__ = ~new_new_n827__ & new_new_n830__;
  assign new_new_n833__ = G18 & G201;
  assign new_new_n834__ = ~new_new_n458__ & ~new_new_n833__;
  assign new_new_n835__ = ~G18 & ~G55;
  assign new_new_n836__ = G18 & G3743;
  assign new_new_n837__ = ~new_new_n835__ & ~new_new_n836__;
  assign new_new_n838__ = ~new_new_n834__ & new_new_n837__;
  assign new_new_n839__ = ~new_new_n832__ & ~new_new_n838__;
  assign new_new_n840__ = ~new_new_n831__ & ~new_new_n839__;
  assign new_new_n841__ = new_new_n834__ & ~new_new_n837__;
  assign new_new_n842__ = ~new_new_n831__ & ~new_new_n841__;
  assign new_new_n843__ = new_new_n839__ & new_new_n842__;
  assign new_new_n844__ = G18 & G202;
  assign new_new_n845__ = ~new_new_n445__ & ~new_new_n844__;
  assign new_new_n846__ = ~G18 & ~G54;
  assign new_new_n847__ = G18 & G3737;
  assign new_new_n848__ = ~new_new_n846__ & ~new_new_n847__;
  assign new_new_n849__ = new_new_n845__ & ~new_new_n848__;
  assign new_new_n850__ = ~new_new_n845__ & new_new_n848__;
  assign new_new_n851__ = G18 & G203;
  assign new_new_n852__ = ~new_new_n451__ & ~new_new_n851__;
  assign new_new_n853__ = ~G18 & ~G53;
  assign new_new_n854__ = G18 & G3729;
  assign new_new_n855__ = ~new_new_n853__ & ~new_new_n854__;
  assign new_new_n856__ = ~new_new_n852__ & new_new_n855__;
  assign new_new_n857__ = ~new_new_n850__ & ~new_new_n856__;
  assign new_new_n858__ = ~new_new_n849__ & ~new_new_n857__;
  assign new_new_n859__ = new_new_n843__ & new_new_n858__;
  assign new_new_n860__ = G18 & G205;
  assign new_new_n861__ = ~new_new_n412__ & ~new_new_n860__;
  assign new_new_n862__ = ~G18 & ~G75;
  assign new_new_n863__ = G18 & G3717;
  assign new_new_n864__ = ~new_new_n862__ & ~new_new_n863__;
  assign new_new_n865__ = ~new_new_n861__ & new_new_n864__;
  assign new_new_n866__ = G18 & G206;
  assign new_new_n867__ = ~new_new_n417__ & ~new_new_n866__;
  assign new_new_n868__ = ~G18 & ~G76;
  assign new_new_n869__ = G18 & G3711;
  assign new_new_n870__ = ~new_new_n868__ & ~new_new_n869__;
  assign new_new_n871__ = new_new_n867__ & ~new_new_n870__;
  assign new_new_n872__ = G18 & G207;
  assign new_new_n873__ = ~new_new_n421__ & ~new_new_n872__;
  assign new_new_n874__ = ~G18 & ~G74;
  assign new_new_n875__ = G18 & G3705;
  assign new_new_n876__ = ~new_new_n874__ & ~new_new_n875__;
  assign new_new_n877__ = ~new_new_n873__ & new_new_n876__;
  assign new_new_n878__ = ~new_new_n867__ & new_new_n870__;
  assign new_new_n879__ = new_new_n873__ & ~new_new_n876__;
  assign new_new_n880__ = ~G18 & ~G70;
  assign new_new_n881__ = new_new_n333__ & ~new_new_n880__;
  assign new_new_n882__ = ~new_new_n879__ & new_new_n881__;
  assign new_new_n883__ = ~new_new_n877__ & ~new_new_n878__;
  assign new_new_n884__ = ~new_new_n882__ & new_new_n883__;
  assign new_new_n885__ = ~new_new_n871__ & ~new_new_n884__;
  assign new_new_n886__ = ~new_new_n865__ & ~new_new_n885__;
  assign new_new_n887__ = G18 & G204;
  assign new_new_n888__ = ~new_new_n408__ & ~new_new_n887__;
  assign new_new_n889__ = ~G18 & ~G73;
  assign new_new_n890__ = G18 & G3723;
  assign new_new_n891__ = ~new_new_n889__ & ~new_new_n890__;
  assign new_new_n892__ = new_new_n888__ & ~new_new_n891__;
  assign new_new_n893__ = new_new_n861__ & ~new_new_n864__;
  assign new_new_n894__ = ~new_new_n892__ & ~new_new_n893__;
  assign new_new_n895__ = ~new_new_n886__ & new_new_n894__;
  assign new_new_n896__ = ~new_new_n888__ & new_new_n891__;
  assign new_new_n897__ = ~new_new_n333__ & new_new_n880__;
  assign new_new_n898__ = G89 & ~new_new_n881__;
  assign new_new_n899__ = ~new_new_n897__ & new_new_n898__;
  assign new_new_n900__ = ~new_new_n865__ & ~new_new_n871__;
  assign new_new_n901__ = ~new_new_n879__ & ~new_new_n892__;
  assign new_new_n902__ = ~new_new_n893__ & ~new_new_n896__;
  assign new_new_n903__ = new_new_n901__ & new_new_n902__;
  assign new_new_n904__ = new_new_n883__ & new_new_n900__;
  assign new_new_n905__ = new_new_n899__ & new_new_n904__;
  assign new_new_n906__ = new_new_n903__ & new_new_n905__;
  assign new_new_n907__ = ~new_new_n896__ & ~new_new_n906__;
  assign new_new_n908__ = ~new_new_n895__ & new_new_n907__;
  assign new_new_n909__ = new_new_n852__ & ~new_new_n855__;
  assign new_new_n910__ = ~new_new_n849__ & ~new_new_n909__;
  assign new_new_n911__ = new_new_n857__ & new_new_n910__;
  assign new_new_n912__ = new_new_n843__ & new_new_n911__;
  assign new_new_n913__ = ~new_new_n908__ & new_new_n912__;
  assign new_new_n914__ = ~new_new_n840__ & ~new_new_n859__;
  assign new_new_n915__ = ~new_new_n913__ & new_new_n914__;
  assign new_new_n916__ = new_new_n781__ & new_new_n825__;
  assign new_new_n917__ = ~new_new_n915__ & new_new_n916__;
  assign new_new_n918__ = ~new_new_n800__ & ~new_new_n815__;
  assign new_new_n919__ = ~new_new_n813__ & ~new_new_n918__;
  assign new_new_n920__ = ~new_new_n816__ & ~new_new_n919__;
  assign new_new_n921__ = ~new_new_n807__ & ~new_new_n920__;
  assign new_new_n922__ = new_new_n818__ & ~new_new_n921__;
  assign new_new_n923__ = ~new_new_n814__ & ~new_new_n922__;
  assign new_new_n924__ = new_new_n781__ & ~new_new_n923__;
  assign new_new_n925__ = ~new_new_n753__ & ~new_new_n775__;
  assign new_new_n926__ = ~new_new_n774__ & new_new_n925__;
  assign new_new_n927__ = new_new_n754__ & new_new_n760__;
  assign new_new_n928__ = new_new_n778__ & new_new_n927__;
  assign new_new_n929__ = ~new_new_n752__ & ~new_new_n926__;
  assign new_new_n930__ = ~new_new_n928__ & new_new_n929__;
  assign new_new_n931__ = ~new_new_n924__ & new_new_n930__;
  assign new_new_n932__ = ~new_new_n917__ & new_new_n931__;
  assign new_new_n933__ = ~new_new_n706__ & ~new_new_n712__;
  assign new_new_n934__ = ~new_new_n713__ & ~new_new_n719__;
  assign new_new_n935__ = ~new_new_n720__ & ~new_new_n721__;
  assign new_new_n936__ = ~new_new_n727__ & ~new_new_n728__;
  assign new_new_n937__ = ~new_new_n734__ & ~new_new_n746__;
  assign new_new_n938__ = new_new_n936__ & new_new_n937__;
  assign new_new_n939__ = new_new_n934__ & new_new_n935__;
  assign new_new_n940__ = new_new_n933__ & new_new_n939__;
  assign new_new_n941__ = new_new_n682__ & new_new_n938__;
  assign new_new_n942__ = new_new_n700__ & new_new_n941__;
  assign new_new_n943__ = new_new_n940__ & new_new_n942__;
  assign new_new_n944__ = ~new_new_n932__ & new_new_n943__;
  assign new_new_n945__ = ~new_new_n679__ & ~new_new_n688__;
  assign new_new_n946__ = ~new_new_n678__ & new_new_n945__;
  assign new_new_n947__ = ~new_new_n689__ & ~new_new_n946__;
  assign new_new_n948__ = ~new_new_n745__ & new_new_n947__;
  assign new_new_n949__ = ~new_new_n944__ & new_new_n948__;
  assign new_new_n950__ = ~new_new_n631__ & ~new_new_n663__;
  assign new_new_n951__ = ~new_new_n664__ & ~new_new_n665__;
  assign new_new_n952__ = new_new_n950__ & new_new_n951__;
  assign new_new_n953__ = new_new_n657__ & new_new_n952__;
  assign new_new_n954__ = ~new_new_n949__ & new_new_n953__;
  assign new_new_n955__ = ~G1455 & ~G2204;
  assign new_new_n956__ = G4528 & new_new_n955__;
  assign new_new_n957__ = G38 & ~new_new_n956__;
  assign new_new_n958__ = new_new_n631__ & new_new_n657__;
  assign new_new_n959__ = new_new_n638__ & ~new_new_n653__;
  assign new_new_n960__ = new_new_n651__ & ~new_new_n959__;
  assign new_new_n961__ = ~new_new_n652__ & ~new_new_n960__;
  assign new_new_n962__ = ~new_new_n958__ & ~new_new_n961__;
  assign new_new_n963__ = ~new_new_n663__ & ~new_new_n962__;
  assign new_new_n964__ = ~new_new_n664__ & ~new_new_n957__;
  assign new_new_n965__ = ~new_new_n963__ & new_new_n964__;
  assign new_new_n966__ = ~new_new_n954__ & new_new_n965__;
  assign new_new_n967__ = G1455 & G2204;
  assign new_new_n968__ = ~G38 & G4528;
  assign new_new_n969__ = ~new_new_n967__ & new_new_n968__;
  assign G258 = ~new_new_n966__ & ~new_new_n969__;
  assign new_new_n971__ = ~new_new_n410__ & ~new_new_n434__;
  assign new_new_n972__ = new_new_n435__ & new_new_n439__;
  assign new_new_n973__ = new_new_n436__ & new_new_n972__;
  assign new_new_n974__ = ~new_new_n432__ & ~new_new_n973__;
  assign new_new_n975__ = new_new_n971__ & ~new_new_n974__;
  assign new_new_n976__ = ~new_new_n971__ & new_new_n974__;
  assign G388 = ~new_new_n975__ & ~new_new_n976__;
  assign new_new_n978__ = ~new_new_n430__ & ~new_new_n972__;
  assign new_new_n979__ = new_new_n436__ & ~new_new_n978__;
  assign new_new_n980__ = ~new_new_n436__ & new_new_n978__;
  assign G391 = ~new_new_n979__ & ~new_new_n980__;
  assign new_new_n982__ = ~new_new_n423__ & ~new_new_n426__;
  assign new_new_n983__ = ~new_new_n439__ & new_new_n982__;
  assign new_new_n984__ = new_new_n435__ & ~new_new_n983__;
  assign new_new_n985__ = ~new_new_n435__ & new_new_n983__;
  assign G394 = ~new_new_n984__ & ~new_new_n985__;
  assign new_new_n987__ = ~new_new_n334__ & ~new_new_n340__;
  assign new_new_n988__ = new_new_n425__ & ~new_new_n987__;
  assign new_new_n989__ = ~new_new_n425__ & new_new_n987__;
  assign G397 = ~new_new_n988__ & ~new_new_n989__;
  assign new_new_n991__ = ~new_new_n443__ & new_new_n456__;
  assign new_new_n992__ = new_new_n473__ & ~new_new_n991__;
  assign new_new_n993__ = ~new_new_n461__ & ~new_new_n992__;
  assign new_new_n994__ = ~new_new_n460__ & ~new_new_n993__;
  assign new_new_n995__ = new_new_n468__ & ~new_new_n994__;
  assign new_new_n996__ = ~new_new_n468__ & new_new_n994__;
  assign G376 = ~new_new_n995__ & ~new_new_n996__;
  assign new_new_n998__ = new_new_n462__ & ~new_new_n992__;
  assign new_new_n999__ = ~new_new_n462__ & new_new_n992__;
  assign G379 = ~new_new_n998__ & ~new_new_n999__;
  assign new_new_n1001__ = ~new_new_n443__ & ~new_new_n454__;
  assign new_new_n1002__ = ~new_new_n453__ & ~new_new_n1001__;
  assign new_new_n1003__ = new_new_n449__ & ~new_new_n1002__;
  assign new_new_n1004__ = ~new_new_n449__ & new_new_n1002__;
  assign G382 = ~new_new_n1003__ & ~new_new_n1004__;
  assign new_new_n1006__ = ~new_new_n443__ & new_new_n455__;
  assign new_new_n1007__ = new_new_n443__ & ~new_new_n455__;
  assign G385 = ~new_new_n1006__ & ~new_new_n1007__;
  assign new_new_n1009__ = new_new_n358__ & ~new_new_n364__;
  assign new_new_n1010__ = ~new_new_n358__ & new_new_n364__;
  assign new_new_n1011__ = ~new_new_n1009__ & ~new_new_n1010__;
  assign new_new_n1012__ = ~G18 & G141;
  assign new_new_n1013__ = G18 & G161;
  assign new_new_n1014__ = ~new_new_n1012__ & ~new_new_n1013__;
  assign new_new_n1015__ = new_new_n352__ & ~new_new_n376__;
  assign new_new_n1016__ = ~new_new_n352__ & new_new_n376__;
  assign new_new_n1017__ = ~new_new_n1015__ & ~new_new_n1016__;
  assign new_new_n1018__ = new_new_n1014__ & new_new_n1017__;
  assign new_new_n1019__ = ~new_new_n1014__ & ~new_new_n1017__;
  assign new_new_n1020__ = ~new_new_n1018__ & ~new_new_n1019__;
  assign new_new_n1021__ = new_new_n389__ & new_new_n395__;
  assign new_new_n1022__ = new_new_n390__ & new_new_n394__;
  assign new_new_n1023__ = ~new_new_n1021__ & ~new_new_n1022__;
  assign new_new_n1024__ = new_new_n385__ & new_new_n400__;
  assign new_new_n1025__ = new_new_n384__ & new_new_n401__;
  assign new_new_n1026__ = ~new_new_n1024__ & ~new_new_n1025__;
  assign new_new_n1027__ = ~new_new_n1023__ & new_new_n1026__;
  assign new_new_n1028__ = new_new_n1023__ & ~new_new_n1026__;
  assign new_new_n1029__ = ~new_new_n1027__ & ~new_new_n1028__;
  assign new_new_n1030__ = new_new_n370__ & ~new_new_n1029__;
  assign new_new_n1031__ = ~new_new_n370__ & new_new_n1029__;
  assign new_new_n1032__ = ~new_new_n1030__ & ~new_new_n1031__;
  assign new_new_n1033__ = ~new_new_n1020__ & new_new_n1032__;
  assign new_new_n1034__ = new_new_n1020__ & ~new_new_n1032__;
  assign new_new_n1035__ = ~new_new_n1033__ & ~new_new_n1034__;
  assign new_new_n1036__ = new_new_n1011__ & ~new_new_n1035__;
  assign new_new_n1037__ = ~new_new_n1011__ & new_new_n1035__;
  assign new_new_n1038__ = ~new_new_n1036__ & ~new_new_n1037__;
  assign new_new_n1039__ = ~new_new_n528__ & new_new_n541__;
  assign new_new_n1040__ = new_new_n528__ & ~new_new_n541__;
  assign new_new_n1041__ = ~new_new_n1039__ & ~new_new_n1040__;
  assign new_new_n1042__ = new_new_n534__ & ~new_new_n547__;
  assign new_new_n1043__ = ~new_new_n534__ & new_new_n547__;
  assign new_new_n1044__ = ~new_new_n1042__ & ~new_new_n1043__;
  assign new_new_n1045__ = new_new_n1041__ & new_new_n1044__;
  assign new_new_n1046__ = ~new_new_n1041__ & ~new_new_n1044__;
  assign new_new_n1047__ = ~new_new_n1045__ & ~new_new_n1046__;
  assign new_new_n1048__ = new_new_n493__ & ~new_new_n1047__;
  assign new_new_n1049__ = ~new_new_n493__ & new_new_n1047__;
  assign new_new_n1050__ = ~new_new_n1048__ & ~new_new_n1049__;
  assign new_new_n1051__ = new_new_n481__ & ~new_new_n497__;
  assign new_new_n1052__ = ~new_new_n481__ & new_new_n497__;
  assign new_new_n1053__ = ~new_new_n1051__ & ~new_new_n1052__;
  assign new_new_n1054__ = new_new_n487__ & new_new_n1053__;
  assign new_new_n1055__ = ~new_new_n487__ & ~new_new_n1053__;
  assign new_new_n1056__ = ~new_new_n1054__ & ~new_new_n1055__;
  assign new_new_n1057__ = G18 & G227;
  assign new_new_n1058__ = ~G18 & G115;
  assign new_new_n1059__ = ~new_new_n1057__ & ~new_new_n1058__;
  assign new_new_n1060__ = new_new_n504__ & ~new_new_n1059__;
  assign new_new_n1061__ = ~new_new_n504__ & new_new_n1059__;
  assign new_new_n1062__ = ~new_new_n1060__ & ~new_new_n1061__;
  assign new_new_n1063__ = new_new_n1056__ & ~new_new_n1062__;
  assign new_new_n1064__ = ~new_new_n1056__ & new_new_n1062__;
  assign new_new_n1065__ = ~new_new_n1063__ & ~new_new_n1064__;
  assign new_new_n1066__ = new_new_n1050__ & new_new_n1065__;
  assign new_new_n1067__ = ~new_new_n1050__ & ~new_new_n1065__;
  assign new_new_n1068__ = new_new_n446__ & ~new_new_n465__;
  assign new_new_n1069__ = ~new_new_n446__ & new_new_n465__;
  assign new_new_n1070__ = ~new_new_n1068__ & ~new_new_n1069__;
  assign new_new_n1071__ = new_new_n452__ & ~new_new_n459__;
  assign new_new_n1072__ = ~new_new_n452__ & new_new_n459__;
  assign new_new_n1073__ = ~new_new_n1071__ & ~new_new_n1072__;
  assign new_new_n1074__ = new_new_n1070__ & new_new_n1073__;
  assign new_new_n1075__ = ~new_new_n1070__ & ~new_new_n1073__;
  assign new_new_n1076__ = ~new_new_n1074__ & ~new_new_n1075__;
  assign new_new_n1077__ = new_new_n413__ & ~new_new_n1076__;
  assign new_new_n1078__ = ~new_new_n413__ & new_new_n1076__;
  assign new_new_n1079__ = ~new_new_n1077__ & ~new_new_n1078__;
  assign new_new_n1080__ = G18 & G239;
  assign new_new_n1081__ = ~G18 & G44;
  assign new_new_n1082__ = ~new_new_n1080__ & ~new_new_n1081__;
  assign new_new_n1083__ = new_new_n418__ & ~new_new_n1082__;
  assign new_new_n1084__ = ~new_new_n418__ & new_new_n1082__;
  assign new_new_n1085__ = ~new_new_n1083__ & ~new_new_n1084__;
  assign new_new_n1086__ = new_new_n422__ & new_new_n1085__;
  assign new_new_n1087__ = ~new_new_n422__ & ~new_new_n1085__;
  assign new_new_n1088__ = ~new_new_n1086__ & ~new_new_n1087__;
  assign new_new_n1089__ = new_new_n336__ & ~new_new_n409__;
  assign new_new_n1090__ = ~new_new_n336__ & new_new_n409__;
  assign new_new_n1091__ = ~new_new_n1089__ & ~new_new_n1090__;
  assign new_new_n1092__ = new_new_n1088__ & ~new_new_n1091__;
  assign new_new_n1093__ = ~new_new_n1088__ & new_new_n1091__;
  assign new_new_n1094__ = ~new_new_n1092__ & ~new_new_n1093__;
  assign new_new_n1095__ = new_new_n1079__ & new_new_n1094__;
  assign new_new_n1096__ = ~new_new_n1079__ & ~new_new_n1094__;
  assign new_new_n1097__ = G211 & G212;
  assign new_new_n1098__ = G18 & ~new_new_n350__;
  assign new_new_n1099__ = ~G211 & ~G212;
  assign new_new_n1100__ = ~new_new_n1097__ & ~new_new_n1099__;
  assign new_new_n1101__ = new_new_n1098__ & new_new_n1100__;
  assign new_new_n1102__ = ~new_new_n350__ & new_new_n593__;
  assign new_new_n1103__ = new_new_n580__ & new_new_n586__;
  assign new_new_n1104__ = new_new_n581__ & new_new_n585__;
  assign new_new_n1105__ = ~new_new_n1103__ & ~new_new_n1104__;
  assign new_new_n1106__ = new_new_n591__ & new_new_n599__;
  assign new_new_n1107__ = new_new_n590__ & new_new_n600__;
  assign new_new_n1108__ = ~new_new_n1106__ & ~new_new_n1107__;
  assign new_new_n1109__ = new_new_n1105__ & ~new_new_n1108__;
  assign new_new_n1110__ = ~new_new_n1105__ & new_new_n1108__;
  assign new_new_n1111__ = ~new_new_n1109__ & ~new_new_n1110__;
  assign new_new_n1112__ = new_new_n1102__ & ~new_new_n1111__;
  assign new_new_n1113__ = ~new_new_n1102__ & new_new_n1111__;
  assign new_new_n1114__ = ~new_new_n1112__ & ~new_new_n1113__;
  assign new_new_n1115__ = new_new_n1101__ & new_new_n1114__;
  assign new_new_n1116__ = ~new_new_n1101__ & ~new_new_n1114__;
  assign new_new_n1117__ = ~new_new_n1115__ & ~new_new_n1116__;
  assign new_new_n1118__ = ~new_new_n1066__ & ~new_new_n1067__;
  assign new_new_n1119__ = ~new_new_n1095__ & ~new_new_n1096__;
  assign new_new_n1120__ = new_new_n1118__ & new_new_n1119__;
  assign new_new_n1121__ = ~new_new_n1117__ & new_new_n1120__;
  assign G412 = new_new_n1038__ | ~new_new_n1121__;
  assign new_new_n1123__ = ~new_new_n630__ & new_new_n662__;
  assign new_new_n1124__ = new_new_n630__ & ~new_new_n662__;
  assign new_new_n1125__ = ~new_new_n1123__ & ~new_new_n1124__;
  assign new_new_n1126__ = new_new_n643__ & new_new_n1125__;
  assign new_new_n1127__ = ~new_new_n643__ & ~new_new_n1125__;
  assign new_new_n1128__ = ~new_new_n1126__ & ~new_new_n1127__;
  assign new_new_n1129__ = ~new_new_n636__ & ~new_new_n649__;
  assign new_new_n1130__ = new_new_n636__ & new_new_n649__;
  assign new_new_n1131__ = ~new_new_n1129__ & ~new_new_n1130__;
  assign new_new_n1132__ = G18 & ~G1459;
  assign new_new_n1133__ = ~G18 & G114;
  assign new_new_n1134__ = ~new_new_n1132__ & ~new_new_n1133__;
  assign new_new_n1135__ = new_new_n1131__ & ~new_new_n1134__;
  assign new_new_n1136__ = ~new_new_n1131__ & new_new_n1134__;
  assign new_new_n1137__ = ~new_new_n1135__ & ~new_new_n1136__;
  assign new_new_n1138__ = ~G1492 & ~G1496;
  assign new_new_n1139__ = G1492 & G1496;
  assign new_new_n1140__ = ~new_new_n1138__ & ~new_new_n1139__;
  assign new_new_n1141__ = G18 & ~new_new_n1140__;
  assign new_new_n1142__ = ~new_new_n955__ & ~new_new_n967__;
  assign new_new_n1143__ = ~G18 & ~new_new_n1142__;
  assign new_new_n1144__ = ~new_new_n1141__ & ~new_new_n1143__;
  assign new_new_n1145__ = ~new_new_n1137__ & new_new_n1144__;
  assign new_new_n1146__ = new_new_n1137__ & ~new_new_n1144__;
  assign new_new_n1147__ = ~new_new_n1145__ & ~new_new_n1146__;
  assign new_new_n1148__ = ~new_new_n1128__ & new_new_n1147__;
  assign new_new_n1149__ = new_new_n1128__ & ~new_new_n1147__;
  assign new_new_n1150__ = ~new_new_n1148__ & ~new_new_n1149__;
  assign new_new_n1151__ = ~G18 & G70;
  assign new_new_n1152__ = G18 & ~G3701;
  assign new_new_n1153__ = ~new_new_n1151__ & ~new_new_n1152__;
  assign new_new_n1154__ = new_new_n870__ & ~new_new_n876__;
  assign new_new_n1155__ = ~new_new_n870__ & new_new_n876__;
  assign new_new_n1156__ = ~new_new_n1154__ & ~new_new_n1155__;
  assign new_new_n1157__ = new_new_n1153__ & new_new_n1156__;
  assign new_new_n1158__ = ~new_new_n1153__ & ~new_new_n1156__;
  assign new_new_n1159__ = ~new_new_n1157__ & ~new_new_n1158__;
  assign new_new_n1160__ = G18 & ~G3698;
  assign new_new_n1161__ = ~G18 & G69;
  assign new_new_n1162__ = ~new_new_n1160__ & ~new_new_n1161__;
  assign new_new_n1163__ = ~new_new_n864__ & ~new_new_n891__;
  assign new_new_n1164__ = new_new_n864__ & new_new_n891__;
  assign new_new_n1165__ = ~new_new_n1163__ & ~new_new_n1164__;
  assign new_new_n1166__ = ~new_new_n830__ & new_new_n848__;
  assign new_new_n1167__ = new_new_n830__ & ~new_new_n848__;
  assign new_new_n1168__ = ~new_new_n1166__ & ~new_new_n1167__;
  assign new_new_n1169__ = ~new_new_n837__ & new_new_n855__;
  assign new_new_n1170__ = new_new_n837__ & ~new_new_n855__;
  assign new_new_n1171__ = ~new_new_n1169__ & ~new_new_n1170__;
  assign new_new_n1172__ = new_new_n1168__ & new_new_n1171__;
  assign new_new_n1173__ = ~new_new_n1168__ & ~new_new_n1171__;
  assign new_new_n1174__ = ~new_new_n1172__ & ~new_new_n1173__;
  assign new_new_n1175__ = new_new_n1165__ & ~new_new_n1174__;
  assign new_new_n1176__ = ~new_new_n1165__ & new_new_n1174__;
  assign new_new_n1177__ = ~new_new_n1175__ & ~new_new_n1176__;
  assign new_new_n1178__ = new_new_n1162__ & new_new_n1177__;
  assign new_new_n1179__ = ~new_new_n1162__ & ~new_new_n1177__;
  assign new_new_n1180__ = ~new_new_n1178__ & ~new_new_n1179__;
  assign new_new_n1181__ = ~new_new_n1159__ & ~new_new_n1180__;
  assign new_new_n1182__ = new_new_n786__ & ~new_new_n792__;
  assign new_new_n1183__ = ~new_new_n786__ & new_new_n792__;
  assign new_new_n1184__ = ~new_new_n1182__ & ~new_new_n1183__;
  assign new_new_n1185__ = new_new_n805__ & new_new_n1184__;
  assign new_new_n1186__ = ~new_new_n805__ & ~new_new_n1184__;
  assign new_new_n1187__ = ~new_new_n1185__ & ~new_new_n1186__;
  assign new_new_n1188__ = G18 & ~G4393;
  assign new_new_n1189__ = ~G18 & G58;
  assign new_new_n1190__ = ~new_new_n1188__ & ~new_new_n1189__;
  assign new_new_n1191__ = ~new_new_n798__ & ~new_new_n812__;
  assign new_new_n1192__ = new_new_n798__ & new_new_n812__;
  assign new_new_n1193__ = ~new_new_n1191__ & ~new_new_n1192__;
  assign new_new_n1194__ = new_new_n766__ & ~new_new_n772__;
  assign new_new_n1195__ = ~new_new_n766__ & new_new_n772__;
  assign new_new_n1196__ = ~new_new_n1194__ & ~new_new_n1195__;
  assign new_new_n1197__ = new_new_n751__ & ~new_new_n759__;
  assign new_new_n1198__ = ~new_new_n751__ & new_new_n759__;
  assign new_new_n1199__ = ~new_new_n1197__ & ~new_new_n1198__;
  assign new_new_n1200__ = new_new_n1196__ & new_new_n1199__;
  assign new_new_n1201__ = ~new_new_n1196__ & ~new_new_n1199__;
  assign new_new_n1202__ = ~new_new_n1200__ & ~new_new_n1201__;
  assign new_new_n1203__ = new_new_n1193__ & ~new_new_n1202__;
  assign new_new_n1204__ = ~new_new_n1193__ & new_new_n1202__;
  assign new_new_n1205__ = ~new_new_n1203__ & ~new_new_n1204__;
  assign new_new_n1206__ = new_new_n1190__ & new_new_n1205__;
  assign new_new_n1207__ = ~new_new_n1190__ & ~new_new_n1205__;
  assign new_new_n1208__ = ~new_new_n1206__ & ~new_new_n1207__;
  assign new_new_n1209__ = ~new_new_n1187__ & new_new_n1208__;
  assign new_new_n1210__ = new_new_n1187__ & ~new_new_n1208__;
  assign new_new_n1211__ = new_new_n1159__ & new_new_n1180__;
  assign new_new_n1212__ = ~new_new_n718__ & ~new_new_n726__;
  assign new_new_n1213__ = new_new_n718__ & new_new_n726__;
  assign new_new_n1214__ = ~new_new_n1212__ & ~new_new_n1213__;
  assign new_new_n1215__ = new_new_n670__ & ~new_new_n676__;
  assign new_new_n1216__ = ~new_new_n670__ & new_new_n676__;
  assign new_new_n1217__ = ~new_new_n1215__ & ~new_new_n1216__;
  assign new_new_n1218__ = new_new_n687__ & ~new_new_n695__;
  assign new_new_n1219__ = ~new_new_n687__ & new_new_n695__;
  assign new_new_n1220__ = ~new_new_n1218__ & ~new_new_n1219__;
  assign new_new_n1221__ = new_new_n1217__ & new_new_n1220__;
  assign new_new_n1222__ = ~new_new_n1217__ & ~new_new_n1220__;
  assign new_new_n1223__ = ~new_new_n1221__ & ~new_new_n1222__;
  assign new_new_n1224__ = new_new_n1214__ & ~new_new_n1223__;
  assign new_new_n1225__ = ~new_new_n1214__ & new_new_n1223__;
  assign new_new_n1226__ = ~new_new_n1224__ & ~new_new_n1225__;
  assign new_new_n1227__ = new_new_n705__ & ~new_new_n733__;
  assign new_new_n1228__ = ~new_new_n705__ & new_new_n733__;
  assign new_new_n1229__ = ~new_new_n1227__ & ~new_new_n1228__;
  assign new_new_n1230__ = new_new_n711__ & new_new_n1229__;
  assign new_new_n1231__ = ~new_new_n711__ & ~new_new_n1229__;
  assign new_new_n1232__ = ~new_new_n1230__ & ~new_new_n1231__;
  assign new_new_n1233__ = G18 & ~G2208;
  assign new_new_n1234__ = ~G18 & G82;
  assign new_new_n1235__ = ~new_new_n1233__ & ~new_new_n1234__;
  assign new_new_n1236__ = new_new_n1232__ & ~new_new_n1235__;
  assign new_new_n1237__ = ~new_new_n1232__ & new_new_n1235__;
  assign new_new_n1238__ = ~new_new_n1236__ & ~new_new_n1237__;
  assign new_new_n1239__ = new_new_n1226__ & new_new_n1238__;
  assign new_new_n1240__ = ~new_new_n1226__ & ~new_new_n1238__;
  assign new_new_n1241__ = ~new_new_n1239__ & ~new_new_n1240__;
  assign new_new_n1242__ = ~new_new_n1150__ & new_new_n1241__;
  assign new_new_n1243__ = ~new_new_n1181__ & new_new_n1242__;
  assign new_new_n1244__ = ~new_new_n1209__ & ~new_new_n1210__;
  assign new_new_n1245__ = ~new_new_n1211__ & new_new_n1244__;
  assign G414 = ~new_new_n1243__ | ~new_new_n1245__;
  assign new_new_n1247__ = G18 & ~G170;
  assign new_new_n1248__ = ~new_new_n658__ & ~new_new_n1247__;
  assign new_new_n1249__ = new_new_n658__ & new_new_n1247__;
  assign new_new_n1250__ = ~new_new_n1248__ & ~new_new_n1249__;
  assign new_new_n1251__ = new_new_n639__ & new_new_n1250__;
  assign new_new_n1252__ = ~new_new_n639__ & ~new_new_n1250__;
  assign new_new_n1253__ = ~new_new_n350__ & ~new_new_n1251__;
  assign new_new_n1254__ = ~new_new_n1252__ & new_new_n1253__;
  assign new_new_n1255__ = new_new_n633__ & new_new_n645__;
  assign new_new_n1256__ = new_new_n632__ & new_new_n646__;
  assign new_new_n1257__ = ~new_new_n1255__ & ~new_new_n1256__;
  assign new_new_n1258__ = G164 & G165;
  assign new_new_n1259__ = ~G164 & ~G165;
  assign new_new_n1260__ = ~new_new_n1258__ & ~new_new_n1259__;
  assign new_new_n1261__ = new_new_n1098__ & new_new_n1260__;
  assign new_new_n1262__ = ~new_new_n1257__ & ~new_new_n1261__;
  assign new_new_n1263__ = new_new_n1257__ & new_new_n1261__;
  assign new_new_n1264__ = ~new_new_n1262__ & ~new_new_n1263__;
  assign new_new_n1265__ = new_new_n1254__ & ~new_new_n1264__;
  assign new_new_n1266__ = ~new_new_n1254__ & new_new_n1264__;
  assign new_new_n1267__ = ~new_new_n1265__ & ~new_new_n1266__;
  assign new_new_n1268__ = new_new_n763__ & ~new_new_n769__;
  assign new_new_n1269__ = ~new_new_n763__ & new_new_n769__;
  assign new_new_n1270__ = ~new_new_n1268__ & ~new_new_n1269__;
  assign new_new_n1271__ = new_new_n748__ & ~new_new_n756__;
  assign new_new_n1272__ = ~new_new_n748__ & new_new_n756__;
  assign new_new_n1273__ = ~new_new_n1271__ & ~new_new_n1272__;
  assign new_new_n1274__ = new_new_n1270__ & new_new_n1273__;
  assign new_new_n1275__ = ~new_new_n1270__ & ~new_new_n1273__;
  assign new_new_n1276__ = ~new_new_n1274__ & ~new_new_n1275__;
  assign new_new_n1277__ = new_new_n795__ & ~new_new_n1276__;
  assign new_new_n1278__ = ~new_new_n795__ & new_new_n1276__;
  assign new_new_n1279__ = ~new_new_n1277__ & ~new_new_n1278__;
  assign new_new_n1280__ = new_new_n783__ & ~new_new_n789__;
  assign new_new_n1281__ = ~new_new_n783__ & new_new_n789__;
  assign new_new_n1282__ = ~new_new_n1280__ & ~new_new_n1281__;
  assign new_new_n1283__ = new_new_n802__ & new_new_n1282__;
  assign new_new_n1284__ = ~new_new_n802__ & ~new_new_n1282__;
  assign new_new_n1285__ = ~new_new_n1283__ & ~new_new_n1284__;
  assign new_new_n1286__ = G18 & G197;
  assign new_new_n1287__ = ~new_new_n1058__ & ~new_new_n1286__;
  assign new_new_n1288__ = new_new_n809__ & ~new_new_n1287__;
  assign new_new_n1289__ = ~new_new_n809__ & new_new_n1287__;
  assign new_new_n1290__ = ~new_new_n1288__ & ~new_new_n1289__;
  assign new_new_n1291__ = new_new_n1285__ & ~new_new_n1290__;
  assign new_new_n1292__ = ~new_new_n1285__ & new_new_n1290__;
  assign new_new_n1293__ = ~new_new_n1291__ & ~new_new_n1292__;
  assign new_new_n1294__ = new_new_n1279__ & new_new_n1293__;
  assign new_new_n1295__ = ~new_new_n1279__ & ~new_new_n1293__;
  assign new_new_n1296__ = ~new_new_n827__ & new_new_n845__;
  assign new_new_n1297__ = new_new_n827__ & ~new_new_n845__;
  assign new_new_n1298__ = ~new_new_n1296__ & ~new_new_n1297__;
  assign new_new_n1299__ = ~new_new_n834__ & new_new_n852__;
  assign new_new_n1300__ = new_new_n834__ & ~new_new_n852__;
  assign new_new_n1301__ = ~new_new_n1299__ & ~new_new_n1300__;
  assign new_new_n1302__ = new_new_n1298__ & new_new_n1301__;
  assign new_new_n1303__ = ~new_new_n1298__ & ~new_new_n1301__;
  assign new_new_n1304__ = ~new_new_n1302__ & ~new_new_n1303__;
  assign new_new_n1305__ = new_new_n861__ & ~new_new_n1304__;
  assign new_new_n1306__ = ~new_new_n861__ & new_new_n1304__;
  assign new_new_n1307__ = ~new_new_n1305__ & ~new_new_n1306__;
  assign new_new_n1308__ = G18 & G208;
  assign new_new_n1309__ = ~new_new_n1081__ & ~new_new_n1308__;
  assign new_new_n1310__ = new_new_n867__ & ~new_new_n1309__;
  assign new_new_n1311__ = ~new_new_n867__ & new_new_n1309__;
  assign new_new_n1312__ = ~new_new_n1310__ & ~new_new_n1311__;
  assign new_new_n1313__ = new_new_n873__ & new_new_n1312__;
  assign new_new_n1314__ = ~new_new_n873__ & ~new_new_n1312__;
  assign new_new_n1315__ = ~new_new_n1313__ & ~new_new_n1314__;
  assign new_new_n1316__ = G18 & G198;
  assign new_new_n1317__ = ~new_new_n333__ & ~new_new_n1316__;
  assign new_new_n1318__ = new_new_n888__ & ~new_new_n1317__;
  assign new_new_n1319__ = ~new_new_n888__ & new_new_n1317__;
  assign new_new_n1320__ = ~new_new_n1318__ & ~new_new_n1319__;
  assign new_new_n1321__ = new_new_n1315__ & ~new_new_n1320__;
  assign new_new_n1322__ = ~new_new_n1315__ & new_new_n1320__;
  assign new_new_n1323__ = ~new_new_n1321__ & ~new_new_n1322__;
  assign new_new_n1324__ = new_new_n1307__ & new_new_n1323__;
  assign new_new_n1325__ = ~new_new_n1307__ & ~new_new_n1323__;
  assign new_new_n1326__ = G18 & G181;
  assign new_new_n1327__ = ~new_new_n1012__ & ~new_new_n1326__;
  assign new_new_n1328__ = new_new_n708__ & ~new_new_n730__;
  assign new_new_n1329__ = ~new_new_n708__ & new_new_n730__;
  assign new_new_n1330__ = ~new_new_n1328__ & ~new_new_n1329__;
  assign new_new_n1331__ = new_new_n1327__ & new_new_n1330__;
  assign new_new_n1332__ = ~new_new_n1327__ & ~new_new_n1330__;
  assign new_new_n1333__ = ~new_new_n1331__ & ~new_new_n1332__;
  assign new_new_n1334__ = new_new_n702__ & ~new_new_n715__;
  assign new_new_n1335__ = ~new_new_n702__ & new_new_n715__;
  assign new_new_n1336__ = ~new_new_n1334__ & ~new_new_n1335__;
  assign new_new_n1337__ = new_new_n672__ & new_new_n692__;
  assign new_new_n1338__ = new_new_n673__ & new_new_n691__;
  assign new_new_n1339__ = ~new_new_n1337__ & ~new_new_n1338__;
  assign new_new_n1340__ = new_new_n667__ & new_new_n683__;
  assign new_new_n1341__ = new_new_n666__ & new_new_n684__;
  assign new_new_n1342__ = ~new_new_n1340__ & ~new_new_n1341__;
  assign new_new_n1343__ = ~new_new_n1339__ & new_new_n1342__;
  assign new_new_n1344__ = new_new_n1339__ & ~new_new_n1342__;
  assign new_new_n1345__ = ~new_new_n1343__ & ~new_new_n1344__;
  assign new_new_n1346__ = new_new_n723__ & ~new_new_n1345__;
  assign new_new_n1347__ = ~new_new_n723__ & new_new_n1345__;
  assign new_new_n1348__ = ~new_new_n1346__ & ~new_new_n1347__;
  assign new_new_n1349__ = new_new_n1336__ & new_new_n1348__;
  assign new_new_n1350__ = ~new_new_n1336__ & ~new_new_n1348__;
  assign new_new_n1351__ = ~new_new_n1349__ & ~new_new_n1350__;
  assign new_new_n1352__ = new_new_n1333__ & ~new_new_n1351__;
  assign new_new_n1353__ = ~new_new_n1333__ & new_new_n1351__;
  assign new_new_n1354__ = ~new_new_n1267__ & ~new_new_n1294__;
  assign new_new_n1355__ = ~new_new_n1295__ & ~new_new_n1324__;
  assign new_new_n1356__ = ~new_new_n1325__ & new_new_n1355__;
  assign new_new_n1357__ = new_new_n1354__ & new_new_n1356__;
  assign new_new_n1358__ = ~new_new_n1352__ & ~new_new_n1353__;
  assign G416 = ~new_new_n1357__ | ~new_new_n1358__;
  assign new_new_n1360__ = new_new_n379__ & ~new_new_n560__;
  assign new_new_n1361__ = ~new_new_n379__ & new_new_n560__;
  assign G295 = ~new_new_n1360__ & ~new_new_n1361__;
  assign new_new_n1363__ = ~new_new_n579__ & new_new_n597__;
  assign new_new_n1364__ = new_new_n579__ & ~new_new_n597__;
  assign G324 = ~new_new_n1363__ & ~new_new_n1364__;
  assign new_new_n1366__ = new_new_n825__ & ~new_new_n915__;
  assign new_new_n1367__ = new_new_n923__ & ~new_new_n1366__;
  assign new_new_n1368__ = new_new_n781__ & ~new_new_n1367__;
  assign G252 = ~new_new_n930__ | new_new_n1368__;
  assign new_new_n1370__ = ~new_new_n382__ & new_new_n573__;
  assign new_new_n1371__ = new_new_n560__ & new_new_n573__;
  assign new_new_n1372__ = ~new_new_n1370__ & ~new_new_n1371__;
  assign new_new_n1373__ = new_new_n355__ & ~new_new_n1372__;
  assign new_new_n1374__ = ~new_new_n355__ & new_new_n1372__;
  assign G310 = new_new_n1373__ | new_new_n1374__;
  assign new_new_n1376__ = new_new_n380__ & ~new_new_n560__;
  assign new_new_n1377__ = new_new_n367__ & new_new_n1376__;
  assign new_new_n1378__ = ~new_new_n571__ & ~new_new_n1377__;
  assign new_new_n1379__ = new_new_n361__ & ~new_new_n1378__;
  assign new_new_n1380__ = ~new_new_n361__ & new_new_n1378__;
  assign G313 = ~new_new_n1379__ & ~new_new_n1380__;
  assign new_new_n1382__ = ~new_new_n371__ & ~new_new_n568__;
  assign new_new_n1383__ = ~new_new_n1376__ & new_new_n1382__;
  assign new_new_n1384__ = new_new_n367__ & ~new_new_n1383__;
  assign new_new_n1385__ = ~new_new_n367__ & new_new_n1383__;
  assign G316 = ~new_new_n1384__ & ~new_new_n1385__;
  assign new_new_n1387__ = ~new_new_n377__ & ~new_new_n1360__;
  assign new_new_n1388__ = new_new_n373__ & ~new_new_n1387__;
  assign new_new_n1389__ = ~new_new_n373__ & new_new_n1387__;
  assign G319 = ~new_new_n1388__ & ~new_new_n1389__;
  assign new_new_n1391__ = new_new_n614__ & ~new_new_n616__;
  assign new_new_n1392__ = ~new_new_n588__ & ~new_new_n1391__;
  assign new_new_n1393__ = ~new_new_n587__ & ~new_new_n1392__;
  assign new_new_n1394__ = ~new_new_n579__ & new_new_n606__;
  assign new_new_n1395__ = new_new_n589__ & new_new_n1394__;
  assign new_new_n1396__ = new_new_n1393__ & ~new_new_n1395__;
  assign new_new_n1397__ = new_new_n584__ & new_new_n1396__;
  assign new_new_n1398__ = ~new_new_n584__ & ~new_new_n1396__;
  assign G327 = new_new_n1397__ | new_new_n1398__;
  assign new_new_n1400__ = new_new_n1391__ & ~new_new_n1394__;
  assign new_new_n1401__ = new_new_n589__ & new_new_n1400__;
  assign new_new_n1402__ = ~new_new_n589__ & ~new_new_n1400__;
  assign G330 = new_new_n1401__ | new_new_n1402__;
  assign new_new_n1404__ = ~new_new_n595__ & ~new_new_n1363__;
  assign new_new_n1405__ = new_new_n611__ & ~new_new_n1404__;
  assign new_new_n1406__ = ~new_new_n604__ & ~new_new_n1405__;
  assign new_new_n1407__ = new_new_n603__ & new_new_n1406__;
  assign new_new_n1408__ = ~new_new_n603__ & ~new_new_n1406__;
  assign G333 = new_new_n1407__ | new_new_n1408__;
  assign new_new_n1410__ = ~new_new_n611__ & new_new_n1404__;
  assign G336 = ~new_new_n1405__ & ~new_new_n1410__;
  assign new_new_n1412__ = ~G404 & ~G406;
  assign new_new_n1413__ = ~G408 & ~G410;
  assign new_new_n1414__ = new_new_n1412__ & new_new_n1413__;
  assign new_new_n1415__ = ~G412 & new_new_n1414__;
  assign new_new_n1416__ = ~G416 & new_new_n1415__;
  assign G418 = G414 | ~new_new_n1416__;
  assign new_new_n1418__ = new_new_n383__ & ~new_new_n560__;
  assign new_new_n1419__ = new_new_n575__ & ~new_new_n1418__;
  assign new_new_n1420__ = new_new_n399__ & ~new_new_n1419__;
  assign new_new_n1421__ = ~new_new_n387__ & new_new_n1420__;
  assign new_new_n1422__ = ~new_new_n566__ & ~new_new_n1421__;
  assign new_new_n1423__ = new_new_n404__ & ~new_new_n1422__;
  assign new_new_n1424__ = ~new_new_n404__ & new_new_n1422__;
  assign G298 = ~new_new_n1423__ & ~new_new_n1424__;
  assign new_new_n1426__ = new_new_n564__ & ~new_new_n1420__;
  assign new_new_n1427__ = new_new_n388__ & ~new_new_n1426__;
  assign new_new_n1428__ = ~new_new_n388__ & new_new_n1426__;
  assign G301 = ~new_new_n1427__ & ~new_new_n1428__;
  assign new_new_n1430__ = ~new_new_n397__ & ~new_new_n1419__;
  assign new_new_n1431__ = ~new_new_n396__ & ~new_new_n1430__;
  assign new_new_n1432__ = new_new_n393__ & ~new_new_n1431__;
  assign new_new_n1433__ = ~new_new_n393__ & new_new_n1431__;
  assign G304 = ~new_new_n1432__ & ~new_new_n1433__;
  assign new_new_n1435__ = new_new_n398__ & ~new_new_n1419__;
  assign new_new_n1436__ = ~new_new_n398__ & new_new_n1419__;
  assign G307 = ~new_new_n1435__ & ~new_new_n1436__;
  assign new_new_n1438__ = ~new_new_n478__ & new_new_n500__;
  assign new_new_n1439__ = new_new_n478__ & ~new_new_n500__;
  assign G344 = ~new_new_n1438__ & ~new_new_n1439__;
  assign new_new_n1441__ = ~new_new_n347__ & new_new_n621__;
  assign new_new_n1442__ = ~new_new_n348__ & ~new_new_n1441__;
  assign new_new_n1443__ = ~new_new_n624__ & ~new_new_n1442__;
  assign new_new_n1444__ = new_new_n624__ & new_new_n1442__;
  assign G422 = new_new_n1443__ | new_new_n1444__;
  assign new_new_n1446__ = ~new_new_n349__ & ~new_new_n621__;
  assign new_new_n1447__ = new_new_n349__ & new_new_n621__;
  assign G419 = new_new_n1446__ | new_new_n1447__;
  assign new_new_n1449__ = new_new_n518__ & ~new_new_n520__;
  assign new_new_n1450__ = ~new_new_n489__ & ~new_new_n1449__;
  assign new_new_n1451__ = ~new_new_n488__ & ~new_new_n1450__;
  assign new_new_n1452__ = ~new_new_n478__ & new_new_n510__;
  assign new_new_n1453__ = new_new_n490__ & new_new_n1452__;
  assign new_new_n1454__ = new_new_n1451__ & ~new_new_n1453__;
  assign new_new_n1455__ = new_new_n484__ & ~new_new_n1454__;
  assign new_new_n1456__ = ~new_new_n484__ & new_new_n1454__;
  assign G359 = ~new_new_n1455__ & ~new_new_n1456__;
  assign new_new_n1458__ = new_new_n1449__ & ~new_new_n1452__;
  assign new_new_n1459__ = new_new_n490__ & ~new_new_n1458__;
  assign new_new_n1460__ = ~new_new_n490__ & new_new_n1458__;
  assign G362 = ~new_new_n1459__ & ~new_new_n1460__;
  assign new_new_n1462__ = ~new_new_n498__ & ~new_new_n1438__;
  assign new_new_n1463__ = new_new_n515__ & ~new_new_n1462__;
  assign new_new_n1464__ = ~new_new_n508__ & ~new_new_n1463__;
  assign new_new_n1465__ = new_new_n507__ & ~new_new_n1464__;
  assign new_new_n1466__ = ~new_new_n507__ & new_new_n1464__;
  assign G365 = ~new_new_n1465__ & ~new_new_n1466__;
  assign new_new_n1468__ = ~new_new_n515__ & new_new_n1462__;
  assign G368 = ~new_new_n1463__ & ~new_new_n1468__;
  assign new_new_n1470__ = ~new_new_n525__ & new_new_n538__;
  assign new_new_n1471__ = ~new_new_n548__ & new_new_n1470__;
  assign new_new_n1472__ = new_new_n557__ & ~new_new_n1471__;
  assign new_new_n1473__ = new_new_n544__ & ~new_new_n1472__;
  assign new_new_n1474__ = ~new_new_n544__ & new_new_n1472__;
  assign G347 = ~new_new_n1473__ & ~new_new_n1474__;
  assign new_new_n1476__ = new_new_n555__ & ~new_new_n1470__;
  assign new_new_n1477__ = new_new_n550__ & ~new_new_n1476__;
  assign new_new_n1478__ = ~new_new_n550__ & new_new_n1476__;
  assign G350 = ~new_new_n1477__ & ~new_new_n1478__;
  assign new_new_n1480__ = ~new_new_n525__ & ~new_new_n536__;
  assign new_new_n1481__ = ~new_new_n535__ & ~new_new_n1480__;
  assign new_new_n1482__ = new_new_n531__ & ~new_new_n1481__;
  assign new_new_n1483__ = ~new_new_n531__ & new_new_n1481__;
  assign G353 = ~new_new_n1482__ & ~new_new_n1483__;
  assign new_new_n1485__ = ~new_new_n525__ & new_new_n537__;
  assign new_new_n1486__ = new_new_n525__ & ~new_new_n537__;
  assign G356 = ~new_new_n1485__ & ~new_new_n1486__;
  assign new_new_n1488__ = ~new_new_n372__ & ~new_new_n377__;
  assign new_new_n1489__ = ~new_new_n371__ & ~new_new_n1488__;
  assign new_new_n1490__ = new_new_n573__ & ~new_new_n1489__;
  assign new_new_n1491__ = ~new_new_n573__ & new_new_n1489__;
  assign new_new_n1492__ = ~new_new_n1490__ & ~new_new_n1491__;
  assign new_new_n1493__ = new_new_n355__ & ~new_new_n1492__;
  assign new_new_n1494__ = ~new_new_n355__ & new_new_n1492__;
  assign new_new_n1495__ = ~new_new_n1493__ & ~new_new_n1494__;
  assign new_new_n1496__ = new_new_n361__ & ~new_new_n367__;
  assign new_new_n1497__ = ~new_new_n361__ & new_new_n367__;
  assign new_new_n1498__ = ~new_new_n1496__ & ~new_new_n1497__;
  assign new_new_n1499__ = new_new_n377__ & ~new_new_n571__;
  assign new_new_n1500__ = ~new_new_n366__ & ~new_new_n377__;
  assign new_new_n1501__ = ~new_new_n569__ & new_new_n1500__;
  assign new_new_n1502__ = new_new_n379__ & ~new_new_n1501__;
  assign new_new_n1503__ = ~new_new_n379__ & new_new_n1501__;
  assign new_new_n1504__ = ~new_new_n1502__ & ~new_new_n1503__;
  assign new_new_n1505__ = ~new_new_n1499__ & new_new_n1504__;
  assign new_new_n1506__ = new_new_n1498__ & ~new_new_n1505__;
  assign new_new_n1507__ = ~new_new_n1498__ & new_new_n1505__;
  assign new_new_n1508__ = ~new_new_n1506__ & ~new_new_n1507__;
  assign new_new_n1509__ = ~new_new_n1495__ & ~new_new_n1508__;
  assign new_new_n1510__ = new_new_n1495__ & new_new_n1508__;
  assign new_new_n1511__ = ~new_new_n1509__ & ~new_new_n1510__;
  assign new_new_n1512__ = new_new_n560__ & ~new_new_n1511__;
  assign new_new_n1513__ = ~new_new_n381__ & ~new_new_n571__;
  assign new_new_n1514__ = ~new_new_n573__ & new_new_n1513__;
  assign new_new_n1515__ = new_new_n360__ & ~new_new_n1513__;
  assign new_new_n1516__ = ~new_new_n1514__ & ~new_new_n1515__;
  assign new_new_n1517__ = ~new_new_n380__ & new_new_n1382__;
  assign new_new_n1518__ = new_new_n355__ & ~new_new_n1517__;
  assign new_new_n1519__ = ~new_new_n355__ & new_new_n1517__;
  assign new_new_n1520__ = ~new_new_n1518__ & ~new_new_n1519__;
  assign new_new_n1521__ = new_new_n1516__ & new_new_n1520__;
  assign new_new_n1522__ = ~new_new_n1516__ & ~new_new_n1520__;
  assign new_new_n1523__ = ~new_new_n1521__ & ~new_new_n1522__;
  assign new_new_n1524__ = ~new_new_n373__ & ~new_new_n377__;
  assign new_new_n1525__ = ~new_new_n568__ & ~new_new_n1524__;
  assign new_new_n1526__ = new_new_n1498__ & new_new_n1525__;
  assign new_new_n1527__ = ~new_new_n1498__ & ~new_new_n1525__;
  assign new_new_n1528__ = ~new_new_n1526__ & ~new_new_n1527__;
  assign new_new_n1529__ = ~new_new_n1523__ & ~new_new_n1528__;
  assign new_new_n1530__ = new_new_n1523__ & new_new_n1528__;
  assign new_new_n1531__ = ~new_new_n1529__ & ~new_new_n1530__;
  assign new_new_n1532__ = ~new_new_n560__ & ~new_new_n1531__;
  assign new_new_n1533__ = ~new_new_n1512__ & ~new_new_n1532__;
  assign new_new_n1534__ = ~new_new_n387__ & ~new_new_n564__;
  assign new_new_n1535__ = ~new_new_n565__ & ~new_new_n1534__;
  assign new_new_n1536__ = new_new_n404__ & new_new_n1535__;
  assign new_new_n1537__ = ~new_new_n404__ & ~new_new_n1535__;
  assign new_new_n1538__ = ~new_new_n1536__ & ~new_new_n1537__;
  assign new_new_n1539__ = new_new_n393__ & ~new_new_n1538__;
  assign new_new_n1540__ = ~new_new_n393__ & new_new_n1538__;
  assign new_new_n1541__ = ~new_new_n1539__ & ~new_new_n1540__;
  assign new_new_n1542__ = new_new_n397__ & ~new_new_n1541__;
  assign new_new_n1543__ = ~new_new_n397__ & new_new_n1541__;
  assign new_new_n1544__ = ~new_new_n1542__ & ~new_new_n1543__;
  assign new_new_n1545__ = new_new_n1419__ & new_new_n1544__;
  assign new_new_n1546__ = ~new_new_n393__ & ~new_new_n396__;
  assign new_new_n1547__ = ~new_new_n563__ & ~new_new_n1546__;
  assign new_new_n1548__ = ~new_new_n399__ & new_new_n564__;
  assign new_new_n1549__ = ~new_new_n386__ & new_new_n1548__;
  assign new_new_n1550__ = ~new_new_n387__ & ~new_new_n1548__;
  assign new_new_n1551__ = ~new_new_n1549__ & ~new_new_n1550__;
  assign new_new_n1552__ = new_new_n404__ & ~new_new_n1551__;
  assign new_new_n1553__ = ~new_new_n404__ & new_new_n1551__;
  assign new_new_n1554__ = ~new_new_n1552__ & ~new_new_n1553__;
  assign new_new_n1555__ = new_new_n1547__ & ~new_new_n1554__;
  assign new_new_n1556__ = ~new_new_n1547__ & new_new_n1554__;
  assign new_new_n1557__ = ~new_new_n1555__ & ~new_new_n1556__;
  assign new_new_n1558__ = ~new_new_n1419__ & new_new_n1557__;
  assign new_new_n1559__ = ~new_new_n1545__ & ~new_new_n1558__;
  assign new_new_n1560__ = new_new_n388__ & ~new_new_n1559__;
  assign new_new_n1561__ = ~new_new_n388__ & new_new_n1559__;
  assign new_new_n1562__ = ~new_new_n1560__ & ~new_new_n1561__;
  assign new_new_n1563__ = new_new_n1533__ & new_new_n1562__;
  assign new_new_n1564__ = ~new_new_n1533__ & ~new_new_n1562__;
  assign G321 = new_new_n1563__ | new_new_n1564__;
  assign new_new_n1566__ = ~new_new_n595__ & ~new_new_n601__;
  assign new_new_n1567__ = ~new_new_n616__ & new_new_n1566__;
  assign new_new_n1568__ = ~new_new_n597__ & new_new_n1567__;
  assign new_new_n1569__ = new_new_n595__ & ~new_new_n1391__;
  assign new_new_n1570__ = ~new_new_n597__ & ~new_new_n1569__;
  assign new_new_n1571__ = ~new_new_n1567__ & ~new_new_n1570__;
  assign new_new_n1572__ = ~new_new_n1568__ & ~new_new_n1571__;
  assign new_new_n1573__ = ~new_new_n589__ & new_new_n603__;
  assign new_new_n1574__ = new_new_n589__ & ~new_new_n603__;
  assign new_new_n1575__ = ~new_new_n1573__ & ~new_new_n1574__;
  assign new_new_n1576__ = ~new_new_n592__ & ~new_new_n595__;
  assign new_new_n1577__ = ~new_new_n604__ & ~new_new_n1576__;
  assign new_new_n1578__ = new_new_n1393__ & ~new_new_n1577__;
  assign new_new_n1579__ = ~new_new_n1393__ & new_new_n1577__;
  assign new_new_n1580__ = ~new_new_n1578__ & ~new_new_n1579__;
  assign new_new_n1581__ = new_new_n584__ & ~new_new_n1580__;
  assign new_new_n1582__ = ~new_new_n584__ & new_new_n1580__;
  assign new_new_n1583__ = ~new_new_n1581__ & ~new_new_n1582__;
  assign new_new_n1584__ = ~new_new_n1575__ & new_new_n1583__;
  assign new_new_n1585__ = new_new_n1575__ & ~new_new_n1583__;
  assign new_new_n1586__ = ~new_new_n1584__ & ~new_new_n1585__;
  assign new_new_n1587__ = new_new_n1572__ & ~new_new_n1586__;
  assign new_new_n1588__ = ~new_new_n1572__ & new_new_n1586__;
  assign new_new_n1589__ = ~new_new_n1587__ & ~new_new_n1588__;
  assign new_new_n1590__ = new_new_n579__ & new_new_n1589__;
  assign new_new_n1591__ = ~new_new_n595__ & ~new_new_n611__;
  assign new_new_n1592__ = ~new_new_n612__ & ~new_new_n1591__;
  assign new_new_n1593__ = new_new_n603__ & new_new_n1592__;
  assign new_new_n1594__ = ~new_new_n603__ & ~new_new_n1592__;
  assign new_new_n1595__ = ~new_new_n1593__ & ~new_new_n1594__;
  assign new_new_n1596__ = ~new_new_n598__ & ~new_new_n604__;
  assign new_new_n1597__ = ~new_new_n612__ & new_new_n1596__;
  assign new_new_n1598__ = new_new_n584__ & ~new_new_n1597__;
  assign new_new_n1599__ = ~new_new_n584__ & new_new_n1597__;
  assign new_new_n1600__ = ~new_new_n1598__ & ~new_new_n1599__;
  assign new_new_n1601__ = ~new_new_n606__ & new_new_n1391__;
  assign new_new_n1602__ = ~new_new_n1393__ & new_new_n1601__;
  assign new_new_n1603__ = new_new_n588__ & ~new_new_n1601__;
  assign new_new_n1604__ = ~new_new_n1602__ & ~new_new_n1603__;
  assign new_new_n1605__ = new_new_n589__ & ~new_new_n1604__;
  assign new_new_n1606__ = ~new_new_n589__ & new_new_n1604__;
  assign new_new_n1607__ = ~new_new_n1605__ & ~new_new_n1606__;
  assign new_new_n1608__ = new_new_n1600__ & new_new_n1607__;
  assign new_new_n1609__ = ~new_new_n1600__ & ~new_new_n1607__;
  assign new_new_n1610__ = ~new_new_n1608__ & ~new_new_n1609__;
  assign new_new_n1611__ = ~new_new_n1595__ & ~new_new_n1610__;
  assign new_new_n1612__ = new_new_n1595__ & new_new_n1610__;
  assign new_new_n1613__ = ~new_new_n1611__ & ~new_new_n1612__;
  assign new_new_n1614__ = ~new_new_n579__ & new_new_n1613__;
  assign new_new_n1615__ = ~new_new_n1590__ & ~new_new_n1614__;
  assign new_new_n1616__ = ~new_new_n343__ & new_new_n1446__;
  assign new_new_n1617__ = ~new_new_n344__ & new_new_n624__;
  assign new_new_n1618__ = new_new_n346__ & new_new_n623__;
  assign new_new_n1619__ = ~new_new_n1617__ & ~new_new_n1618__;
  assign new_new_n1620__ = ~new_new_n1446__ & new_new_n1619__;
  assign new_new_n1621__ = ~new_new_n1616__ & ~new_new_n1620__;
  assign new_new_n1622__ = new_new_n1615__ & ~new_new_n1621__;
  assign new_new_n1623__ = ~new_new_n1615__ & new_new_n1621__;
  assign G338 = ~new_new_n1622__ & ~new_new_n1623__;
  assign new_new_n1625__ = ~new_new_n490__ & new_new_n507__;
  assign new_new_n1626__ = new_new_n490__ & ~new_new_n507__;
  assign new_new_n1627__ = ~new_new_n1625__ & ~new_new_n1626__;
  assign new_new_n1628__ = ~new_new_n498__ & ~new_new_n505__;
  assign new_new_n1629__ = ~new_new_n520__ & new_new_n1628__;
  assign new_new_n1630__ = ~new_new_n500__ & new_new_n1629__;
  assign new_new_n1631__ = new_new_n498__ & ~new_new_n1449__;
  assign new_new_n1632__ = ~new_new_n500__ & ~new_new_n1631__;
  assign new_new_n1633__ = ~new_new_n1629__ & ~new_new_n1632__;
  assign new_new_n1634__ = ~new_new_n1630__ & ~new_new_n1633__;
  assign new_new_n1635__ = ~new_new_n494__ & ~new_new_n498__;
  assign new_new_n1636__ = ~new_new_n508__ & ~new_new_n1635__;
  assign new_new_n1637__ = new_new_n1451__ & ~new_new_n1636__;
  assign new_new_n1638__ = ~new_new_n1451__ & new_new_n1636__;
  assign new_new_n1639__ = ~new_new_n1637__ & ~new_new_n1638__;
  assign new_new_n1640__ = new_new_n484__ & ~new_new_n1639__;
  assign new_new_n1641__ = ~new_new_n484__ & new_new_n1639__;
  assign new_new_n1642__ = ~new_new_n1640__ & ~new_new_n1641__;
  assign new_new_n1643__ = new_new_n1634__ & new_new_n1642__;
  assign new_new_n1644__ = ~new_new_n1634__ & ~new_new_n1642__;
  assign new_new_n1645__ = ~new_new_n1643__ & ~new_new_n1644__;
  assign new_new_n1646__ = ~new_new_n1627__ & new_new_n1645__;
  assign new_new_n1647__ = new_new_n1627__ & ~new_new_n1645__;
  assign new_new_n1648__ = ~new_new_n1646__ & ~new_new_n1647__;
  assign new_new_n1649__ = new_new_n478__ & ~new_new_n1648__;
  assign new_new_n1650__ = ~new_new_n510__ & new_new_n1449__;
  assign new_new_n1651__ = ~new_new_n1451__ & new_new_n1650__;
  assign new_new_n1652__ = new_new_n489__ & ~new_new_n1650__;
  assign new_new_n1653__ = ~new_new_n1651__ & ~new_new_n1652__;
  assign new_new_n1654__ = ~new_new_n501__ & ~new_new_n508__;
  assign new_new_n1655__ = ~new_new_n516__ & new_new_n1654__;
  assign new_new_n1656__ = new_new_n484__ & ~new_new_n1655__;
  assign new_new_n1657__ = ~new_new_n484__ & new_new_n1655__;
  assign new_new_n1658__ = ~new_new_n1656__ & ~new_new_n1657__;
  assign new_new_n1659__ = new_new_n1653__ & new_new_n1658__;
  assign new_new_n1660__ = ~new_new_n1653__ & ~new_new_n1658__;
  assign new_new_n1661__ = ~new_new_n1659__ & ~new_new_n1660__;
  assign new_new_n1662__ = ~new_new_n498__ & ~new_new_n515__;
  assign new_new_n1663__ = ~new_new_n516__ & ~new_new_n1662__;
  assign new_new_n1664__ = new_new_n1627__ & new_new_n1663__;
  assign new_new_n1665__ = ~new_new_n1627__ & ~new_new_n1663__;
  assign new_new_n1666__ = ~new_new_n1664__ & ~new_new_n1665__;
  assign new_new_n1667__ = ~new_new_n1661__ & ~new_new_n1666__;
  assign new_new_n1668__ = new_new_n1661__ & new_new_n1666__;
  assign new_new_n1669__ = ~new_new_n478__ & ~new_new_n1667__;
  assign new_new_n1670__ = ~new_new_n1668__ & new_new_n1669__;
  assign new_new_n1671__ = ~new_new_n1649__ & ~new_new_n1670__;
  assign new_new_n1672__ = ~new_new_n549__ & new_new_n555__;
  assign new_new_n1673__ = ~new_new_n556__ & ~new_new_n1672__;
  assign new_new_n1674__ = new_new_n544__ & ~new_new_n1673__;
  assign new_new_n1675__ = ~new_new_n544__ & new_new_n1673__;
  assign new_new_n1676__ = ~new_new_n1674__ & ~new_new_n1675__;
  assign new_new_n1677__ = ~new_new_n536__ & new_new_n1676__;
  assign new_new_n1678__ = new_new_n536__ & ~new_new_n1676__;
  assign new_new_n1679__ = ~new_new_n1677__ & ~new_new_n1678__;
  assign new_new_n1680__ = new_new_n531__ & new_new_n1679__;
  assign new_new_n1681__ = ~new_new_n531__ & ~new_new_n1679__;
  assign new_new_n1682__ = ~new_new_n1680__ & ~new_new_n1681__;
  assign new_new_n1683__ = new_new_n525__ & new_new_n1682__;
  assign new_new_n1684__ = ~new_new_n531__ & ~new_new_n535__;
  assign new_new_n1685__ = ~new_new_n554__ & ~new_new_n1684__;
  assign new_new_n1686__ = ~new_new_n538__ & new_new_n555__;
  assign new_new_n1687__ = ~new_new_n549__ & new_new_n1686__;
  assign new_new_n1688__ = ~new_new_n548__ & ~new_new_n1686__;
  assign new_new_n1689__ = ~new_new_n1687__ & ~new_new_n1688__;
  assign new_new_n1690__ = ~new_new_n544__ & ~new_new_n1689__;
  assign new_new_n1691__ = new_new_n544__ & new_new_n1689__;
  assign new_new_n1692__ = ~new_new_n1690__ & ~new_new_n1691__;
  assign new_new_n1693__ = new_new_n1685__ & new_new_n1692__;
  assign new_new_n1694__ = ~new_new_n1685__ & ~new_new_n1692__;
  assign new_new_n1695__ = ~new_new_n1693__ & ~new_new_n1694__;
  assign new_new_n1696__ = ~new_new_n525__ & new_new_n1695__;
  assign new_new_n1697__ = ~new_new_n1683__ & ~new_new_n1696__;
  assign new_new_n1698__ = new_new_n550__ & ~new_new_n1697__;
  assign new_new_n1699__ = ~new_new_n550__ & new_new_n1697__;
  assign new_new_n1700__ = ~new_new_n1698__ & ~new_new_n1699__;
  assign new_new_n1701__ = new_new_n1671__ & new_new_n1700__;
  assign new_new_n1702__ = ~new_new_n1671__ & ~new_new_n1700__;
  assign G370 = ~new_new_n1701__ & ~new_new_n1702__;
  assign new_new_n1704__ = new_new_n435__ & new_new_n438__;
  assign new_new_n1705__ = ~new_new_n414__ & new_new_n1704__;
  assign new_new_n1706__ = ~new_new_n432__ & ~new_new_n1705__;
  assign new_new_n1707__ = new_new_n971__ & ~new_new_n1706__;
  assign new_new_n1708__ = ~new_new_n971__ & new_new_n1706__;
  assign new_new_n1709__ = ~new_new_n1707__ & ~new_new_n1708__;
  assign new_new_n1710__ = ~new_new_n338__ & new_new_n1704__;
  assign new_new_n1711__ = ~new_new_n430__ & ~new_new_n1710__;
  assign new_new_n1712__ = new_new_n334__ & ~new_new_n338__;
  assign new_new_n1713__ = ~new_new_n1711__ & new_new_n1712__;
  assign new_new_n1714__ = new_new_n1711__ & ~new_new_n1712__;
  assign new_new_n1715__ = ~new_new_n1713__ & ~new_new_n1714__;
  assign new_new_n1716__ = new_new_n339__ & ~new_new_n424__;
  assign new_new_n1717__ = new_new_n982__ & ~new_new_n1716__;
  assign new_new_n1718__ = new_new_n425__ & ~new_new_n1717__;
  assign new_new_n1719__ = ~new_new_n425__ & new_new_n1717__;
  assign new_new_n1720__ = ~new_new_n1718__ & ~new_new_n1719__;
  assign new_new_n1721__ = new_new_n1715__ & ~new_new_n1720__;
  assign new_new_n1722__ = ~new_new_n1715__ & new_new_n1720__;
  assign new_new_n1723__ = ~new_new_n1721__ & ~new_new_n1722__;
  assign new_new_n1724__ = new_new_n1709__ & ~new_new_n1723__;
  assign new_new_n1725__ = ~new_new_n1709__ & new_new_n1723__;
  assign new_new_n1726__ = ~new_new_n1724__ & ~new_new_n1725__;
  assign new_new_n1727__ = G4526 & ~new_new_n1726__;
  assign new_new_n1728__ = new_new_n432__ & ~new_new_n971__;
  assign new_new_n1729__ = ~new_new_n432__ & new_new_n971__;
  assign new_new_n1730__ = ~new_new_n1728__ & ~new_new_n1729__;
  assign new_new_n1731__ = new_new_n334__ & ~new_new_n430__;
  assign new_new_n1732__ = ~new_new_n334__ & ~new_new_n419__;
  assign new_new_n1733__ = ~new_new_n428__ & new_new_n1732__;
  assign new_new_n1734__ = new_new_n339__ & ~new_new_n1733__;
  assign new_new_n1735__ = ~new_new_n339__ & new_new_n1733__;
  assign new_new_n1736__ = ~new_new_n1734__ & ~new_new_n1735__;
  assign new_new_n1737__ = ~new_new_n1731__ & new_new_n1736__;
  assign new_new_n1738__ = ~new_new_n334__ & ~new_new_n424__;
  assign new_new_n1739__ = ~new_new_n423__ & ~new_new_n1738__;
  assign new_new_n1740__ = new_new_n1737__ & ~new_new_n1739__;
  assign new_new_n1741__ = ~new_new_n1737__ & new_new_n1739__;
  assign new_new_n1742__ = ~new_new_n1740__ & ~new_new_n1741__;
  assign new_new_n1743__ = new_new_n1730__ & ~new_new_n1742__;
  assign new_new_n1744__ = ~new_new_n1730__ & new_new_n1742__;
  assign new_new_n1745__ = ~new_new_n1743__ & ~new_new_n1744__;
  assign new_new_n1746__ = ~G4526 & ~new_new_n1745__;
  assign new_new_n1747__ = ~new_new_n1727__ & ~new_new_n1746__;
  assign new_new_n1748__ = ~new_new_n435__ & ~new_new_n436__;
  assign new_new_n1749__ = ~new_new_n437__ & ~new_new_n1748__;
  assign new_new_n1750__ = new_new_n461__ & new_new_n473__;
  assign new_new_n1751__ = new_new_n460__ & ~new_new_n473__;
  assign new_new_n1752__ = ~new_new_n1750__ & ~new_new_n1751__;
  assign new_new_n1753__ = new_new_n468__ & ~new_new_n1752__;
  assign new_new_n1754__ = ~new_new_n468__ & new_new_n1752__;
  assign new_new_n1755__ = ~new_new_n1753__ & ~new_new_n1754__;
  assign new_new_n1756__ = ~new_new_n449__ & new_new_n454__;
  assign new_new_n1757__ = new_new_n449__ & ~new_new_n454__;
  assign new_new_n1758__ = ~new_new_n1756__ & ~new_new_n1757__;
  assign new_new_n1759__ = ~new_new_n1755__ & ~new_new_n1758__;
  assign new_new_n1760__ = new_new_n1755__ & new_new_n1758__;
  assign new_new_n1761__ = ~new_new_n1759__ & ~new_new_n1760__;
  assign new_new_n1762__ = new_new_n443__ & ~new_new_n1761__;
  assign new_new_n1763__ = ~new_new_n449__ & ~new_new_n453__;
  assign new_new_n1764__ = ~new_new_n472__ & ~new_new_n1763__;
  assign new_new_n1765__ = ~new_new_n462__ & ~new_new_n468__;
  assign new_new_n1766__ = ~new_new_n469__ & ~new_new_n1765__;
  assign new_new_n1767__ = new_new_n1764__ & ~new_new_n1766__;
  assign new_new_n1768__ = ~new_new_n1764__ & new_new_n1766__;
  assign new_new_n1769__ = ~new_new_n1767__ & ~new_new_n1768__;
  assign new_new_n1770__ = ~new_new_n447__ & ~new_new_n1757__;
  assign new_new_n1771__ = ~new_new_n460__ & new_new_n1770__;
  assign new_new_n1772__ = ~new_new_n461__ & ~new_new_n1770__;
  assign new_new_n1773__ = ~new_new_n1771__ & ~new_new_n1772__;
  assign new_new_n1774__ = ~new_new_n1769__ & ~new_new_n1773__;
  assign new_new_n1775__ = new_new_n1769__ & new_new_n1773__;
  assign new_new_n1776__ = ~new_new_n1774__ & ~new_new_n1775__;
  assign new_new_n1777__ = ~new_new_n443__ & new_new_n1776__;
  assign new_new_n1778__ = ~new_new_n1762__ & ~new_new_n1777__;
  assign new_new_n1779__ = new_new_n1749__ & ~new_new_n1778__;
  assign new_new_n1780__ = ~new_new_n1749__ & new_new_n1778__;
  assign new_new_n1781__ = ~new_new_n1779__ & ~new_new_n1780__;
  assign new_new_n1782__ = new_new_n1747__ & new_new_n1781__;
  assign new_new_n1783__ = ~new_new_n1747__ & ~new_new_n1781__;
  assign G399 = ~new_new_n1782__ & ~new_new_n1783__;
  assign G279 = ~G15;
  assign G339 = \IN-G339 ;
  // assign G2 = G1;
  // assign G3 = G1;
  // assign G450 = G1459;
  // assign G448 = G1469;
  // assign G444 = G1480;
  // assign G442 = G1486;
  // assign G440 = G1492;
  // assign G438 = G1496;
  // assign G496 = G2208;
  // assign G494 = G2218;
  // assign G492 = G2224;
  // assign G490 = G2230;
  // assign G488 = G2236;
  // assign G486 = G2239;
  // assign G484 = G2247;
  // assign G482 = G2253;
  // assign G480 = G2256;
  // assign G560 = G3698;
  // assign G542 = G3701;
  // assign G558 = G3705;
  // assign G556 = G3711;
  // assign G554 = G3717;
  // assign G552 = G3723;
  // assign G550 = G3729;
  // assign G548 = G3737;
  // assign G546 = G3743;
  // assign G544 = G3749;
  // assign G540 = G4393;
  // assign G538 = G4400;
  // assign G536 = G4405;
  // assign G534 = G4410;
  // assign G532 = G4415;
  // assign G530 = G4420;
  // assign G528 = G4427;
  // assign G526 = G4432;
  // assign G524 = G4437;
  // assign G436 = G1462;
  // assign G478 = G2211;
  // assign G522 = G4394;
  // assign G432 = G1;
  // assign G446 = G106;
  // assign G286 = G279;
  // assign G289 = G284;
  // assign G341 = G279;
  // assign G281 = G292;
  // assign G453 = G1;
  // assign G264 = G258;
  // assign G270 = G246;
  // assign G249 = G258;
  // assign G276 = G246;
  // assign G273 = G246;
  // assign G469 = G422;
  // assign G471 = G419;
endmodule


