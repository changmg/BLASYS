module max_34_1(pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 , po0 , po1 , po2 , po3 , po4 );
  input pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 ;
  output po0 , po1 , po2 , po3 , po4 ;
  wire new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36, new_n37, new_n38, new_n39;
  assign new_n12 = ~pi01 & pi03 ;
  assign new_n13 = ~pi00 & pi02 ;
  assign new_n14 = ~pi09 & ~new_n13 ;
  assign new_n15 = pi01 & ~pi03 ;
  assign new_n16 = pi00 & ~pi02 ;
  assign new_n17 = ~new_n15 & ~new_n16 ;
  assign new_n18 = ~new_n14 & new_n17 ;
  assign new_n19 = ~new_n12 & ~new_n18 ;
  assign new_n20 = pi00 & pi04 ;
  assign new_n21 = pi02 & ~pi04 ;
  assign new_n22 = ~new_n20 & ~new_n21 ;
  assign new_n23 = pi05 & ~new_n22 ;
  assign new_n24 = pi01 & pi04 ;
  assign new_n25 = pi03 & ~pi04 ;
  assign new_n26 = ~new_n24 & ~new_n25 ;
  assign new_n27 = ~pi06 & new_n26 ;
  assign new_n28 = ~pi05 & new_n22 ;
  assign new_n29 = ~new_n27 & ~new_n28 ;
  assign new_n30 = ~pi10 & new_n29 ;
  assign new_n31 = pi06 & ~new_n26 ;
  assign new_n32 = ~pi07 & ~new_n31 ;
  assign new_n33 = ~new_n30 & new_n32 ;
  assign new_n34 = pi08 & ~new_n22 ;
  assign new_n35 = ~pi05 & ~pi08 ;
  assign new_n36 = ~new_n34 & ~new_n35 ;
  assign new_n37 = pi08 & ~new_n26 ;
  assign new_n38 = ~pi06 & ~pi08 ;
  assign new_n39 = ~new_n37 & ~new_n38 ;
  assign po0 = new_n19 ;
  assign po1 = new_n23 ;
  assign po2 = new_n33 ;
  assign po3 = new_n36 ;
  assign po4 = new_n39 ;
endmodule
