module max(pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020
, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041
, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062
, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083
, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104
, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125
, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146
, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167
, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188
, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209
, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230
, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251
, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272
, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293
, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314
, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335
, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356
, pi357, pi358, pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377
, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398
, pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419
, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440
, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459, pi460, pi461
, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479, pi480, pi481, pi482
, pi483, pi484, pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503
, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511, po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012
, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033
, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054
, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075
, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096
, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117
, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129);
  input pi000;
  input pi001;
  input pi002;
  input pi003;
  input pi004;
  input pi005;
  input pi006;
  input pi007;
  input pi008;
  input pi009;
  input pi010;
  input pi011;
  input pi012;
  input pi013;
  input pi014;
  input pi015;
  input pi016;
  input pi017;
  input pi018;
  input pi019;
  input pi020;
  input pi021;
  input pi022;
  input pi023;
  input pi024;
  input pi025;
  input pi026;
  input pi027;
  input pi028;
  input pi029;
  input pi030;
  input pi031;
  input pi032;
  input pi033;
  input pi034;
  input pi035;
  input pi036;
  input pi037;
  input pi038;
  input pi039;
  input pi040;
  input pi041;
  input pi042;
  input pi043;
  input pi044;
  input pi045;
  input pi046;
  input pi047;
  input pi048;
  input pi049;
  input pi050;
  input pi051;
  input pi052;
  input pi053;
  input pi054;
  input pi055;
  input pi056;
  input pi057;
  input pi058;
  input pi059;
  input pi060;
  input pi061;
  input pi062;
  input pi063;
  input pi064;
  input pi065;
  input pi066;
  input pi067;
  input pi068;
  input pi069;
  input pi070;
  input pi071;
  input pi072;
  input pi073;
  input pi074;
  input pi075;
  input pi076;
  input pi077;
  input pi078;
  input pi079;
  input pi080;
  input pi081;
  input pi082;
  input pi083;
  input pi084;
  input pi085;
  input pi086;
  input pi087;
  input pi088;
  input pi089;
  input pi090;
  input pi091;
  input pi092;
  input pi093;
  input pi094;
  input pi095;
  input pi096;
  input pi097;
  input pi098;
  input pi099;
  input pi100;
  input pi101;
  input pi102;
  input pi103;
  input pi104;
  input pi105;
  input pi106;
  input pi107;
  input pi108;
  input pi109;
  input pi110;
  input pi111;
  input pi112;
  input pi113;
  input pi114;
  input pi115;
  input pi116;
  input pi117;
  input pi118;
  input pi119;
  input pi120;
  input pi121;
  input pi122;
  input pi123;
  input pi124;
  input pi125;
  input pi126;
  input pi127;
  input pi128;
  input pi129;
  input pi130;
  input pi131;
  input pi132;
  input pi133;
  input pi134;
  input pi135;
  input pi136;
  input pi137;
  input pi138;
  input pi139;
  input pi140;
  input pi141;
  input pi142;
  input pi143;
  input pi144;
  input pi145;
  input pi146;
  input pi147;
  input pi148;
  input pi149;
  input pi150;
  input pi151;
  input pi152;
  input pi153;
  input pi154;
  input pi155;
  input pi156;
  input pi157;
  input pi158;
  input pi159;
  input pi160;
  input pi161;
  input pi162;
  input pi163;
  input pi164;
  input pi165;
  input pi166;
  input pi167;
  input pi168;
  input pi169;
  input pi170;
  input pi171;
  input pi172;
  input pi173;
  input pi174;
  input pi175;
  input pi176;
  input pi177;
  input pi178;
  input pi179;
  input pi180;
  input pi181;
  input pi182;
  input pi183;
  input pi184;
  input pi185;
  input pi186;
  input pi187;
  input pi188;
  input pi189;
  input pi190;
  input pi191;
  input pi192;
  input pi193;
  input pi194;
  input pi195;
  input pi196;
  input pi197;
  input pi198;
  input pi199;
  input pi200;
  input pi201;
  input pi202;
  input pi203;
  input pi204;
  input pi205;
  input pi206;
  input pi207;
  input pi208;
  input pi209;
  input pi210;
  input pi211;
  input pi212;
  input pi213;
  input pi214;
  input pi215;
  input pi216;
  input pi217;
  input pi218;
  input pi219;
  input pi220;
  input pi221;
  input pi222;
  input pi223;
  input pi224;
  input pi225;
  input pi226;
  input pi227;
  input pi228;
  input pi229;
  input pi230;
  input pi231;
  input pi232;
  input pi233;
  input pi234;
  input pi235;
  input pi236;
  input pi237;
  input pi238;
  input pi239;
  input pi240;
  input pi241;
  input pi242;
  input pi243;
  input pi244;
  input pi245;
  input pi246;
  input pi247;
  input pi248;
  input pi249;
  input pi250;
  input pi251;
  input pi252;
  input pi253;
  input pi254;
  input pi255;
  input pi256;
  input pi257;
  input pi258;
  input pi259;
  input pi260;
  input pi261;
  input pi262;
  input pi263;
  input pi264;
  input pi265;
  input pi266;
  input pi267;
  input pi268;
  input pi269;
  input pi270;
  input pi271;
  input pi272;
  input pi273;
  input pi274;
  input pi275;
  input pi276;
  input pi277;
  input pi278;
  input pi279;
  input pi280;
  input pi281;
  input pi282;
  input pi283;
  input pi284;
  input pi285;
  input pi286;
  input pi287;
  input pi288;
  input pi289;
  input pi290;
  input pi291;
  input pi292;
  input pi293;
  input pi294;
  input pi295;
  input pi296;
  input pi297;
  input pi298;
  input pi299;
  input pi300;
  input pi301;
  input pi302;
  input pi303;
  input pi304;
  input pi305;
  input pi306;
  input pi307;
  input pi308;
  input pi309;
  input pi310;
  input pi311;
  input pi312;
  input pi313;
  input pi314;
  input pi315;
  input pi316;
  input pi317;
  input pi318;
  input pi319;
  input pi320;
  input pi321;
  input pi322;
  input pi323;
  input pi324;
  input pi325;
  input pi326;
  input pi327;
  input pi328;
  input pi329;
  input pi330;
  input pi331;
  input pi332;
  input pi333;
  input pi334;
  input pi335;
  input pi336;
  input pi337;
  input pi338;
  input pi339;
  input pi340;
  input pi341;
  input pi342;
  input pi343;
  input pi344;
  input pi345;
  input pi346;
  input pi347;
  input pi348;
  input pi349;
  input pi350;
  input pi351;
  input pi352;
  input pi353;
  input pi354;
  input pi355;
  input pi356;
  input pi357;
  input pi358;
  input pi359;
  input pi360;
  input pi361;
  input pi362;
  input pi363;
  input pi364;
  input pi365;
  input pi366;
  input pi367;
  input pi368;
  input pi369;
  input pi370;
  input pi371;
  input pi372;
  input pi373;
  input pi374;
  input pi375;
  input pi376;
  input pi377;
  input pi378;
  input pi379;
  input pi380;
  input pi381;
  input pi382;
  input pi383;
  input pi384;
  input pi385;
  input pi386;
  input pi387;
  input pi388;
  input pi389;
  input pi390;
  input pi391;
  input pi392;
  input pi393;
  input pi394;
  input pi395;
  input pi396;
  input pi397;
  input pi398;
  input pi399;
  input pi400;
  input pi401;
  input pi402;
  input pi403;
  input pi404;
  input pi405;
  input pi406;
  input pi407;
  input pi408;
  input pi409;
  input pi410;
  input pi411;
  input pi412;
  input pi413;
  input pi414;
  input pi415;
  input pi416;
  input pi417;
  input pi418;
  input pi419;
  input pi420;
  input pi421;
  input pi422;
  input pi423;
  input pi424;
  input pi425;
  input pi426;
  input pi427;
  input pi428;
  input pi429;
  input pi430;
  input pi431;
  input pi432;
  input pi433;
  input pi434;
  input pi435;
  input pi436;
  input pi437;
  input pi438;
  input pi439;
  input pi440;
  input pi441;
  input pi442;
  input pi443;
  input pi444;
  input pi445;
  input pi446;
  input pi447;
  input pi448;
  input pi449;
  input pi450;
  input pi451;
  input pi452;
  input pi453;
  input pi454;
  input pi455;
  input pi456;
  input pi457;
  input pi458;
  input pi459;
  input pi460;
  input pi461;
  input pi462;
  input pi463;
  input pi464;
  input pi465;
  input pi466;
  input pi467;
  input pi468;
  input pi469;
  input pi470;
  input pi471;
  input pi472;
  input pi473;
  input pi474;
  input pi475;
  input pi476;
  input pi477;
  input pi478;
  input pi479;
  input pi480;
  input pi481;
  input pi482;
  input pi483;
  input pi484;
  input pi485;
  input pi486;
  input pi487;
  input pi488;
  input pi489;
  input pi490;
  input pi491;
  input pi492;
  input pi493;
  input pi494;
  input pi495;
  input pi496;
  input pi497;
  input pi498;
  input pi499;
  input pi500;
  input pi501;
  input pi502;
  input pi503;
  input pi504;
  input pi505;
  input pi506;
  input pi507;
  input pi508;
  input pi509;
  input pi510;
  input pi511;
  output po000;
  output po001;
  output po002;
  output po003;
  output po004;
  output po005;
  output po006;
  output po007;
  output po008;
  output po009;
  output po010;
  output po011;
  output po012;
  output po013;
  output po014;
  output po015;
  output po016;
  output po017;
  output po018;
  output po019;
  output po020;
  output po021;
  output po022;
  output po023;
  output po024;
  output po025;
  output po026;
  output po027;
  output po028;
  output po029;
  output po030;
  output po031;
  output po032;
  output po033;
  output po034;
  output po035;
  output po036;
  output po037;
  output po038;
  output po039;
  output po040;
  output po041;
  output po042;
  output po043;
  output po044;
  output po045;
  output po046;
  output po047;
  output po048;
  output po049;
  output po050;
  output po051;
  output po052;
  output po053;
  output po054;
  output po055;
  output po056;
  output po057;
  output po058;
  output po059;
  output po060;
  output po061;
  output po062;
  output po063;
  output po064;
  output po065;
  output po066;
  output po067;
  output po068;
  output po069;
  output po070;
  output po071;
  output po072;
  output po073;
  output po074;
  output po075;
  output po076;
  output po077;
  output po078;
  output po079;
  output po080;
  output po081;
  output po082;
  output po083;
  output po084;
  output po085;
  output po086;
  output po087;
  output po088;
  output po089;
  output po090;
  output po091;
  output po092;
  output po093;
  output po094;
  output po095;
  output po096;
  output po097;
  output po098;
  output po099;
  output po100;
  output po101;
  output po102;
  output po103;
  output po104;
  output po105;
  output po106;
  output po107;
  output po108;
  output po109;
  output po110;
  output po111;
  output po112;
  output po113;
  output po114;
  output po115;
  output po116;
  output po117;
  output po118;
  output po119;
  output po120;
  output po121;
  output po122;
  output po123;
  output po124;
  output po125;
  output po126;
  output po127;
  output po128;
  output po129;
  top U0 ( .pi000( pi000 ) , .pi001( pi001 ) , .pi002( pi002 ) , .pi003( pi003 ) , .pi004( pi004 ) , .pi005( pi005 ) , .pi006( pi006 ) , .pi007( pi007 ) , .pi008( pi008 ) , .pi009( pi009 ) , .pi010( pi010 ) , .pi011( pi011 ) , .pi012( pi012 ) , .pi013( pi013 ) , .pi014( pi014 ) , .pi015( pi015 ) , .pi016( pi016 ) , .pi017( pi017 ) , .pi018( pi018 ) , .pi019( pi019 ) , .pi020( pi020 ) , .pi021( pi021 ) , .pi022( pi022 ) , .pi023( pi023 ) , .pi024( pi024 ) , .pi025( pi025 ) , .pi026( pi026 ) , .pi027( pi027 ) , .pi028( pi028 ) , .pi029( pi029 ) , .pi030( pi030 ) , .pi031( pi031 ) , .pi032( pi032 ) , .pi033( pi033 ) , .pi034( pi034 ) , .pi035( pi035 ) , .pi036( pi036 ) , .pi037( pi037 ) , .pi038( pi038 ) , .pi039( pi039 ) , .pi040( pi040 ) , .pi041( pi041 ) , .pi042( pi042 ) , .pi043( pi043 ) , .pi044( pi044 ) , .pi045( pi045 ) , .pi046( pi046 ) , .pi047( pi047 ) , .pi048( pi048 ) , .pi049( pi049 ) , .pi050( pi050 ) , .pi051( pi051 ) , .pi052( pi052 ) , .pi053( pi053 ) , .pi054( pi054 ) , .pi055( pi055 ) , .pi056( pi056 ) , .pi057( pi057 ) , .pi058( pi058 ) , .pi059( pi059 ) , .pi060( pi060 ) , .pi061( pi061 ) , .pi062( pi062 ) , .pi063( pi063 ) , .pi064( pi064 ) , .pi065( pi065 ) , .pi066( pi066 ) , .pi067( pi067 ) , .pi068( pi068 ) , .pi069( pi069 ) , .pi070( pi070 ) , .pi071( pi071 ) , .pi072( pi072 ) , .pi073( pi073 ) , .pi074( pi074 ) , .pi075( pi075 ) , .pi076( pi076 ) , .pi077( pi077 ) , .pi078( pi078 ) , .pi079( pi079 ) , .pi080( pi080 ) , .pi081( pi081 ) , .pi082( pi082 ) , .pi083( pi083 ) , .pi084( pi084 ) , .pi085( pi085 ) , .pi086( pi086 ) , .pi087( pi087 ) , .pi088( pi088 ) , .pi089( pi089 ) , .pi090( pi090 ) , .pi091( pi091 ) , .pi092( pi092 ) , .pi093( pi093 ) , .pi094( pi094 ) , .pi095( pi095 ) , .pi096( pi096 ) , .pi097( pi097 ) , .pi098( pi098 ) , .pi099( pi099 ) , .pi100( pi100 ) , .pi101( pi101 ) , .pi102( pi102 ) , .pi103( pi103 ) , .pi104( pi104 ) , .pi105( pi105 ) , .pi106( pi106 ) , .pi107( pi107 ) , .pi108( pi108 ) , .pi109( pi109 ) , .pi110( pi110 ) , .pi111( pi111 ) , .pi112( pi112 ) , .pi113( pi113 ) , .pi114( pi114 ) , .pi115( pi115 ) , .pi116( pi116 ) , .pi117( pi117 ) , .pi118( pi118 ) , .pi119( pi119 ) , .pi120( pi120 ) , .pi121( pi121 ) , .pi122( pi122 ) , .pi123( pi123 ) , .pi124( pi124 ) , .pi125( pi125 ) , .pi126( pi126 ) , .pi127( pi127 ) , .pi128( pi128 ) , .pi129( pi129 ) , .pi130( pi130 ) , .pi131( pi131 ) , .pi132( pi132 ) , .pi133( pi133 ) , .pi134( pi134 ) , .pi135( pi135 ) , .pi136( pi136 ) , .pi137( pi137 ) , .pi138( pi138 ) , .pi139( pi139 ) , .pi140( pi140 ) , .pi141( pi141 ) , .pi142( pi142 ) , .pi143( pi143 ) , .pi144( pi144 ) , .pi145( pi145 ) , .pi146( pi146 ) , .pi147( pi147 ) , .pi148( pi148 ) , .pi149( pi149 ) , .pi150( pi150 ) , .pi151( pi151 ) , .pi152( pi152 ) , .pi153( pi153 ) , .pi154( pi154 ) , .pi155( pi155 ) , .pi156( pi156 ) , .pi157( pi157 ) , .pi158( pi158 ) , .pi159( pi159 ) , .pi160( pi160 ) , .pi161( pi161 ) , .pi162( pi162 ) , .pi163( pi163 ) , .pi164( pi164 ) , .pi165( pi165 ) , .pi166( pi166 ) , .pi167( pi167 ) , .pi168( pi168 ) , .pi169( pi169 ) , .pi170( pi170 ) , .pi171( pi171 ) , .pi172( pi172 ) , .pi173( pi173 ) , .pi174( pi174 ) , .pi175( pi175 ) , .pi176( pi176 ) , .pi177( pi177 ) , .pi178( pi178 ) , .pi179( pi179 ) , .pi180( pi180 ) , .pi181( pi181 ) , .pi182( pi182 ) , .pi183( pi183 ) , .pi184( pi184 ) , .pi185( pi185 ) , .pi186( pi186 ) , .pi187( pi187 ) , .pi188( pi188 ) , .pi189( pi189 ) , .pi190( pi190 ) , .pi191( pi191 ) , .pi192( pi192 ) , .pi193( pi193 ) , .pi194( pi194 ) , .pi195( pi195 ) , .pi196( pi196 ) , .pi197( pi197 ) , .pi198( pi198 ) , .pi199( pi199 ) , .pi200( pi200 ) , .pi201( pi201 ) , .pi202( pi202 ) , .pi203( pi203 ) , .pi204( pi204 ) , .pi205( pi205 ) , .pi206( pi206 ) , .pi207( pi207 ) , .pi208( pi208 ) , .pi209( pi209 ) , .pi210( pi210 ) , .pi211( pi211 ) , .pi212( pi212 ) , .pi213( pi213 ) , .pi214( pi214 ) , .pi215( pi215 ) , .pi216( pi216 ) , .pi217( pi217 ) , .pi218( pi218 ) , .pi219( pi219 ) , .pi220( pi220 ) , .pi221( pi221 ) , .pi222( pi222 ) , .pi223( pi223 ) , .pi224( pi224 ) , .pi225( pi225 ) , .pi226( pi226 ) , .pi227( pi227 ) , .pi228( pi228 ) , .pi229( pi229 ) , .pi230( pi230 ) , .pi231( pi231 ) , .pi232( pi232 ) , .pi233( pi233 ) , .pi234( pi234 ) , .pi235( pi235 ) , .pi236( pi236 ) , .pi237( pi237 ) , .pi238( pi238 ) , .pi239( pi239 ) , .pi240( pi240 ) , .pi241( pi241 ) , .pi242( pi242 ) , .pi243( pi243 ) , .pi244( pi244 ) , .pi245( pi245 ) , .pi246( pi246 ) , .pi247( pi247 ) , .pi248( pi248 ) , .pi249( pi249 ) , .pi250( pi250 ) , .pi251( pi251 ) , .pi252( pi252 ) , .pi253( pi253 ) , .pi254( pi254 ) , .pi255( pi255 ) , .pi256( pi256 ) , .pi257( pi257 ) , .pi258( pi258 ) , .pi259( pi259 ) , .pi260( pi260 ) , .pi261( pi261 ) , .pi262( pi262 ) , .pi263( pi263 ) , .pi264( pi264 ) , .pi265( pi265 ) , .pi266( pi266 ) , .pi267( pi267 ) , .pi268( pi268 ) , .pi269( pi269 ) , .pi270( pi270 ) , .pi271( pi271 ) , .pi272( pi272 ) , .pi273( pi273 ) , .pi274( pi274 ) , .pi275( pi275 ) , .pi276( pi276 ) , .pi277( pi277 ) , .pi278( pi278 ) , .pi279( pi279 ) , .pi280( pi280 ) , .pi281( pi281 ) , .pi282( pi282 ) , .pi283( pi283 ) , .pi284( pi284 ) , .pi285( pi285 ) , .pi286( pi286 ) , .pi287( pi287 ) , .pi288( pi288 ) , .pi289( pi289 ) , .pi290( pi290 ) , .pi291( pi291 ) , .pi292( pi292 ) , .pi293( pi293 ) , .pi294( pi294 ) , .pi295( pi295 ) , .pi296( pi296 ) , .pi297( pi297 ) , .pi298( pi298 ) , .pi299( pi299 ) , .pi300( pi300 ) , .pi301( pi301 ) , .pi302( pi302 ) , .pi303( pi303 ) , .pi304( pi304 ) , .pi305( pi305 ) , .pi306( pi306 ) , .pi307( pi307 ) , .pi308( pi308 ) , .pi309( pi309 ) , .pi310( pi310 ) , .pi311( pi311 ) , .pi312( pi312 ) , .pi313( pi313 ) , .pi314( pi314 ) , .pi315( pi315 ) , .pi316( pi316 ) , .pi317( pi317 ) , .pi318( pi318 ) , .pi319( pi319 ) , .pi320( pi320 ) , .pi321( pi321 ) , .pi322( pi322 ) , .pi323( pi323 ) , .pi324( pi324 ) , .pi325( pi325 ) , .pi326( pi326 ) , .pi327( pi327 ) , .pi328( pi328 ) , .pi329( pi329 ) , .pi330( pi330 ) , .pi331( pi331 ) , .pi332( pi332 ) , .pi333( pi333 ) , .pi334( pi334 ) , .pi335( pi335 ) , .pi336( pi336 ) , .pi337( pi337 ) , .pi338( pi338 ) , .pi339( pi339 ) , .pi340( pi340 ) , .pi341( pi341 ) , .pi342( pi342 ) , .pi343( pi343 ) , .pi344( pi344 ) , .pi345( pi345 ) , .pi346( pi346 ) , .pi347( pi347 ) , .pi348( pi348 ) , .pi349( pi349 ) , .pi350( pi350 ) , .pi351( pi351 ) , .pi352( pi352 ) , .pi353( pi353 ) , .pi354( pi354 ) , .pi355( pi355 ) , .pi356( pi356 ) , .pi357( pi357 ) , .pi358( pi358 ) , .pi359( pi359 ) , .pi360( pi360 ) , .pi361( pi361 ) , .pi362( pi362 ) , .pi363( pi363 ) , .pi364( pi364 ) , .pi365( pi365 ) , .pi366( pi366 ) , .pi367( pi367 ) , .pi368( pi368 ) , .pi369( pi369 ) , .pi370( pi370 ) , .pi371( pi371 ) , .pi372( pi372 ) , .pi373( pi373 ) , .pi374( pi374 ) , .pi375( pi375 ) , .pi376( pi376 ) , .pi377( pi377 ) , .pi378( pi378 ) , .pi379( pi379 ) , .pi380( pi380 ) , .pi381( pi381 ) , .pi382( pi382 ) , .pi383( pi383 ) , .pi384( pi384 ) , .pi385( pi385 ) , .pi386( pi386 ) , .pi387( pi387 ) , .pi388( pi388 ) , .pi389( pi389 ) , .pi390( pi390 ) , .pi391( pi391 ) , .pi392( pi392 ) , .pi393( pi393 ) , .pi394( pi394 ) , .pi395( pi395 ) , .pi396( pi396 ) , .pi397( pi397 ) , .pi398( pi398 ) , .pi399( pi399 ) , .pi400( pi400 ) , .pi401( pi401 ) , .pi402( pi402 ) , .pi403( pi403 ) , .pi404( pi404 ) , .pi405( pi405 ) , .pi406( pi406 ) , .pi407( pi407 ) , .pi408( pi408 ) , .pi409( pi409 ) , .pi410( pi410 ) , .pi411( pi411 ) , .pi412( pi412 ) , .pi413( pi413 ) , .pi414( pi414 ) , .pi415( pi415 ) , .pi416( pi416 ) , .pi417( pi417 ) , .pi418( pi418 ) , .pi419( pi419 ) , .pi420( pi420 ) , .pi421( pi421 ) , .pi422( pi422 ) , .pi423( pi423 ) , .pi424( pi424 ) , .pi425( pi425 ) , .pi426( pi426 ) , .pi427( pi427 ) , .pi428( pi428 ) , .pi429( pi429 ) , .pi430( pi430 ) , .pi431( pi431 ) , .pi432( pi432 ) , .pi433( pi433 ) , .pi434( pi434 ) , .pi435( pi435 ) , .pi436( pi436 ) , .pi437( pi437 ) , .pi438( pi438 ) , .pi439( pi439 ) , .pi440( pi440 ) , .pi441( pi441 ) , .pi442( pi442 ) , .pi443( pi443 ) , .pi444( pi444 ) , .pi445( pi445 ) , .pi446( pi446 ) , .pi447( pi447 ) , .pi448( pi448 ) , .pi449( pi449 ) , .pi450( pi450 ) , .pi451( pi451 ) , .pi452( pi452 ) , .pi453( pi453 ) , .pi454( pi454 ) , .pi455( pi455 ) , .pi456( pi456 ) , .pi457( pi457 ) , .pi458( pi458 ) , .pi459( pi459 ) , .pi460( pi460 ) , .pi461( pi461 ) , .pi462( pi462 ) , .pi463( pi463 ) , .pi464( pi464 ) , .pi465( pi465 ) , .pi466( pi466 ) , .pi467( pi467 ) , .pi468( pi468 ) , .pi469( pi469 ) , .pi470( pi470 ) , .pi471( pi471 ) , .pi472( pi472 ) , .pi473( pi473 ) , .pi474( pi474 ) , .pi475( pi475 ) , .pi476( pi476 ) , .pi477( pi477 ) , .pi478( pi478 ) , .pi479( pi479 ) , .pi480( pi480 ) , .pi481( pi481 ) , .pi482( pi482 ) , .pi483( pi483 ) , .pi484( pi484 ) , .pi485( pi485 ) , .pi486( pi486 ) , .pi487( pi487 ) , .pi488( pi488 ) , .pi489( pi489 ) , .pi490( pi490 ) , .pi491( pi491 ) , .pi492( pi492 ) , .pi493( pi493 ) , .pi494( pi494 ) , .pi495( pi495 ) , .pi496( pi496 ) , .pi497( pi497 ) , .pi498( pi498 ) , .pi499( pi499 ) , .pi500( pi500 ) , .pi501( pi501 ) , .pi502( pi502 ) , .pi503( pi503 ) , .pi504( pi504 ) , .pi505( pi505 ) , .pi506( pi506 ) , .pi507( pi507 ) , .pi508( pi508 ) , .pi509( pi509 ) , .pi510( pi510 ) , .pi511( pi511 ) , .po000( po000 ) , .po001( po001 ) , .po002( po002 ) , .po003( po003 ) , .po004( po004 ) , .po005( po005 ) , .po006( po006 ) , .po007( po007 ) , .po008( po008 ) , .po009( po009 ) , .po010( po010 ) , .po011( po011 ) , .po012( po012 ) , .po013( po013 ) , .po014( po014 ) , .po015( po015 ) , .po016( po016 ) , .po017( po017 ) , .po018( po018 ) , .po019( po019 ) , .po020( po020 ) , .po021( po021 ) , .po022( po022 ) , .po023( po023 ) , .po024( po024 ) , .po025( po025 ) , .po026( po026 ) , .po027( po027 ) , .po028( po028 ) , .po029( po029 ) , .po030( po030 ) , .po031( po031 ) , .po032( po032 ) , .po033( po033 ) , .po034( po034 ) , .po035( po035 ) , .po036( po036 ) , .po037( po037 ) , .po038( po038 ) , .po039( po039 ) , .po040( po040 ) , .po041( po041 ) , .po042( po042 ) , .po043( po043 ) , .po044( po044 ) , .po045( po045 ) , .po046( po046 ) , .po047( po047 ) , .po048( po048 ) , .po049( po049 ) , .po050( po050 ) , .po051( po051 ) , .po052( po052 ) , .po053( po053 ) , .po054( po054 ) , .po055( po055 ) , .po056( po056 ) , .po057( po057 ) , .po058( po058 ) , .po059( po059 ) , .po060( po060 ) , .po061( po061 ) , .po062( po062 ) , .po063( po063 ) , .po064( po064 ) , .po065( po065 ) , .po066( po066 ) , .po067( po067 ) , .po068( po068 ) , .po069( po069 ) , .po070( po070 ) , .po071( po071 ) , .po072( po072 ) , .po073( po073 ) , .po074( po074 ) , .po075( po075 ) , .po076( po076 ) , .po077( po077 ) , .po078( po078 ) , .po079( po079 ) , .po080( po080 ) , .po081( po081 ) , .po082( po082 ) , .po083( po083 ) , .po084( po084 ) , .po085( po085 ) , .po086( po086 ) , .po087( po087 ) , .po088( po088 ) , .po089( po089 ) , .po090( po090 ) , .po091( po091 ) , .po092( po092 ) , .po093( po093 ) , .po094( po094 ) , .po095( po095 ) , .po096( po096 ) , .po097( po097 ) , .po098( po098 ) , .po099( po099 ) , .po100( po100 ) , .po101( po101 ) , .po102( po102 ) , .po103( po103 ) , .po104( po104 ) , .po105( po105 ) , .po106( po106 ) , .po107( po107 ) , .po108( po108 ) , .po109( po109 ) , .po110( po110 ) , .po111( po111 ) , .po112( po112 ) , .po113( po113 ) , .po114( po114 ) , .po115( po115 ) , .po116( po116 ) , .po117( po117 ) , .po118( po118 ) , .po119( po119 ) , .po120( po120 ) , .po121( po121 ) , .po122( po122 ) , .po123( po123 ) , .po124( po124 ) , .po125( po125 ) , .po126( po126 ) , .po127( po127 ) , .po128( po128 ) , .po129( po129 ) );
endmodule

module top(pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511, po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129);
  input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129;
  wire n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, tpo000, tpo001, tpo002, tpo003, tpo004, tpo005, tpo006, tpo007, tpo008, tpo009, tpo010, tpo011, tpo012, tpo013, tpo014, tpo015, tpo016, tpo017, tpo018, tpo019, tpo020, tpo021, tpo022, tpo023, tpo024, tpo025, tpo026, tpo027, tpo028, tpo029, tpo030, tpo031, tpo032, tpo033, tpo034, tpo035, tpo036, tpo037, tpo038, tpo039, tpo040, tpo041, tpo042, tpo043, tpo044, tpo045, tpo046, tpo047, tpo048, tpo049, tpo050, tpo051, tpo052, tpo053, tpo054, tpo055, tpo056, tpo057, tpo058, tpo059, tpo060, tpo061, tpo062, tpo063, tpo064, tpo065, tpo066, tpo067, tpo068, tpo069, tpo070, tpo071, tpo072, tpo073, tpo074, tpo075, tpo076, tpo077, tpo078, tpo079, tpo080, tpo081, tpo082, tpo083, tpo084, tpo085, tpo086, tpo087, tpo088, tpo089, tpo090, tpo091, tpo092, tpo093, tpo094, tpo095, tpo096, tpo097, tpo098, tpo099, tpo100, tpo101, tpo102, tpo103, tpo104, tpo105, tpo106, tpo107, tpo108, tpo109, tpo110, tpo111, tpo112, tpo113, tpo114, tpo115, tpo116, tpo117, tpo118, tpo119, tpo120, tpo121, tpo122, tpo123, tpo124, tpo125, tpo126, tpo127, tpo128, tpo129;
  assign po000 = ~tpo000;
  assign po001 = ~tpo001;
  assign po002 = ~tpo002;
  assign po003 = ~tpo003;
  assign po004 = ~tpo004;
  assign po005 = ~tpo005;
  assign po006 = ~tpo006;
  assign po007 = ~tpo007;
  assign po008 = ~tpo008;
  assign po009 = ~tpo009;
  assign po010 = ~tpo010;
  assign po011 = ~tpo011;
  assign po012 = ~tpo012;
  assign po013 = ~tpo013;
  assign po014 = ~tpo014;
  assign po015 = ~tpo015;
  assign po016 = ~tpo016;
  assign po017 = ~tpo017;
  assign po018 = ~tpo018;
  assign po019 = ~tpo019;
  assign po020 = ~tpo020;
  assign po021 = ~tpo021;
  assign po022 = ~tpo022;
  assign po023 = ~tpo023;
  assign po024 = ~tpo024;
  assign po025 = ~tpo025;
  assign po026 = ~tpo026;
  assign po027 = ~tpo027;
  assign po028 = ~tpo028;
  assign po029 = ~tpo029;
  assign po030 = ~tpo030;
  assign po031 = ~tpo031;
  assign po032 = ~tpo032;
  assign po033 = ~tpo033;
  assign po034 = ~tpo034;
  assign po035 = ~tpo035;
  assign po036 = ~tpo036;
  assign po037 = ~tpo037;
  assign po038 = ~tpo038;
  assign po039 = ~tpo039;
  assign po040 = ~tpo040;
  assign po041 = ~tpo041;
  assign po042 = ~tpo042;
  assign po043 = ~tpo043;
  assign po044 = ~tpo044;
  assign po045 = ~tpo045;
  assign po046 = ~tpo046;
  assign po047 = ~tpo047;
  assign po048 = ~tpo048;
  assign po049 = ~tpo049;
  assign po050 = ~tpo050;
  assign po051 = ~tpo051;
  assign po052 = ~tpo052;
  assign po053 = ~tpo053;
  assign po054 = ~tpo054;
  assign po055 = ~tpo055;
  assign po056 = ~tpo056;
  assign po057 = ~tpo057;
  assign po058 = ~tpo058;
  assign po059 = ~tpo059;
  assign po060 = ~tpo060;
  assign po061 = ~tpo061;
  assign po062 = ~tpo062;
  assign po063 = ~tpo063;
  assign po064 = ~tpo064;
  assign po065 = ~tpo065;
  assign po066 = ~tpo066;
  assign po067 = ~tpo067;
  assign po068 = ~tpo068;
  assign po069 = ~tpo069;
  assign po070 = ~tpo070;
  assign po071 = ~tpo071;
  assign po072 = ~tpo072;
  assign po073 = ~tpo073;
  assign po074 = ~tpo074;
  assign po075 = ~tpo075;
  assign po076 = ~tpo076;
  assign po077 = ~tpo077;
  assign po078 = ~tpo078;
  assign po079 = ~tpo079;
  assign po080 = ~tpo080;
  assign po081 = ~tpo081;
  assign po082 = ~tpo082;
  assign po083 = ~tpo083;
  assign po084 = ~tpo084;
  assign po085 = ~tpo085;
  assign po086 = ~tpo086;
  assign po087 = ~tpo087;
  assign po088 = ~tpo088;
  assign po089 = ~tpo089;
  assign po090 = ~tpo090;
  assign po091 = ~tpo091;
  assign po092 = ~tpo092;
  assign po093 = ~tpo093;
  assign po094 = ~tpo094;
  assign po095 = ~tpo095;
  assign po096 = ~tpo096;
  assign po097 = ~tpo097;
  assign po098 = ~tpo098;
  assign po099 = ~tpo099;
  assign po100 = ~tpo100;
  assign po101 = ~tpo101;
  assign po102 = ~tpo102;
  assign po103 = ~tpo103;
  assign po104 = ~tpo104;
  assign po105 = ~tpo105;
  assign po106 = ~tpo106;
  assign po107 = ~tpo107;
  assign po108 = ~tpo108;
  assign po109 = ~tpo109;
  assign po110 = ~tpo110;
  assign po111 = ~tpo111;
  assign po112 = ~tpo112;
  assign po113 = ~tpo113;
  assign po114 = ~tpo114;
  assign po115 = ~tpo115;
  assign po116 = ~tpo116;
  assign po117 = ~tpo117;
  assign po118 = ~tpo118;
  assign po119 = ~tpo119;
  assign po120 = ~tpo120;
  assign po121 = ~tpo121;
  assign po122 = ~tpo122;
  assign po123 = ~tpo123;
  assign po124 = ~tpo124;
  assign po125 = ~tpo125;
  assign po126 = ~tpo126;
  assign po127 = tpo127;
  assign po128 = ~tpo128;
  assign po129 = ~tpo129;
  max_0 U0 ( .pi00( pi321 ), .pi01( pi322 ), .pi02( pi323 ), .pi03( pi449 ), .pi04( pi450 ), .pi05( pi451 ), .pi06( n75 ), .pi07( n97 ), .pi08( n211 ), .pi09( n212 ), .pi10( n213 ), .pi11( n214 ), .pi12( n215 ), .pi13( n217 ), .pi14( tpo129 ), .po0( n76 ), .po1( n77 ), .po2( n218 ), .po3( tpo065 ), .po4( tpo066 ), .po5( tpo067 ) );
  max_1 U1 ( .pi00( pi324 ), .pi01( pi325 ), .pi02( pi326 ), .pi03( pi327 ), .pi04( pi452 ), .pi05( pi453 ), .pi06( pi454 ), .pi07( pi455 ), .pi08( n76 ), .pi09( n77 ), .pi10( n97 ), .pi11( n216 ), .pi12( n218 ), .pi13( n219 ), .pi14( n220 ), .pi15( n221 ), .pi16( n223 ), .pi17( tpo129 ), .po0( n78 ), .po1( n217 ), .po2( n224 ), .po3( tpo068 ), .po4( tpo069 ), .po5( tpo070 ), .po6( tpo071 ) );
  max_2 U2 ( .pi0( pi194 ), .po0(  ) );
  max_3 U3 ( .pi00( pi065 ), .pi01( pi066 ), .pi02( pi067 ), .pi03( pi068 ), .pi04( pi069 ), .pi05( pi070 ), .pi06( pi071 ), .pi07( pi193 ), .pi08( pi194 ), .pi09( pi195 ), .pi10( pi196 ), .pi11( pi197 ), .pi12( pi198 ), .pi13( pi199 ), .pi14( n21 ), .pi15( n22 ), .pi16( n23 ), .pi17( n47 ), .po0( n24 ), .po1( n213 ), .po2( n214 ), .po3( n215 ), .po4( n216 ), .po5( n219 ), .po6( n220 ), .po7( n221 ) );
  max_4 U4 ( .pi00( pi332 ), .pi01( pi333 ), .pi02( pi334 ), .pi03( pi335 ), .pi04( pi460 ), .pi05( pi461 ), .pi06( pi462 ), .pi07( pi463 ), .pi08( n79 ), .pi09( n80 ), .pi10( n97 ), .po0( n81 ), .po1( n117 ), .po2( n118 ), .po3( n119 ), .po4( n229 ) );
  max_5 U5 ( .pi00( pi077 ), .pi01( pi078 ), .pi02( pi079 ), .pi03( pi205 ), .pi04( pi206 ), .pi05( pi207 ), .pi06( n25 ), .pi07( n26 ), .pi08( n47 ), .pi09( n117 ), .pi10( n118 ), .pi11( n228 ), .pi12( n229 ), .pi13( tpo129 ), .po0( n27 ), .po1( n28 ), .po2( n230 ), .po3( tpo077 ), .po4( tpo078 ), .po5( tpo079 ) );
  max_6 U6 ( .pi00( pi328 ), .pi01( pi329 ), .pi02( pi330 ), .pi03( pi331 ), .pi04( pi456 ), .pi05( pi457 ), .pi06( pi458 ), .pi07( pi459 ), .pi08( n78 ), .pi09( n97 ), .pi10( n119 ), .pi11( n120 ), .pi12( n222 ), .pi13( n224 ), .pi14( n225 ), .pi15( n226 ), .pi16( n227 ), .pi17( tpo129 ), .po0( n79 ), .po1( n223 ), .po2( n228 ), .po3( tpo072 ), .po4( tpo073 ), .po5( tpo074 ), .po6( tpo075 ), .po7( tpo076 ) );
  max_7 U7 ( .pi00( pi072 ), .pi01( pi073 ), .pi02( pi074 ), .pi03( pi075 ), .pi04( pi076 ), .pi05( pi200 ), .pi06( pi201 ), .pi07( pi202 ), .pi08( pi203 ), .pi09( pi204 ), .pi10( n24 ), .pi11( n47 ), .po0( n23 ), .po1( n25 ), .po2( n26 ), .po3( n120 ), .po4( n222 ), .po5( n225 ), .po6( n226 ), .po7( n227 ) );
  max_8 U8 ( .pi00( pi084 ), .pi01( pi085 ), .pi02( pi086 ), .pi03( pi212 ), .pi04( pi213 ), .pi05( pi214 ), .pi06( n29 ), .pi07( n30 ), .pi08( n47 ), .pi09( n115 ), .pi10( n234 ), .pi11( n235 ), .pi12( n236 ), .pi13( n237 ), .pi14( tpo129 ), .po0( n31 ), .po1( n238 ), .po2( tpo084 ), .po3( tpo085 ), .po4( tpo086 ) );
  max_9 U9 ( .pi00( pi340 ), .pi01( pi341 ), .pi02( pi342 ), .pi03( pi343 ), .pi04( pi468 ), .pi05( pi469 ), .pi06( pi470 ), .pi07( pi471 ), .pi08( n82 ), .pi09( n97 ), .po0( n83 ), .po1( n114 ), .po2( n115 ), .po3( n236 ), .po4( n237 ) );
  max_10 U10 ( .pi00( pi080 ), .pi01( pi081 ), .pi02( pi082 ), .pi03( pi083 ), .pi04( pi208 ), .pi05( pi209 ), .pi06( pi210 ), .pi07( pi211 ), .pi08( n27 ), .pi09( n28 ), .pi10( n47 ), .pi11( n97 ), .pi12( tpo129 ), .po0( n29 ), .po1( n30 ), .po2( n116 ), .po3( n231 ), .po4( n232 ), .po5( n233 ), .po6( tpo128 ) );
  max_11 U11 ( .pi00( pi336 ), .pi01( pi337 ), .pi02( pi338 ), .pi03( pi339 ), .pi04( pi464 ), .pi05( pi465 ), .pi06( pi466 ), .pi07( pi467 ), .pi08( n81 ), .pi09( n97 ), .pi10( n116 ), .pi11( n230 ), .pi12( n231 ), .pi13( n232 ), .pi14( n233 ), .pi15( tpo129 ), .po0( n80 ), .po1( n82 ), .po2( n234 ), .po3( n235 ), .po4( tpo080 ), .po5( tpo081 ), .po6( tpo082 ), .po7( tpo083 ) );
  max_12 U12 ( .pi00( pi087 ), .pi01( pi088 ), .pi02( pi089 ), .pi03( pi090 ), .pi04( pi215 ), .pi05( pi216 ), .pi06( pi217 ), .pi07( pi218 ), .pi08( n31 ), .pi09( n47 ), .pi10( n113 ), .pi11( n114 ), .pi12( n238 ), .pi13( n239 ), .pi14( n240 ), .pi15( n242 ), .pi16( tpo129 ), .po0( n32 ), .po1( n243 ), .po2( tpo087 ), .po3( tpo088 ), .po4( tpo089 ), .po5( tpo090 ) );
  max_13 U13 ( .pi0( pi344 ), .pi1( pi345 ), .pi2( pi346 ), .pi3( pi472 ), .pi4( pi473 ), .pi5( pi474 ), .pi6( n83 ), .pi7( n84 ), .pi8( n97 ), .po0( n85 ), .po1( n113 ), .po2( n239 ), .po3( n240 ) );
  max_14 U14 ( .pi00( pi347 ), .pi01( pi348 ), .pi02( pi349 ), .pi03( pi350 ), .pi04( pi475 ), .pi05( pi476 ), .pi06( pi477 ), .pi07( pi478 ), .pi08( n85 ), .pi09( n86 ), .pi10( n97 ), .pi11( n241 ), .pi12( n243 ), .pi13( n244 ), .pi14( n245 ), .pi15( n246 ), .pi16( n247 ), .pi17( tpo129 ), .po0( n84 ), .po1( n87 ), .po2( n242 ), .po3( n248 ), .po4( tpo091 ), .po5( tpo092 ), .po6( tpo093 ), .po7( tpo094 ) );
  max_15 U15 ( .pi00( pi091 ), .pi01( pi092 ), .pi02( pi093 ), .pi03( pi094 ), .pi04( pi219 ), .pi05( pi220 ), .pi06( pi221 ), .pi07( pi222 ), .pi08( n32 ), .pi09( n47 ), .po0( n33 ), .po1( n241 ), .po2( n244 ), .po3( n245 ), .po4( n246 ) );
  max_16 U16 ( .pi00( pi095 ), .pi01( pi096 ), .pi02( pi097 ), .pi03( pi098 ), .pi04( pi099 ), .pi05( pi223 ), .pi06( pi224 ), .pi07( pi225 ), .pi08( pi226 ), .pi09( pi227 ), .pi10( n33 ), .pi11( n47 ), .pi12( n112 ), .pi13( n248 ), .pi14( tpo129 ), .po0( n34 ), .po1( n35 ), .po2( n110 ), .po3( n111 ), .po4( n247 ), .po5( n249 ), .po6( n250 ), .po7( n251 ), .po8( tpo095 ) );
  max_17 U17 ( .pi00( pi351 ), .pi01( pi352 ), .pi02( pi353 ), .pi03( pi354 ), .pi04( pi355 ), .pi05( pi479 ), .pi06( pi480 ), .pi07( pi481 ), .pi08( pi482 ), .pi09( pi483 ), .pi10( n87 ), .pi11( n97 ), .pi12( n110 ), .pi13( n111 ), .pi14( n249 ), .pi15( n250 ), .pi16( n251 ), .pi17( tpo129 ), .po0( n86 ), .po1( n88 ), .po2( n112 ), .po3( n252 ), .po4( tpo096 ), .po5( tpo097 ), .po6( tpo098 ), .po7( tpo099 ) );
  max_18 U18 ( .pi00( pi356 ), .pi01( pi357 ), .pi02( pi358 ), .pi03( pi359 ), .pi04( pi484 ), .pi05( pi485 ), .pi06( pi486 ), .pi07( pi487 ), .pi08( n88 ), .pi09( n97 ), .pi10( n108 ), .pi11( n109 ), .pi12( n252 ), .pi13( n253 ), .pi14( n254 ), .pi15( tpo129 ), .po0( n89 ), .po1( n255 ), .po2( tpo100 ), .po3( tpo101 ), .po4( tpo102 ), .po5( tpo103 ) );
  max_19 U19 ( .pi00( pi100 ), .pi01( pi101 ), .pi02( pi102 ), .pi03( pi103 ), .pi04( pi228 ), .pi05( pi229 ), .pi06( pi230 ), .pi07( pi231 ), .pi08( n34 ), .pi09( n35 ), .pi10( n47 ), .po0( n36 ), .po1( n37 ), .po2( n108 ), .po3( n109 ), .po4( n253 ), .po5( n254 ) );
  max_20 U20 ( .pi00( pi104 ), .pi01( pi105 ), .pi02( pi106 ), .pi03( pi107 ), .pi04( pi232 ), .pi05( pi233 ), .pi06( pi234 ), .pi07( pi235 ), .pi08( n36 ), .pi09( n37 ), .pi10( n47 ), .po0( n38 ), .po1( n39 ), .po2( n105 ), .po3( n106 ), .po4( n107 ), .po5( n256 ) );
  max_21 U21 ( .pi00( pi360 ), .pi01( pi361 ), .pi02( pi362 ), .pi03( pi363 ), .pi04( pi488 ), .pi05( pi489 ), .pi06( pi490 ), .pi07( pi491 ), .pi08( n89 ), .pi09( n97 ), .pi10( n105 ), .pi11( n106 ), .pi12( n107 ), .pi13( n255 ), .pi14( n256 ), .pi15( tpo129 ), .po0( n90 ), .po1( n257 ), .po2( n258 ), .po3( tpo104 ), .po4( tpo105 ), .po5( tpo106 ), .po6( tpo107 ) );
  max_22 U22 ( .pi00( pi108 ), .pi01( pi109 ), .pi02( pi110 ), .pi03( pi111 ), .pi04( pi236 ), .pi05( pi237 ), .pi06( pi238 ), .pi07( pi239 ), .pi08( n38 ), .pi09( n39 ), .pi10( n47 ), .po0( n40 ), .po1( n41 ), .po2( n103 ), .po3( n104 ), .po4( n259 ), .po5( n260 ) );
  max_23 U23 ( .pi00( pi364 ), .pi01( pi365 ), .pi02( pi366 ), .pi03( pi367 ), .pi04( pi492 ), .pi05( pi493 ), .pi06( pi494 ), .pi07( pi495 ), .pi08( n90 ), .pi09( n97 ), .pi10( n103 ), .pi11( n104 ), .pi12( n257 ), .pi13( n258 ), .pi14( n259 ), .pi15( n260 ), .pi16( tpo129 ), .po0( n91 ), .po1( n261 ), .po2( n262 ), .po3( tpo108 ), .po4( tpo109 ), .po5( tpo110 ), .po6( tpo111 ) );
  max_24 U24 ( .pi00( pi116 ), .pi01( pi117 ), .pi02( pi118 ), .pi03( pi244 ), .pi04( pi245 ), .pi05( pi246 ), .pi06( pi372 ), .pi07( pi373 ), .pi08( pi374 ), .pi09( pi500 ), .pi10( pi501 ), .pi11( pi502 ), .pi12( n42 ), .pi13( n43 ), .pi14( n47 ), .pi15( n92 ), .pi16( n93 ), .pi17( n97 ), .pi18( n265 ), .pi19( n266 ), .pi20( tpo129 ), .po0( n44 ), .po1( n94 ), .po2( n267 ), .po3( n268 ), .po4( n269 ), .po5( tpo117 ), .po6( tpo118 ) );
  max_25 U25 ( .pi0( n267 ), .pi1( n268 ), .pi2( tpo129 ), .po0( tpo116 ) );
  max_26 U26 ( .pi00( pi368 ), .pi01( pi369 ), .pi02( pi370 ), .pi03( pi371 ), .pi04( pi496 ), .pi05( pi497 ), .pi06( pi498 ), .pi07( pi499 ), .pi08( n91 ), .pi09( n97 ), .pi10( n101 ), .pi11( n102 ), .pi12( n261 ), .pi13( n262 ), .pi14( n263 ), .pi15( n264 ), .pi16( tpo129 ), .po0( n92 ), .po1( n93 ), .po2( n265 ), .po3( n266 ), .po4( tpo112 ), .po5( tpo113 ), .po6( tpo114 ), .po7( tpo115 ) );
  max_27 U27 ( .pi00( pi112 ), .pi01( pi113 ), .pi02( pi114 ), .pi03( pi115 ), .pi04( pi240 ), .pi05( pi241 ), .pi06( pi242 ), .pi07( pi243 ), .pi08( n40 ), .pi09( n41 ), .pi10( n47 ), .po0( n42 ), .po1( n101 ), .po2( n102 ), .po3( n263 ), .po4( n264 ) );
  max_28 U28 ( .pi00( pi379 ), .pi01( pi380 ), .pi02( pi381 ), .pi03( pi382 ), .pi04( pi383 ), .pi05( pi507 ), .pi06( pi508 ), .pi07( pi509 ), .pi08( pi510 ), .pi09( pi511 ), .pi10( n49 ), .pi11( n96 ), .pi12( n98 ), .pi13( n272 ), .pi14( n274 ), .pi15( n275 ), .pi16( n276 ), .po0( n95 ), .po1( n97 ), .po2( n273 ), .po3( tpo129 ), .po4( tpo123 ), .po5( tpo125 ), .po6( tpo126 ), .po7( tpo127 ) );
  max_29 U29 ( .pi00( pi123 ), .pi01( pi124 ), .pi02( pi125 ), .pi03( pi126 ), .pi04( pi127 ), .pi05( pi251 ), .pi06( pi252 ), .pi07( pi253 ), .pi08( pi254 ), .pi09( pi255 ), .pi10( n46 ), .pi11( n273 ), .pi12( tpo129 ), .po0( n45 ), .po1( n47 ), .po2( n49 ), .po3( n98 ), .po4( n274 ), .po5( n275 ), .po6( n276 ), .po7( tpo124 ) );
  max_30 U30 ( .pi00( pi375 ), .pi01( pi376 ), .pi02( pi377 ), .pi03( pi378 ), .pi04( pi503 ), .pi05( pi504 ), .pi06( pi505 ), .pi07( pi506 ), .pi08( n94 ), .pi09( n95 ), .pi10( n97 ), .po0( n96 ), .po1( n99 ), .po2( n100 ), .po3( n270 ), .po4( n271 ) );
  max_31 U31 ( .pi00( pi119 ), .pi01( pi120 ), .pi02( pi121 ), .pi03( pi122 ), .pi04( pi247 ), .pi05( pi248 ), .pi06( pi249 ), .pi07( pi250 ), .pi08( n44 ), .pi09( n45 ), .pi10( n47 ), .pi11( n99 ), .pi12( n100 ), .pi13( n269 ), .pi14( n270 ), .pi15( n271 ), .pi16( tpo129 ), .po0( n43 ), .po1( n46 ), .po2( n272 ), .po3( tpo119 ), .po4( tpo120 ), .po5( tpo121 ), .po6( tpo122 ) );
  max_32 U32 ( .pi00( pi264 ), .pi01( pi265 ), .pi02( pi266 ), .pi03( pi392 ), .pi04( pi393 ), .pi05( pi394 ), .pi06( n52 ), .pi07( n53 ), .pi08( n97 ), .pi09( n131 ), .pi10( n140 ), .pi11( n142 ), .pi12( n143 ), .pi13( tpo129 ), .po0( n54 ), .po1( n141 ), .po2( n144 ), .po3( tpo008 ), .po4( tpo009 ), .po5( tpo010 ) );
  max_33 U33 ( .pi00( pi008 ), .pi01( pi009 ), .pi02( pi010 ), .pi03( pi011 ), .pi04( pi136 ), .pi05( pi137 ), .pi06( pi138 ), .pi07( pi139 ), .pi08( n2 ), .pi09( n47 ), .po0( n3 ), .po1( n130 ), .po2( n131 ), .po3( n140 ), .po4( n143 ) );
  max_34 U34 ( .pi00( pi012 ), .pi01( pi013 ), .pi02( pi014 ), .pi03( pi015 ), .pi04( pi140 ), .pi05( pi141 ), .pi06( pi142 ), .pi07( pi143 ), .pi08( n3 ), .pi09( n47 ), .pi10( n129 ), .pi11( n130 ), .pi12( n144 ), .pi13( n145 ), .pi14( n146 ), .pi15( n147 ), .pi16( n148 ), .pi17( n150 ), .pi18( tpo129 ), .po0( n4 ), .po1( n151 ), .po2( tpo011 ), .po3( tpo012 ), .po4( tpo013 ), .po5( tpo014 ), .po6( tpo015 ) );
  max_35 U35 ( .pi00( pi267 ), .pi01( pi268 ), .pi02( pi269 ), .pi03( pi270 ), .pi04( pi271 ), .pi05( pi395 ), .pi06( pi396 ), .pi07( pi397 ), .pi08( pi398 ), .pi09( pi399 ), .pi10( n54 ), .pi11( n97 ), .po0( n55 ), .po1( n56 ), .po2( n129 ), .po3( n145 ), .po4( n146 ), .po5( n147 ), .po6( n148 ) );
  max_36 U36 ( .pi00( pi000 ), .pi01( pi001 ), .pi02( pi002 ), .pi03( pi003 ), .pi04( pi128 ), .pi05( pi129 ), .pi06( pi130 ), .pi07( pi131 ), .pi08( n0 ), .pi09( n47 ), .po0( n1 ), .po1( n48 ), .po2( n133 ), .po3( n134 ), .po4( n135 ) );
  max_37 U37 ( .pi00( pi256 ), .pi01( pi257 ), .pi02( pi258 ), .pi03( pi259 ), .pi04( pi384 ), .pi05( pi385 ), .pi06( pi386 ), .pi07( pi387 ), .pi08( n48 ), .pi09( n97 ), .pi10( n133 ), .pi11( n134 ), .pi12( n135 ), .pi13( tpo129 ), .po0( n50 ), .po1( n51 ), .po2( n136 ), .po3( tpo000 ), .po4( tpo001 ), .po5( tpo002 ), .po6( tpo003 ) );
  max_38 U38 ( .pi00( pi004 ), .pi01( pi005 ), .pi02( pi006 ), .pi03( pi007 ), .pi04( pi132 ), .pi05( pi133 ), .pi06( pi134 ), .pi07( pi135 ), .pi08( n1 ), .pi09( n47 ), .pi10( n132 ), .pi11( n136 ), .pi12( n137 ), .pi13( n138 ), .pi14( n139 ), .pi15( n141 ), .pi16( tpo129 ), .po0( n0 ), .po1( n2 ), .po2( n142 ), .po3( tpo004 ), .po4( tpo005 ), .po5( tpo006 ), .po6( tpo007 ) );
  max_39 U39 ( .pi00( pi260 ), .pi01( pi261 ), .pi02( pi262 ), .pi03( pi263 ), .pi04( pi388 ), .pi05( pi389 ), .pi06( pi390 ), .pi07( pi391 ), .pi08( n50 ), .pi09( n51 ), .pi10( n97 ), .po0( n52 ), .po1( n53 ), .po2( n132 ), .po3( n137 ), .po4( n138 ), .po5( n139 ) );
  max_40 U40 ( .pi00( pi272 ), .pi01( pi273 ), .pi02( pi274 ), .pi03( pi275 ), .pi04( pi276 ), .pi05( pi400 ), .pi06( pi401 ), .pi07( pi402 ), .pi08( pi403 ), .pi09( pi404 ), .pi10( n55 ), .pi11( n56 ), .pi12( n97 ), .po0( n57 ), .po1( n127 ), .po2( n128 ), .po3( n149 ), .po4( n152 ), .po5( n153 ) );
  max_41 U41 ( .pi00( pi016 ), .pi01( pi017 ), .pi02( pi018 ), .pi03( pi019 ), .pi04( pi020 ), .pi05( pi144 ), .pi06( pi145 ), .pi07( pi146 ), .pi08( pi147 ), .pi09( pi148 ), .pi10( n4 ), .pi11( n47 ), .pi12( n127 ), .pi13( n128 ), .pi14( n149 ), .pi15( n151 ), .pi16( n152 ), .pi17( n153 ), .pi18( tpo129 ), .po0( n5 ), .po1( n150 ), .po2( n154 ), .po3( n155 ), .po4( tpo016 ), .po5( tpo017 ), .po6( tpo018 ), .po7( tpo019 ) );
  max_42 U42 ( .pi00( pi021 ), .pi01( pi022 ), .pi02( pi023 ), .pi03( pi149 ), .pi04( pi150 ), .pi05( pi151 ), .pi06( pi277 ), .pi07( pi278 ), .pi08( pi279 ), .pi09( pi405 ), .pi10( pi406 ), .pi11( pi407 ), .pi12( n5 ), .pi13( n47 ), .pi14( n57 ), .pi15( n58 ), .pi16( n97 ), .pi17( n155 ), .pi18( n156 ), .pi19( tpo129 ), .po0( n6 ), .po1( n7 ), .po2( n59 ), .po3( n157 ), .po4( n158 ), .po5( tpo021 ), .po6( tpo022 ), .po7( tpo023 ) );
  max_43 U43 ( .pi0( n153 ), .pi1( n154 ), .pi2( tpo129 ), .po0( n156 ), .po1( tpo020 ) );
  max_44 U44 ( .pi00( pi027 ), .pi01( pi028 ), .pi02( pi029 ), .pi03( pi030 ), .pi04( pi031 ), .pi05( pi155 ), .pi06( pi156 ), .pi07( pi157 ), .pi08( pi158 ), .pi09( pi159 ), .pi10( n8 ), .pi11( n47 ), .pi12( n161 ), .pi13( n163 ), .pi14( n164 ), .pi15( n165 ), .pi16( n166 ), .pi17( n167 ), .pi18( tpo129 ), .po0( n9 ), .po1( n10 ), .po2( n162 ), .po3( n168 ), .po4( n169 ), .po5( tpo028 ), .po6( tpo029 ), .po7( tpo030 ), .po8( tpo031 ) );
  max_45 U45 ( .pi00( pi283 ), .pi01( pi284 ), .pi02( pi285 ), .pi03( pi286 ), .pi04( pi287 ), .pi05( pi411 ), .pi06( pi412 ), .pi07( pi413 ), .pi08( pi414 ), .pi09( pi415 ), .pi10( n60 ), .pi11( n97 ), .po0( n61 ), .po1( n161 ), .po2( n164 ), .po3( n165 ), .po4( n166 ), .po5( n167 ) );
  max_46 U46 ( .pi0( pi024 ), .pi1( pi025 ), .pi2( pi026 ), .pi3( pi152 ), .pi4( pi153 ), .pi5( pi154 ), .pi6( n6 ), .pi7( n7 ), .pi8( n47 ), .po0( n8 ), .po1( n126 ), .po2( n159 ), .po3( n160 ) );
  max_47 U47 ( .pi00( pi280 ), .pi01( pi281 ), .pi02( pi282 ), .pi03( pi408 ), .pi04( pi409 ), .pi05( pi410 ), .pi06( n59 ), .pi07( n97 ), .pi08( n126 ), .pi09( n157 ), .pi10( n158 ), .pi11( n159 ), .pi12( n160 ), .pi13( n161 ), .pi14( n162 ), .pi15( tpo129 ), .po0( n58 ), .po1( n60 ), .po2( n163 ), .po3( tpo024 ), .po4( tpo025 ), .po5( tpo026 ), .po6( tpo027 ) );
  max_48 U48 ( .pi00( pi313 ), .pi01( pi314 ), .pi02( pi315 ), .pi03( pi441 ), .pi04( pi442 ), .pi05( pi443 ), .pi06( n72 ), .pi07( n97 ), .pi08( n122 ), .pi09( n123 ), .pi10( n202 ), .pi11( n203 ), .pi12( n204 ), .pi13( n205 ), .pi14( n206 ), .pi15( n207 ), .pi16( tpo129 ), .po0( n71 ), .po1( n73 ), .po2( n74 ), .po3( n208 ), .po4( tpo057 ), .po5( tpo058 ), .po6( tpo059 ), .po7( tpo060 ), .po8( tpo061 ) );
  max_49 U49 ( .pi00( pi316 ), .pi01( pi317 ), .pi02( pi318 ), .pi03( pi319 ), .pi04( pi320 ), .pi05( pi444 ), .pi06( pi445 ), .pi07( pi446 ), .pi08( pi447 ), .pi09( pi448 ), .pi10( n73 ), .pi11( n74 ), .pi12( n97 ), .po0( n75 ), .po1( n121 ), .po2( n122 ), .po3( n207 ), .po4( n209 ), .po5( n210 ) );
  max_50 U50 ( .pi00( pi060 ), .pi01( pi061 ), .pi02( pi062 ), .pi03( pi063 ), .pi04( pi064 ), .pi05( pi188 ), .pi06( pi189 ), .pi07( pi190 ), .pi08( pi191 ), .pi09( pi192 ), .pi10( n19 ), .pi11( n20 ), .pi12( n47 ), .pi13( n121 ), .pi14( n208 ), .pi15( n209 ), .pi16( n210 ), .pi17( tpo129 ), .po0( n21 ), .po1( n22 ), .po2( n123 ), .po3( n206 ), .po4( n211 ), .po5( n212 ), .po6( tpo062 ), .po7( tpo063 ), .po8( tpo064 ) );
  max_51 U51 ( .pi0( pi057 ), .pi1( pi058 ), .pi2( pi059 ), .pi3( pi185 ), .pi4( pi186 ), .pi5( pi187 ), .pi6( n18 ), .pi7( n47 ), .po0( n19 ), .po1( n20 ), .po2( n203 ), .po3( n204 ), .po4( n205 ) );
  max_52 U52 ( .pi00( pi052 ), .pi01( pi053 ), .pi02( pi054 ), .pi03( pi055 ), .pi04( pi056 ), .pi05( pi180 ), .pi06( pi181 ), .pi07( pi182 ), .pi08( pi183 ), .pi09( pi184 ), .pi10( n17 ), .pi11( n47 ), .pi12( n124 ), .pi13( n195 ), .pi14( n198 ), .pi15( n199 ), .pi16( n200 ), .pi17( n201 ), .pi18( tpo129 ), .po0( n18 ), .po1( n196 ), .po2( n202 ), .po3( tpo053 ), .po4( tpo054 ), .po5( tpo055 ), .po6( tpo056 ) );
  max_53 U53 ( .pi00( pi308 ), .pi01( pi309 ), .pi02( pi310 ), .pi03( pi311 ), .pi04( pi312 ), .pi05( pi436 ), .pi06( pi437 ), .pi07( pi438 ), .pi08( pi439 ), .pi09( pi440 ), .pi10( n70 ), .pi11( n71 ), .pi12( n97 ), .po0( n72 ), .po1( n124 ), .po2( n195 ), .po3( n199 ), .po4( n200 ), .po5( n201 ) );
  max_54 U54 ( .pi00( pi049 ), .pi01( pi050 ), .pi02( pi051 ), .pi03( pi177 ), .pi04( pi178 ), .pi05( pi179 ), .pi06( pi305 ), .pi07( pi306 ), .pi08( pi307 ), .pi09( pi433 ), .pi10( pi434 ), .pi11( pi435 ), .pi12( n16 ), .pi13( n47 ), .pi14( n69 ), .pi15( n97 ), .pi16( n194 ), .pi17( n197 ), .pi18( tpo129 ), .po0( n15 ), .po1( n17 ), .po2( n70 ), .po3( n193 ), .po4( n198 ), .po5( tpo049 ), .po6( tpo050 ), .po7( tpo051 ) );
  max_55 U55 ( .pi0( n195 ), .pi1( n196 ), .pi2( tpo129 ), .po0( n197 ), .po1( tpo052 ) );
  max_56 U56 ( .pi0( n175 ), .pi1( n176 ), .pi2( tpo129 ), .po0( tpo038 ) );
  max_57 U57 ( .pi00( pi036 ), .pi01( pi037 ), .pi02( pi038 ), .pi03( pi164 ), .pi04( pi165 ), .pi05( pi166 ), .pi06( pi292 ), .pi07( pi293 ), .pi08( pi294 ), .pi09( pi420 ), .pi10( pi421 ), .pi11( pi422 ), .pi12( n11 ), .pi13( n47 ), .pi14( n62 ), .pi15( n63 ), .pi16( n97 ), .pi17( n173 ), .pi18( n174 ), .pi19( n178 ), .pi20( tpo129 ), .po0( n12 ), .po1( n64 ), .po2( n175 ), .po3( n176 ), .po4( n179 ), .po5( tpo036 ), .po6( tpo037 ) );
  max_58 U58 ( .pi00( pi032 ), .pi01( pi033 ), .pi02( pi034 ), .pi03( pi035 ), .pi04( pi160 ), .pi05( pi161 ), .pi06( pi162 ), .pi07( pi163 ), .pi08( n9 ), .pi09( n10 ), .pi10( n47 ), .po0( n11 ), .po1( n125 ), .po2( n170 ), .po3( n171 ), .po4( n172 ) );
  max_59 U59 ( .pi00( pi288 ), .pi01( pi289 ), .pi02( pi290 ), .pi03( pi291 ), .pi04( pi416 ), .pi05( pi417 ), .pi06( pi418 ), .pi07( pi419 ), .pi08( n61 ), .pi09( n97 ), .pi10( n125 ), .pi11( n168 ), .pi12( n169 ), .pi13( n170 ), .pi14( n171 ), .pi15( n172 ), .pi16( tpo129 ), .po0( n62 ), .po1( n173 ), .po2( n174 ), .po3( tpo032 ), .po4( tpo033 ), .po5( tpo034 ), .po6( tpo035 ) );
  max_60 U60 ( .pi00( pi039 ), .pi01( pi040 ), .pi02( pi041 ), .pi03( pi042 ), .pi04( pi043 ), .pi05( pi167 ), .pi06( pi168 ), .pi07( pi169 ), .pi08( pi170 ), .pi09( pi171 ), .pi10( n12 ), .pi11( n47 ), .po0( n13 ), .po1( n14 ), .po2( n177 ), .po3( n180 ), .po4( n181 ), .po5( n182 ), .po6( n183 ) );
  max_61 U61 ( .pi00( pi295 ), .pi01( pi296 ), .pi02( pi297 ), .pi03( pi298 ), .pi04( pi423 ), .pi05( pi424 ), .pi06( pi425 ), .pi07( pi426 ), .pi08( n64 ), .pi09( n65 ), .pi10( n97 ), .pi11( n177 ), .pi12( n179 ), .pi13( n180 ), .pi14( n181 ), .pi15( n182 ), .pi16( n184 ), .pi17( tpo129 ), .po0( n63 ), .po1( n66 ), .po2( n178 ), .po3( n185 ), .po4( tpo039 ), .po5( tpo040 ), .po6( tpo041 ), .po7( tpo042 ) );
  max_62 U62 ( .pi00( pi044 ), .pi01( pi045 ), .pi02( pi046 ), .pi03( pi047 ), .pi04( pi048 ), .pi05( pi172 ), .pi06( pi173 ), .pi07( pi174 ), .pi08( pi175 ), .pi09( pi176 ), .pi10( n13 ), .pi11( n14 ), .pi12( n15 ), .pi13( n47 ), .po0( n16 ), .po1( n186 ), .po2( n187 ), .po3( n188 ), .po4( n191 ), .po5( n192 ) );
  max_63 U63 ( .pi00( pi299 ), .pi01( pi300 ), .pi02( pi301 ), .pi03( pi302 ), .pi04( pi427 ), .pi05( pi428 ), .pi06( pi429 ), .pi07( pi430 ), .pi08( n66 ), .pi09( n67 ), .pi10( n97 ), .pi11( n183 ), .pi12( n185 ), .pi13( n186 ), .pi14( n187 ), .pi15( n188 ), .pi16( tpo129 ), .po0( n65 ), .po1( n68 ), .po2( n184 ), .po3( n189 ), .po4( n190 ), .po5( tpo043 ), .po6( tpo044 ), .po7( tpo045 ), .po8( tpo046 ) );
  max_64 U64 ( .pi00( pi303 ), .pi01( pi304 ), .pi02( pi431 ), .pi03( pi432 ), .pi04( n68 ), .pi05( n97 ), .pi06( n189 ), .pi07( n190 ), .pi08( n191 ), .pi09( n192 ), .pi10( n193 ), .pi11( tpo129 ), .po0( n67 ), .po1( n69 ), .po2( n194 ), .po3( tpo047 ), .po4( tpo048 ) );
endmodule
module max_63(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, po0, po1, po2, po3, po4, po5, po6, po7, po8);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8;
  wire n0, n1, n2, n3, n4, n5, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7, tpo8;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = tpo7;
  assign po8 = tpo8;
  max_63_0 U0 ( .pi0( pi00 ), .pi1( pi04 ), .pi2( pi10 ), .pi3( pi11 ), .pi4( pi16 ), .po0(  ), .po1(  ), .po2( tpo0 ), .po3( n0 ), .po4( tpo2 ), .po5( n2 ), .po6( tpo5 ) );
  max_63_1 U1 ( .pi00( pi01 ), .pi01( pi02 ), .pi02( pi03 ), .pi03( pi05 ), .pi04( pi06 ), .pi05( pi07 ), .pi06( pi08 ), .pi07( pi09 ), .pi08( pi10 ), .pi09( n0 ), .po0( tpo1 ), .po1( n1 ), .po2( n3 ), .po3( n4 ), .po4( n5 ) );
  max_63_2 U2 ( .pi00( pi12 ), .pi01( pi13 ), .pi02( pi14 ), .pi03( pi15 ), .pi04( pi16 ), .pi05( n1 ), .pi06( n2 ), .pi07( n3 ), .pi08( n4 ), .pi09( n5 ), .po0( tpo3 ), .po1( tpo4 ), .po2( tpo6 ), .po3( tpo7 ), .po4( tpo8 ) );
endmodule
module max_61(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, po0, po1, po2, po3, po4, po5, po6, po7);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n0, n1, n2, n3, n4, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = tpo7;
  max_61_0 U0 ( .pi0( pi00 ), .pi1( pi04 ), .pi2( pi10 ), .pi3( pi11 ), .pi4( pi17 ), .po0(  ), .po1(  ), .po2( tpo0 ), .po3( n0 ), .po4( tpo2 ), .po5( n1 ), .po6( tpo4 ) );
  max_61_1 U1 ( .pi00( pi01 ), .pi01( pi02 ), .pi02( pi03 ), .pi03( pi05 ), .pi04( pi06 ), .pi05( pi07 ), .pi06( pi08 ), .pi07( pi09 ), .pi08( pi10 ), .pi09( n0 ), .po0( tpo1 ), .po1( n2 ), .po2( n3 ), .po3( n4 ) );
  max_61_2 U2 ( .pi00( pi12 ), .pi01( pi13 ), .pi02( pi14 ), .pi03( pi15 ), .pi04( pi16 ), .pi05( pi17 ), .pi06( n1 ), .pi07( n2 ), .pi08( n3 ), .pi09( n4 ), .po0( tpo3 ), .po1( tpo5 ), .po2( tpo6 ), .po3( tpo7 ) );
endmodule
module max_59(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, po0, po1, po2, po3, po4, po5, po6);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16;
  output po0, po1, po2, po3, po4, po5, po6;
  wire n0, n1, n2, n3, n4, n5, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  max_59_0 U0 ( .pi0( pi10 ), .pi1( pi11 ), .pi2( pi12 ), .pi3( pi16 ), .pi4( n0 ), .po0(  ), .po1( n1 ), .po2( tpo3 ) );
  max_59_1 U1 ( .pi00( pi00 ), .pi01( pi01 ), .pi02( pi02 ), .pi03( pi03 ), .pi04( pi04 ), .pi05( pi05 ), .pi06( pi06 ), .pi07( pi07 ), .pi08( pi08 ), .pi09( pi09 ), .po0( tpo0 ), .po1( n0 ), .po2( n2 ), .po3( n3 ), .po4( n4 ), .po5( n5 ) );
  max_59_2 U2 ( .pi0( pi13 ), .pi1( pi14 ), .pi2( pi15 ), .pi3( pi16 ), .pi4( n1 ), .pi5( n2 ), .pi6( n3 ), .pi7( n4 ), .pi8( n5 ), .po0( tpo1 ), .po1( tpo2 ), .po2( tpo4 ), .po3( tpo5 ), .po4( tpo6 ) );
endmodule
module max_57(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, po0, po1, po2, po3, po4, po5, po6);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20;
  output po0, po1, po2, po3, po4, po5, po6;
  wire n0, n1, n2, n3, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  max_57_0 U0 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi02 ), .pi3( pi03 ), .pi4( pi04 ), .pi5( pi05 ), .pi6( pi12 ), .pi7( pi13 ), .po0( tpo0 ), .po1( tpo2 ), .po2( n1 ), .po3( n2 ) );
  max_57_1 U1 ( .pi0( pi06 ), .pi1( pi07 ), .pi2( pi08 ), .pi3( pi09 ), .pi4( pi10 ), .pi5( pi11 ), .pi6( pi14 ), .pi7( pi15 ), .pi8( pi16 ), .po0( tpo1 ), .po1( tpo3 ), .po2( n0 ), .po3( n3 ) );
  max_57_2 U2 ( .pi00( pi17 ), .pi01( pi18 ), .pi02( pi19 ), .pi03( pi20 ), .pi04( tpo2 ), .pi05( tpo3 ), .pi06( n0 ), .pi07( n1 ), .pi08( n2 ), .pi09( n3 ), .po0( tpo4 ), .po1( tpo5 ), .po2( tpo6 ) );
endmodule
module max_54(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, po0, po1, po2, po3, po4, po5, po6, po7);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n0, n1, n2, n3, n4, n5, n6, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = tpo7;
  max_54_0 U0 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi02 ), .pi3( pi03 ), .pi4( pi04 ), .pi5( pi05 ), .pi6( pi12 ), .pi7( pi13 ), .po0( tpo0 ), .po1( tpo1 ), .po2( n0 ), .po3( n3 ), .po4( n6 ) );
  max_54_1 U1 ( .pi0( pi06 ), .pi1( pi07 ), .pi2( pi08 ), .pi3( pi09 ), .pi4( pi10 ), .pi5( pi11 ), .pi6( pi14 ), .pi7( pi15 ), .po0( tpo2 ), .po1( n1 ), .po2( n2 ), .po3( n4 ), .po4( n5 ) );
  max_54_2 U2 ( .pi00( pi16 ), .pi01( pi17 ), .pi02( pi18 ), .pi03( n0 ), .pi04( n1 ), .pi05( n2 ), .pi06( n3 ), .pi07( n4 ), .pi08( n5 ), .pi09( n6 ), .po0( tpo3 ), .po1( tpo4 ), .po2( tpo5 ), .po3( tpo6 ), .po4( tpo7 ) );
endmodule
module max_52(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, po0, po1, po2, po3, po4, po5, po6);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18;
  output po0, po1, po2, po3, po4, po5, po6;
  wire n0, n1, n2, n3, n4, n5, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  max_52_0 U0 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi05 ), .pi3( pi06 ), .pi4( pi10 ), .pi5( pi11 ), .pi6( n0 ), .po0(  ), .po1( n1 ), .po2( tpo1 ), .po3( n3 ) );
  max_52_1 U1 ( .pi00( pi12 ), .pi01( pi13 ), .pi02( pi14 ), .pi03( pi15 ), .pi04( pi16 ), .pi05( pi17 ), .pi06( pi18 ), .pi07( tpo1 ), .pi08( n2 ), .pi09( n3 ), .pi10( n4 ), .pi11( n5 ), .po0( tpo2 ), .po1( tpo3 ), .po2( tpo4 ), .po3( tpo5 ), .po4( tpo6 ) );
  max_52_2 U2 ( .pi0( pi02 ), .pi1( pi03 ), .pi2( pi04 ), .pi3( pi07 ), .pi4( pi08 ), .pi5( pi09 ), .pi6( pi11 ), .pi7( n1 ), .po0( n0 ), .po1( tpo0 ), .po2( n2 ), .po3( n4 ), .po4( n5 ) );
endmodule
module max_50(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, po0, po1, po2, po3, po4, po5, po6, po7, po8);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8;
  wire n0, n1, n2, n3, n4, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7, tpo8;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = tpo7;
  assign po8 = tpo8;
  max_50_0 U0 ( .pi0( pi13 ), .pi1( pi14 ), .pi2( pi15 ), .pi3( pi16 ), .pi4( pi17 ), .pi5( n2 ), .pi6( n3 ), .pi7( n4 ), .po0( tpo4 ), .po1( tpo5 ), .po2( tpo6 ), .po3( tpo7 ), .po4( tpo8 ) );
  max_50_1 U1 ( .pi00( pi00 ), .pi01( pi01 ), .pi02( pi02 ), .pi03( pi05 ), .pi04( pi06 ), .pi05( pi07 ), .pi06( pi10 ), .pi07( pi11 ), .pi08( pi12 ), .pi09( n0 ), .po0( n1 ), .po1( tpo2 ), .po2( tpo3 ), .po3( n2 ) );
  max_50_2 U2 ( .pi0( pi03 ), .pi1( pi04 ), .pi2( pi08 ), .pi3( pi09 ), .pi4( pi12 ), .pi5( n1 ), .po0(  ), .po1( n0 ), .po2( tpo0 ), .po3( tpo1 ), .po4( n3 ), .po5( n4 ) );
endmodule
module max_48(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, po0, po1, po2, po3, po4, po5, po6, po7, po8);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8;
  wire n0, n1, n2, n3, n4, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7, tpo8;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = tpo7;
  assign po8 = tpo8;
  max_48_0 U0 ( .pi0( pi08 ), .pi1( pi09 ), .pi2( pi14 ), .pi3( pi15 ), .pi4( pi16 ), .pi5( n3 ), .pi6( n4 ), .po0(  ), .po1( tpo3 ), .po2( tpo7 ), .po3( tpo8 ) );
  max_48_1 U1 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi02 ), .pi3( pi03 ), .pi4( pi04 ), .pi5( pi05 ), .pi6( pi06 ), .pi7( pi07 ), .po0( tpo0 ), .po1( tpo1 ), .po2( tpo2 ), .po3( n0 ), .po4( n1 ), .po5( n2 ) );
  max_48_2 U2 ( .pi0( pi10 ), .pi1( pi11 ), .pi2( pi12 ), .pi3( pi13 ), .pi4( pi16 ), .pi5( n0 ), .pi6( n1 ), .pi7( n2 ), .po0( n3 ), .po1( n4 ), .po2( tpo4 ), .po3( tpo5 ), .po4( tpo6 ) );
endmodule
module max_44(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, po0, po1, po2, po3, po4, po5, po6, po7, po8);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8;
  wire n0, n1, n2, n3, n4, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7, tpo8;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = tpo7;
  assign po8 = tpo8;
  max_44_0 U0 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi02 ), .pi3( pi05 ), .pi4( pi06 ), .pi5( pi07 ), .pi6( pi10 ), .pi7( pi11 ), .po0( n0 ), .po1( tpo2 ), .po2( n1 ), .po3( n2 ) );
  max_44_1 U1 ( .pi00( pi12 ), .pi01( pi13 ), .pi02( pi14 ), .pi03( pi15 ), .pi04( pi16 ), .pi05( pi18 ), .pi06( tpo2 ), .pi07( n1 ), .pi08( n2 ), .pi09( n3 ), .pi10( n4 ), .po0( tpo3 ), .po1( tpo5 ), .po2( tpo6 ), .po3( tpo7 ) );
  max_44_2 U2 ( .pi0( pi03 ), .pi1( pi04 ), .pi2( pi08 ), .pi3( pi09 ), .pi4( pi11 ), .pi5( pi17 ), .pi6( pi18 ), .pi7( n0 ), .po0(  ), .po1(  ), .po2( tpo0 ), .po3( tpo1 ), .po4( n3 ), .po5( n4 ), .po6( tpo4 ), .po7( tpo8 ) );
endmodule
module max_42(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, po0, po1, po2, po3, po4, po5, po6, po7);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n0, n1, n2, n3, n4, n5, n6, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = tpo7;
  max_42_0 U0 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi02 ), .pi3( pi03 ), .pi4( pi04 ), .pi5( pi05 ), .pi6( pi12 ), .pi7( pi13 ), .po0( tpo0 ), .po1( tpo1 ), .po2( n0 ), .po3( n2 ), .po4( n4 ) );
  max_42_1 U1 ( .pi0( pi06 ), .pi1( pi07 ), .pi2( pi08 ), .pi3( pi09 ), .pi4( pi10 ), .pi5( pi11 ), .pi6( pi14 ), .pi7( pi15 ), .pi8( pi16 ), .po0( tpo2 ), .po1( n1 ), .po2( n3 ), .po3( n5 ), .po4( n6 ) );
  max_42_2 U2 ( .pi00( pi17 ), .pi01( pi18 ), .pi02( pi19 ), .pi03( n0 ), .pi04( n1 ), .pi05( n2 ), .pi06( n3 ), .pi07( n4 ), .pi08( n5 ), .pi09( n6 ), .po0( tpo3 ), .po1( tpo4 ), .po2( tpo5 ), .po3( tpo6 ), .po4( tpo7 ) );
endmodule
module max_41(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, po0, po1, po2, po3, po4, po5, po6, po7);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n0, n1, n2, n3, n4, n5, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = tpo7;
  max_41_0 U0 ( .pi0( pi03 ), .pi1( pi04 ), .pi2( pi08 ), .pi3( pi09 ), .pi4( pi11 ), .pi5( n0 ), .pi6( n1 ), .po0(  ), .po1( tpo0 ), .po2( tpo2 ), .po3( n2 ) );
  max_41_1 U1 ( .pi00( pi12 ), .pi01( pi13 ), .pi02( pi15 ), .pi03( pi16 ), .pi04( pi17 ), .pi05( pi18 ), .pi06( tpo2 ), .pi07( n2 ), .pi08( n3 ), .pi09( n4 ), .pi10( n5 ), .po0(  ), .po1( tpo3 ), .po2( tpo5 ), .po3( tpo6 ), .po4( tpo7 ) );
  max_41_2 U2 ( .pi00( pi00 ), .pi01( pi01 ), .pi02( pi02 ), .pi03( pi05 ), .pi04( pi06 ), .pi05( pi07 ), .pi06( pi10 ), .pi07( pi11 ), .pi08( pi14 ), .pi09( pi18 ), .po0( n0 ), .po1( n1 ), .po2( tpo1 ), .po3( n3 ), .po4( n4 ), .po5( n5 ), .po6( tpo4 ) );
endmodule
module max_38(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, po0, po1, po2, po3, po4, po5, po6);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16;
  output po0, po1, po2, po3, po4, po5, po6;
  wire n0, n1, n2, n3, n4, n5, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  max_38_0 U0 ( .pi0( pi02 ), .pi1( pi03 ), .pi2( pi06 ), .pi3( pi07 ), .pi4( pi08 ), .pi5( pi09 ), .pi6( n0 ), .pi7( n1 ), .po0(  ), .po1( tpo1 ), .po2( n4 ), .po3( n5 ) );
  max_38_1 U1 ( .pi00( pi10 ), .pi01( pi11 ), .pi02( pi12 ), .pi03( pi13 ), .pi04( pi14 ), .pi05( pi15 ), .pi06( pi16 ), .pi07( n2 ), .pi08( n3 ), .pi09( n4 ), .pi10( n5 ), .po0( tpo2 ), .po1( tpo3 ), .po2( tpo4 ), .po3( tpo5 ), .po4( tpo6 ) );
  max_38_2 U2 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi04 ), .pi3( pi05 ), .pi4( pi09 ), .po0( tpo0 ), .po1( n0 ), .po2( n1 ), .po3( n2 ), .po4( n3 ) );
endmodule
module max_34(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, po0, po1, po2, po3, po4, po5, po6);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18;
  output po0, po1, po2, po3, po4, po5, po6;
  wire n0, n1, n2, n3, n4, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  max_34_0 U0 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi04 ), .pi3( pi05 ), .pi4( pi08 ), .pi5( pi09 ), .po0(  ), .po1( n0 ), .po2( n1 ), .po3( n2 ) );
  max_34_1 U1 ( .pi00( pi02 ), .pi01( pi03 ), .pi02( pi06 ), .pi03( pi07 ), .pi04( pi09 ), .pi05( pi15 ), .pi06( pi16 ), .pi07( pi17 ), .pi08( pi18 ), .pi09( n0 ), .pi10( n4 ), .po0( tpo0 ), .po1( n3 ), .po2( tpo1 ), .po3( tpo5 ), .po4( tpo6 ) );
  max_34_2 U2 ( .pi0( pi10 ), .pi1( pi11 ), .pi2( pi12 ), .pi3( pi13 ), .pi4( pi14 ), .pi5( pi18 ), .pi6( n1 ), .pi7( n2 ), .pi8( n3 ), .po0(  ), .po1( n4 ), .po2( tpo2 ), .po3( tpo3 ), .po4( tpo4 ) );
endmodule
module max_31(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, po0, po1, po2, po3, po4, po5, po6);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16;
  output po0, po1, po2, po3, po4, po5, po6;
  wire n0, n1, n2, n3, n4, n5, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  max_31_0 U0 ( .pi0( pi03 ), .pi1( pi07 ), .pi2( pi09 ), .pi3( pi10 ), .pi4( n0 ), .pi5( n1 ), .po0(  ), .po1( tpo1 ), .po2( n2 ) );
  max_31_1 U1 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi02 ), .pi3( pi04 ), .pi4( pi05 ), .pi5( pi06 ), .pi6( pi08 ), .pi7( pi10 ), .po0( tpo0 ), .po1( n0 ), .po2( n1 ), .po3( n3 ), .po4( n4 ), .po5( n5 ) );
  max_31_2 U2 ( .pi00( pi11 ), .pi01( pi12 ), .pi02( pi13 ), .pi03( pi14 ), .pi04( pi15 ), .pi05( pi16 ), .pi06( n2 ), .pi07( n3 ), .pi08( n4 ), .pi09( n5 ), .po0( tpo2 ), .po1( tpo3 ), .po2( tpo4 ), .po3( tpo5 ), .po4( tpo6 ) );
endmodule
module max_28(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, po0, po1, po2, po3, po4, po5, po6, po7);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n0, n1, n2, n3, n4, n5, n6, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = tpo7;
  max_28_0 U0 ( .pi0( pi00 ), .pi1( pi05 ), .pi2( pi12 ), .pi3( pi13 ), .pi4( pi14 ), .pi5( tpo1 ), .pi6( tpo2 ), .pi7( n4 ), .pi8( tpo3 ), .po0( tpo0 ), .po1( n1 ), .po2( n5 ), .po3( tpo4 ) );
  max_28_1 U1 ( .pi00( pi01 ), .pi01( pi02 ), .pi02( pi06 ), .pi03( pi07 ), .pi04( pi11 ), .pi05( pi15 ), .pi06( n0 ), .pi07( n1 ), .pi08( tpo1 ), .pi09( tpo3 ), .po0( n2 ), .po1( n3 ), .po2( tpo2 ), .po3( n4 ), .po4( n6 ), .po5( tpo5 ) );
  max_28_2 U2 ( .pi00( pi03 ), .pi01( pi04 ), .pi02( pi08 ), .pi03( pi09 ), .pi04( pi10 ), .pi05( pi16 ), .pi06( n2 ), .pi07( n3 ), .pi08( n5 ), .pi09( n6 ), .po0( n0 ), .po1( tpo1 ), .po2( tpo3 ), .po3( tpo6 ), .po4( tpo7 ) );
endmodule
module max_26(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, po0, po1, po2, po3, po4, po5, po6, po7);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n0, n1, n2, n3, n4, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = tpo7;
  max_26_0 U0 ( .pi0( pi03 ), .pi1( pi07 ), .pi2( pi09 ), .pi3( pi15 ), .pi4( pi16 ), .po0(  ), .po1(  ), .po2( n0 ), .po3( tpo1 ), .po4( n4 ), .po5( tpo3 ), .po6( tpo7 ) );
  max_26_1 U1 ( .pi00( pi10 ), .pi01( pi11 ), .pi02( pi12 ), .pi03( pi13 ), .pi04( pi14 ), .pi05( pi16 ), .pi06( n1 ), .pi07( n2 ), .pi08( n3 ), .pi09( n4 ), .po0( tpo2 ), .po1( tpo4 ), .po2( tpo5 ), .po3( tpo6 ) );
  max_26_2 U2 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi02 ), .pi3( pi04 ), .pi4( pi05 ), .pi5( pi06 ), .pi6( pi08 ), .pi7( pi09 ), .pi8( n0 ), .po0( tpo0 ), .po1( n1 ), .po2( n2 ), .po3( n3 ) );
endmodule
module max_24(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, po0, po1, po2, po3, po4, po5, po6);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20;
  output po0, po1, po2, po3, po4, po5, po6;
  wire n0, n1, n2, n3, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  max_24_0 U0 ( .pi0( pi06 ), .pi1( pi07 ), .pi2( pi08 ), .pi3( pi09 ), .pi4( pi10 ), .pi5( pi11 ), .pi6( pi15 ), .pi7( pi16 ), .pi8( pi17 ), .po0( tpo1 ), .po1( tpo3 ), .po2( n0 ), .po3( n3 ) );
  max_24_1 U1 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi02 ), .pi3( pi03 ), .pi4( pi04 ), .pi5( pi05 ), .pi6( pi12 ), .pi7( pi13 ), .pi8( pi14 ), .po0( tpo0 ), .po1( tpo2 ), .po2( n1 ), .po3( n2 ) );
  max_24_2 U2 ( .pi0( pi18 ), .pi1( pi19 ), .pi2( pi20 ), .pi3( tpo2 ), .pi4( tpo3 ), .pi5( n0 ), .pi6( n1 ), .pi7( n2 ), .pi8( n3 ), .po0( tpo4 ), .po1( tpo5 ), .po2( tpo6 ) );
endmodule
module max_23(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, po0, po1, po2, po3, po4, po5, po6);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16;
  output po0, po1, po2, po3, po4, po5, po6;
  wire n0, n1, n2, n3, n4, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  max_23_0 U0 ( .pi0( pi11 ), .pi1( pi12 ), .pi2( pi13 ), .pi3( pi14 ), .pi4( pi16 ), .pi5( n2 ), .pi6( n3 ), .po0(  ), .po1( n4 ), .po2( tpo3 ), .po3( tpo4 ) );
  max_23_1 U1 ( .pi00( pi02 ), .pi01( pi03 ), .pi02( pi06 ), .pi03( pi07 ), .pi04( pi09 ), .pi05( pi10 ), .pi06( pi15 ), .pi07( pi16 ), .pi08( n1 ), .pi09( n4 ), .po0( n0 ), .po1( tpo0 ), .po2( tpo1 ), .po3( tpo2 ), .po4( tpo5 ), .po5( tpo6 ) );
  max_23_2 U2 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi04 ), .pi3( pi05 ), .pi4( pi08 ), .pi5( pi09 ), .pi6( n0 ), .po0(  ), .po1( n1 ), .po2( n2 ), .po3( n3 ) );
endmodule
module max_17(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, po0, po1, po2, po3, po4, po5, po6, po7);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n0, n1, n2, n3, n4, n5, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = tpo7;
  max_17_0 U0 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi05 ), .pi3( pi06 ), .pi4( pi10 ), .pi5( pi11 ), .pi6( n0 ), .po0(  ), .po1( tpo0 ), .po2( n1 ), .po3( tpo2 ), .po4( n3 ) );
  max_17_1 U1 ( .pi00( pi12 ), .pi01( pi13 ), .pi02( pi14 ), .pi03( pi15 ), .pi04( pi16 ), .pi05( pi17 ), .pi06( n2 ), .pi07( n3 ), .pi08( n4 ), .pi09( n5 ), .po0( tpo3 ), .po1( tpo4 ), .po2( tpo5 ), .po3( tpo6 ), .po4( tpo7 ) );
  max_17_2 U2 ( .pi0( pi02 ), .pi1( pi03 ), .pi2( pi04 ), .pi3( pi07 ), .pi4( pi08 ), .pi5( pi09 ), .pi6( pi11 ), .pi7( n1 ), .po0( n0 ), .po1( tpo1 ), .po2( n2 ), .po3( n4 ), .po4( n5 ) );
endmodule
module max_14(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, po0, po1, po2, po3, po4, po5, po6, po7);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n0, n1, n2, n3, n4, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = tpo7;
  max_14_0 U0 ( .pi0( pi00 ), .pi1( pi04 ), .pi2( pi10 ), .pi3( pi11 ), .pi4( pi17 ), .po0(  ), .po1(  ), .po2( tpo0 ), .po3( n0 ), .po4( tpo2 ), .po5( n2 ), .po6( tpo4 ) );
  max_14_1 U1 ( .pi00( pi01 ), .pi01( pi02 ), .pi02( pi03 ), .pi03( pi05 ), .pi04( pi06 ), .pi05( pi07 ), .pi06( pi08 ), .pi07( pi09 ), .pi08( pi10 ), .pi09( n0 ), .po0( tpo1 ), .po1( n1 ), .po2( n3 ), .po3( n4 ) );
  max_14_2 U2 ( .pi00( pi12 ), .pi01( pi13 ), .pi02( pi14 ), .pi03( pi15 ), .pi04( pi16 ), .pi05( pi17 ), .pi06( n1 ), .pi07( n2 ), .pi08( n3 ), .pi09( n4 ), .po0( tpo3 ), .po1( tpo5 ), .po2( tpo6 ), .po3( tpo7 ) );
endmodule
module max_12(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, po0, po1, po2, po3, po4, po5);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16;
  output po0, po1, po2, po3, po4, po5;
  wire n0, n1, n2, n3, n4, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  max_12_0 U0 ( .pi0( pi13 ), .pi1( pi14 ), .pi2( pi15 ), .pi3( pi16 ), .pi4( n2 ), .pi5( n3 ), .pi6( n4 ), .po0(  ), .po1( tpo1 ), .po2( tpo4 ), .po3( tpo5 ) );
  max_12_1 U1 ( .pi0( pi02 ), .pi1( pi03 ), .pi2( pi06 ), .pi3( pi07 ), .pi4( pi09 ), .pi5( n0 ), .pi6( n1 ), .po0(  ), .po1( tpo0 ), .po2( n3 ), .po3( n4 ) );
  max_12_2 U2 ( .pi00( pi00 ), .pi01( pi01 ), .pi02( pi04 ), .pi03( pi05 ), .pi04( pi08 ), .pi05( pi09 ), .pi06( pi10 ), .pi07( pi11 ), .pi08( pi12 ), .pi09( pi16 ), .po0( n0 ), .po1( n1 ), .po2( n2 ), .po3( tpo2 ), .po4( tpo3 ) );
endmodule
module max_6(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, po0, po1, po2, po3, po4, po5, po6, po7);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n0, n1, n2, n3, n4, n5, n6, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = tpo7;
  max_6_0 U0 ( .pi0( pi10 ), .pi1( pi11 ), .pi2( pi16 ), .pi3( pi17 ), .pi4( n4 ), .pi5( n5 ), .pi6( n6 ), .po0(  ), .po1( tpo2 ), .po2( tpo6 ), .po3( tpo7 ) );
  max_6_1 U1 ( .pi0( pi12 ), .pi1( pi13 ), .pi2( pi14 ), .pi3( pi15 ), .pi4( pi17 ), .pi5( n0 ), .pi6( n1 ), .pi7( n2 ), .pi8( n3 ), .po0( tpo1 ), .po1( n4 ), .po2( n5 ), .po3( tpo3 ), .po4( tpo4 ), .po5( tpo5 ) );
  max_6_2 U2 ( .pi00( pi00 ), .pi01( pi01 ), .pi02( pi02 ), .pi03( pi03 ), .pi04( pi04 ), .pi05( pi05 ), .pi06( pi06 ), .pi07( pi07 ), .pi08( pi08 ), .pi09( pi09 ), .po0( tpo0 ), .po1( n0 ), .po2( n1 ), .po3( n2 ), .po4( n3 ), .po5( n6 ) );
endmodule
module max_3(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, po0, po1, po2, po3, po4, po5, po6, po7);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n0, n1, n2, n3, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = tpo7;
  max_3_0 U0 ( .pi0( pi00 ), .pi1( pi07 ), .pi2( pi14 ), .pi3( pi15 ), .pi4( pi17 ), .po0(  ), .po1( n0 ), .po2( tpo1 ) );
  max_3_1 U1 ( .pi0( pi01 ), .pi1( pi02 ), .pi2( pi03 ), .pi3( pi08 ), .pi4( pi09 ), .pi5( pi10 ), .pi6( pi17 ), .pi7( n0 ), .pi8( n1 ), .po0( n2 ), .po1( n3 ), .po2( tpo2 ), .po3( tpo3 ), .po4( tpo4 ) );
  max_3_2 U2 ( .pi00( pi04 ), .pi01( pi05 ), .pi02( pi06 ), .pi03( pi11 ), .pi04( pi12 ), .pi05( pi13 ), .pi06( pi16 ), .pi07( pi17 ), .pi08( n2 ), .pi09( n3 ), .po0( n1 ), .po1( tpo0 ), .po2( tpo5 ), .po3( tpo6 ), .po4( tpo7 ) );
endmodule
module max_1(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, po0, po1, po2, po3, po4, po5, po6);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17;
  output po0, po1, po2, po3, po4, po5, po6;
  wire n0, n1, n2, n3, n4, n5, n6, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  max_1_0 U0 ( .pi0( pi12 ), .pi1( pi14 ), .pi2( pi15 ), .pi3( pi16 ), .pi4( pi17 ), .pi5( n3 ), .pi6( n4 ), .pi7( n5 ), .pi8( n6 ), .po0(  ), .po1( tpo2 ), .po2( tpo5 ), .po3( tpo6 ) );
  max_1_1 U1 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi04 ), .pi3( pi05 ), .pi4( pi10 ), .pi5( pi11 ), .pi6( pi13 ), .pi7( pi17 ), .po0( n0 ), .po1( n1 ), .po2( n2 ), .po3( tpo1 ), .po4( n3 ), .po5( n5 ), .po6( tpo3 ), .po7( tpo4 ) );
  max_1_2 U2 ( .pi00( pi02 ), .pi01( pi03 ), .pi02( pi06 ), .pi03( pi07 ), .pi04( pi08 ), .pi05( pi09 ), .pi06( pi10 ), .pi07( n0 ), .pi08( n1 ), .pi09( n2 ), .po0(  ), .po1( tpo0 ), .po2( n4 ), .po3( n6 ) );
endmodule
