// Benchmark "mult8" written by ABC on Fri Jul  1 13:51:55 2022

module mult8 ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \B[0] ,
    \B[1] , \B[2] , \B[3] , \B[4] , \B[5] , \B[6] , \B[7] ,
    \O[0] , \O[1] , \O[2] , \O[3] , \O[4] , \O[5] , \O[6] , \O[7] , \O[8] ,
    \O[9] , \O[10] , \O[11] , \O[12] , \O[13] , \O[14] , \O[15]   );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \B[0] , \B[1] , \B[2] , \B[3] , \B[4] , \B[5] , \B[6] , \B[7] ;
  output \O[0] , \O[1] , \O[2] , \O[3] , \O[4] , \O[5] , \O[6] , \O[7] ,
    \O[8] , \O[9] , \O[10] , \O[11] , \O[12] , \O[13] , \O[14] , \O[15] ;
  wire new_new_n34__, new_new_n35__, new_new_n36__, new_new_n37__,
    new_new_n39__, new_new_n40__, new_new_n41__, new_new_n42__,
    new_new_n43__, new_new_n44__, new_new_n45__, new_new_n46__,
    new_new_n47__, new_new_n48__, new_new_n49__, new_new_n51__,
    new_new_n52__, new_new_n53__, new_new_n54__, new_new_n55__,
    new_new_n56__, new_new_n57__, new_new_n58__, new_new_n59__,
    new_new_n60__, new_new_n61__, new_new_n62__, new_new_n63__,
    new_new_n64__, new_new_n65__, new_new_n66__, new_new_n67__,
    new_new_n68__, new_new_n69__, new_new_n70__, new_new_n72__,
    new_new_n73__, new_new_n74__, new_new_n75__, new_new_n76__,
    new_new_n77__, new_new_n78__, new_new_n79__, new_new_n80__,
    new_new_n81__, new_new_n82__, new_new_n83__, new_new_n84__,
    new_new_n85__, new_new_n86__, new_new_n87__, new_new_n88__,
    new_new_n89__, new_new_n90__, new_new_n91__, new_new_n92__,
    new_new_n93__, new_new_n94__, new_new_n95__, new_new_n96__,
    new_new_n97__, new_new_n98__, new_new_n99__, new_new_n100__,
    new_new_n102__, new_new_n103__, new_new_n104__, new_new_n105__,
    new_new_n106__, new_new_n107__, new_new_n108__, new_new_n109__,
    new_new_n110__, new_new_n111__, new_new_n112__, new_new_n113__,
    new_new_n114__, new_new_n115__, new_new_n116__, new_new_n117__,
    new_new_n118__, new_new_n119__, new_new_n120__, new_new_n121__,
    new_new_n122__, new_new_n123__, new_new_n124__, new_new_n125__,
    new_new_n126__, new_new_n127__, new_new_n128__, new_new_n129__,
    new_new_n130__, new_new_n131__, new_new_n132__, new_new_n133__,
    new_new_n134__, new_new_n135__, new_new_n136__, new_new_n137__,
    new_new_n138__, new_new_n139__, new_new_n141__, new_new_n142__,
    new_new_n143__, new_new_n144__, new_new_n145__, new_new_n146__,
    new_new_n147__, new_new_n148__, new_new_n149__, new_new_n150__,
    new_new_n151__, new_new_n152__, new_new_n153__, new_new_n154__,
    new_new_n155__, new_new_n156__, new_new_n157__, new_new_n158__,
    new_new_n159__, new_new_n160__, new_new_n161__, new_new_n162__,
    new_new_n163__, new_new_n164__, new_new_n165__, new_new_n166__,
    new_new_n167__, new_new_n168__, new_new_n169__, new_new_n170__,
    new_new_n171__, new_new_n172__, new_new_n173__, new_new_n174__,
    new_new_n175__, new_new_n176__, new_new_n177__, new_new_n178__,
    new_new_n179__, new_new_n180__, new_new_n181__, new_new_n182__,
    new_new_n183__, new_new_n184__, new_new_n185__, new_new_n186__,
    new_new_n187__, new_new_n189__, new_new_n190__, new_new_n191__,
    new_new_n192__, new_new_n193__, new_new_n194__, new_new_n195__,
    new_new_n196__, new_new_n197__, new_new_n198__, new_new_n199__,
    new_new_n200__, new_new_n201__, new_new_n202__, new_new_n203__,
    new_new_n204__, new_new_n205__, new_new_n206__, new_new_n207__,
    new_new_n208__, new_new_n209__, new_new_n210__, new_new_n211__,
    new_new_n212__, new_new_n213__, new_new_n214__, new_new_n215__,
    new_new_n216__, new_new_n217__, new_new_n218__, new_new_n219__,
    new_new_n220__, new_new_n221__, new_new_n222__, new_new_n223__,
    new_new_n224__, new_new_n225__, new_new_n226__, new_new_n227__,
    new_new_n228__, new_new_n229__, new_new_n230__, new_new_n231__,
    new_new_n232__, new_new_n233__, new_new_n234__, new_new_n235__,
    new_new_n236__, new_new_n237__, new_new_n238__, new_new_n239__,
    new_new_n240__, new_new_n241__, new_new_n242__, new_new_n243__,
    new_new_n244__, new_new_n246__, new_new_n247__, new_new_n248__,
    new_new_n249__, new_new_n250__, new_new_n251__, new_new_n252__,
    new_new_n253__, new_new_n254__, new_new_n255__, new_new_n256__,
    new_new_n257__, new_new_n258__, new_new_n259__, new_new_n260__,
    new_new_n261__, new_new_n262__, new_new_n263__, new_new_n264__,
    new_new_n265__, new_new_n266__, new_new_n267__, new_new_n268__,
    new_new_n269__, new_new_n270__, new_new_n271__, new_new_n272__,
    new_new_n273__, new_new_n274__, new_new_n275__, new_new_n276__,
    new_new_n277__, new_new_n278__, new_new_n279__, new_new_n280__,
    new_new_n281__, new_new_n282__, new_new_n283__, new_new_n284__,
    new_new_n285__, new_new_n286__, new_new_n287__, new_new_n288__,
    new_new_n289__, new_new_n290__, new_new_n291__, new_new_n292__,
    new_new_n293__, new_new_n294__, new_new_n295__, new_new_n296__,
    new_new_n297__, new_new_n298__, new_new_n299__, new_new_n300__,
    new_new_n301__, new_new_n302__, new_new_n304__, new_new_n305__,
    new_new_n306__, new_new_n307__, new_new_n308__, new_new_n309__,
    new_new_n310__, new_new_n311__, new_new_n312__, new_new_n313__,
    new_new_n314__, new_new_n315__, new_new_n316__, new_new_n317__,
    new_new_n318__, new_new_n319__, new_new_n320__, new_new_n321__,
    new_new_n322__, new_new_n323__, new_new_n324__, new_new_n325__,
    new_new_n326__, new_new_n327__, new_new_n328__, new_new_n329__,
    new_new_n330__, new_new_n331__, new_new_n332__, new_new_n333__,
    new_new_n334__, new_new_n335__, new_new_n336__, new_new_n337__,
    new_new_n338__, new_new_n339__, new_new_n340__, new_new_n341__,
    new_new_n342__, new_new_n343__, new_new_n344__, new_new_n345__,
    new_new_n346__, new_new_n347__, new_new_n348__, new_new_n349__,
    new_new_n350__, new_new_n351__, new_new_n352__, new_new_n353__,
    new_new_n354__, new_new_n356__, new_new_n357__, new_new_n358__,
    new_new_n359__, new_new_n360__, new_new_n361__, new_new_n362__,
    new_new_n363__, new_new_n364__, new_new_n365__, new_new_n366__,
    new_new_n367__, new_new_n368__, new_new_n369__, new_new_n370__,
    new_new_n371__, new_new_n372__, new_new_n373__, new_new_n374__,
    new_new_n375__, new_new_n376__, new_new_n377__, new_new_n378__,
    new_new_n379__, new_new_n380__, new_new_n381__, new_new_n382__,
    new_new_n383__, new_new_n384__, new_new_n385__, new_new_n386__,
    new_new_n387__, new_new_n388__, new_new_n389__, new_new_n390__,
    new_new_n391__, new_new_n392__, new_new_n393__, new_new_n394__,
    new_new_n395__, new_new_n396__, new_new_n397__, new_new_n398__,
    new_new_n399__, new_new_n400__, new_new_n401__, new_new_n403__,
    new_new_n404__, new_new_n405__, new_new_n406__, new_new_n407__,
    new_new_n408__, new_new_n409__, new_new_n410__, new_new_n411__,
    new_new_n412__, new_new_n413__, new_new_n414__, new_new_n415__,
    new_new_n416__, new_new_n417__, new_new_n418__, new_new_n419__,
    new_new_n420__, new_new_n421__, new_new_n422__, new_new_n423__,
    new_new_n424__, new_new_n425__, new_new_n426__, new_new_n427__,
    new_new_n428__, new_new_n429__, new_new_n430__, new_new_n431__,
    new_new_n432__, new_new_n433__, new_new_n434__, new_new_n435__,
    new_new_n436__, new_new_n437__, new_new_n438__, new_new_n439__,
    new_new_n441__, new_new_n442__, new_new_n443__, new_new_n444__,
    new_new_n445__, new_new_n446__, new_new_n447__, new_new_n448__,
    new_new_n449__, new_new_n450__, new_new_n451__, new_new_n452__,
    new_new_n453__, new_new_n454__, new_new_n455__, new_new_n456__,
    new_new_n457__, new_new_n458__, new_new_n459__, new_new_n460__,
    new_new_n461__, new_new_n462__, new_new_n463__, new_new_n464__,
    new_new_n465__, new_new_n466__, new_new_n467__, new_new_n468__,
    new_new_n470__, new_new_n471__, new_new_n472__, new_new_n473__,
    new_new_n474__, new_new_n475__, new_new_n476__, new_new_n477__,
    new_new_n478__, new_new_n479__, new_new_n480__, new_new_n481__,
    new_new_n482__, new_new_n483__, new_new_n484__, new_new_n485__,
    new_new_n486__, new_new_n487__, new_new_n488__, new_new_n490__,
    new_new_n491__, new_new_n492__, new_new_n493__, new_new_n494__,
    new_new_n495__, new_new_n496__, new_new_n497__, new_new_n498__,
    new_new_n499__, new_new_n501__;
  assign \O[0]  = \A[0]  & \B[0] ;
  assign new_new_n34__ = \A[0]  & \B[1] ;
  assign new_new_n35__ = \A[1]  & \B[0] ;
  assign new_new_n36__ = ~new_new_n34__ & ~new_new_n35__;
  assign new_new_n37__ = new_new_n34__ & new_new_n35__;
  assign \O[1]  = ~new_new_n36__ & ~new_new_n37__;
  assign new_new_n39__ = \A[0]  & \B[2] ;
  assign new_new_n40__ = \A[1]  & \B[1] ;
  assign new_new_n41__ = \A[2]  & \B[0] ;
  assign new_new_n42__ = ~new_new_n40__ & ~new_new_n41__;
  assign new_new_n43__ = new_new_n40__ & new_new_n41__;
  assign new_new_n44__ = ~new_new_n42__ & ~new_new_n43__;
  assign new_new_n45__ = ~new_new_n37__ & ~new_new_n44__;
  assign new_new_n46__ = new_new_n37__ & ~new_new_n43__;
  assign new_new_n47__ = ~new_new_n45__ & ~new_new_n46__;
  assign new_new_n48__ = new_new_n39__ & ~new_new_n47__;
  assign new_new_n49__ = ~new_new_n39__ & new_new_n47__;
  assign \O[2]  = new_new_n48__ | new_new_n49__;
  assign new_new_n51__ = \A[0]  & \B[3] ;
  assign new_new_n52__ = new_new_n39__ & ~new_new_n45__;
  assign new_new_n53__ = ~new_new_n46__ & ~new_new_n52__;
  assign new_new_n54__ = \A[1]  & \B[2] ;
  assign new_new_n55__ = \A[2]  & \B[1] ;
  assign new_new_n56__ = \A[3]  & \B[0] ;
  assign new_new_n57__ = ~new_new_n55__ & ~new_new_n56__;
  assign new_new_n58__ = new_new_n55__ & new_new_n56__;
  assign new_new_n59__ = ~new_new_n57__ & ~new_new_n58__;
  assign new_new_n60__ = ~new_new_n43__ & ~new_new_n59__;
  assign new_new_n61__ = new_new_n43__ & ~new_new_n58__;
  assign new_new_n62__ = ~new_new_n60__ & ~new_new_n61__;
  assign new_new_n63__ = new_new_n54__ & ~new_new_n62__;
  assign new_new_n64__ = ~new_new_n54__ & new_new_n62__;
  assign new_new_n65__ = ~new_new_n63__ & ~new_new_n64__;
  assign new_new_n66__ = ~new_new_n53__ & ~new_new_n65__;
  assign new_new_n67__ = new_new_n53__ & new_new_n65__;
  assign new_new_n68__ = ~new_new_n66__ & ~new_new_n67__;
  assign new_new_n69__ = new_new_n51__ & ~new_new_n68__;
  assign new_new_n70__ = ~new_new_n51__ & new_new_n68__;
  assign \O[3]  = new_new_n69__ | new_new_n70__;
  assign new_new_n72__ = \A[0]  & \B[4] ;
  assign new_new_n73__ = new_new_n51__ & ~new_new_n67__;
  assign new_new_n74__ = ~new_new_n66__ & ~new_new_n73__;
  assign new_new_n75__ = \A[1]  & \B[3] ;
  assign new_new_n76__ = new_new_n54__ & ~new_new_n60__;
  assign new_new_n77__ = ~new_new_n61__ & ~new_new_n76__;
  assign new_new_n78__ = \A[2]  & \B[2] ;
  assign new_new_n79__ = \A[3]  & \B[1] ;
  assign new_new_n80__ = \A[4]  & \B[0] ;
  assign new_new_n81__ = ~new_new_n79__ & ~new_new_n80__;
  assign new_new_n82__ = new_new_n79__ & new_new_n80__;
  assign new_new_n83__ = ~new_new_n81__ & ~new_new_n82__;
  assign new_new_n84__ = ~new_new_n58__ & ~new_new_n83__;
  assign new_new_n85__ = new_new_n58__ & ~new_new_n82__;
  assign new_new_n86__ = ~new_new_n84__ & ~new_new_n85__;
  assign new_new_n87__ = new_new_n78__ & ~new_new_n86__;
  assign new_new_n88__ = ~new_new_n78__ & new_new_n86__;
  assign new_new_n89__ = ~new_new_n87__ & ~new_new_n88__;
  assign new_new_n90__ = ~new_new_n77__ & ~new_new_n89__;
  assign new_new_n91__ = new_new_n77__ & new_new_n89__;
  assign new_new_n92__ = ~new_new_n90__ & ~new_new_n91__;
  assign new_new_n93__ = new_new_n75__ & ~new_new_n92__;
  assign new_new_n94__ = ~new_new_n75__ & new_new_n92__;
  assign new_new_n95__ = ~new_new_n93__ & ~new_new_n94__;
  assign new_new_n96__ = ~new_new_n74__ & ~new_new_n95__;
  assign new_new_n97__ = new_new_n74__ & new_new_n95__;
  assign new_new_n98__ = ~new_new_n96__ & ~new_new_n97__;
  assign new_new_n99__ = new_new_n72__ & new_new_n98__;
  assign new_new_n100__ = ~new_new_n72__ & ~new_new_n98__;
  assign \O[4]  = ~new_new_n99__ & ~new_new_n100__;
  assign new_new_n102__ = \A[0]  & \B[5] ;
  assign new_new_n103__ = new_new_n72__ & ~new_new_n97__;
  assign new_new_n104__ = ~new_new_n96__ & ~new_new_n103__;
  assign new_new_n105__ = \A[1]  & \B[4] ;
  assign new_new_n106__ = new_new_n75__ & ~new_new_n91__;
  assign new_new_n107__ = ~new_new_n90__ & ~new_new_n106__;
  assign new_new_n108__ = \A[2]  & \B[3] ;
  assign new_new_n109__ = new_new_n78__ & ~new_new_n84__;
  assign new_new_n110__ = ~new_new_n85__ & ~new_new_n109__;
  assign new_new_n111__ = \A[3]  & \B[2] ;
  assign new_new_n112__ = \A[4]  & \B[1] ;
  assign new_new_n113__ = \A[5]  & \B[0] ;
  assign new_new_n114__ = ~new_new_n112__ & ~new_new_n113__;
  assign new_new_n115__ = new_new_n112__ & new_new_n113__;
  assign new_new_n116__ = ~new_new_n114__ & ~new_new_n115__;
  assign new_new_n117__ = ~new_new_n82__ & ~new_new_n116__;
  assign new_new_n118__ = new_new_n82__ & ~new_new_n115__;
  assign new_new_n119__ = ~new_new_n117__ & ~new_new_n118__;
  assign new_new_n120__ = new_new_n111__ & ~new_new_n119__;
  assign new_new_n121__ = ~new_new_n111__ & new_new_n119__;
  assign new_new_n122__ = ~new_new_n120__ & ~new_new_n121__;
  assign new_new_n123__ = ~new_new_n110__ & ~new_new_n122__;
  assign new_new_n124__ = new_new_n110__ & new_new_n122__;
  assign new_new_n125__ = ~new_new_n123__ & ~new_new_n124__;
  assign new_new_n126__ = new_new_n108__ & ~new_new_n125__;
  assign new_new_n127__ = ~new_new_n108__ & new_new_n125__;
  assign new_new_n128__ = ~new_new_n126__ & ~new_new_n127__;
  assign new_new_n129__ = ~new_new_n107__ & ~new_new_n128__;
  assign new_new_n130__ = new_new_n107__ & new_new_n128__;
  assign new_new_n131__ = ~new_new_n129__ & ~new_new_n130__;
  assign new_new_n132__ = new_new_n105__ & new_new_n131__;
  assign new_new_n133__ = ~new_new_n105__ & ~new_new_n131__;
  assign new_new_n134__ = ~new_new_n132__ & ~new_new_n133__;
  assign new_new_n135__ = ~new_new_n104__ & new_new_n134__;
  assign new_new_n136__ = new_new_n104__ & ~new_new_n134__;
  assign new_new_n137__ = ~new_new_n135__ & ~new_new_n136__;
  assign new_new_n138__ = new_new_n102__ & ~new_new_n137__;
  assign new_new_n139__ = ~new_new_n102__ & new_new_n137__;
  assign \O[5]  = new_new_n138__ | new_new_n139__;
  assign new_new_n141__ = \A[0]  & \B[6] ;
  assign new_new_n142__ = new_new_n102__ & ~new_new_n136__;
  assign new_new_n143__ = ~new_new_n135__ & ~new_new_n142__;
  assign new_new_n144__ = \A[1]  & \B[5] ;
  assign new_new_n145__ = new_new_n105__ & ~new_new_n130__;
  assign new_new_n146__ = ~new_new_n129__ & ~new_new_n145__;
  assign new_new_n147__ = \A[2]  & \B[4] ;
  assign new_new_n148__ = new_new_n108__ & ~new_new_n124__;
  assign new_new_n149__ = ~new_new_n123__ & ~new_new_n148__;
  assign new_new_n150__ = \A[3]  & \B[3] ;
  assign new_new_n151__ = new_new_n111__ & ~new_new_n117__;
  assign new_new_n152__ = ~new_new_n118__ & ~new_new_n151__;
  assign new_new_n153__ = \A[4]  & \B[2] ;
  assign new_new_n154__ = \A[5]  & \B[1] ;
  assign new_new_n155__ = \A[6]  & \B[0] ;
  assign new_new_n156__ = ~new_new_n154__ & ~new_new_n155__;
  assign new_new_n157__ = new_new_n154__ & new_new_n155__;
  assign new_new_n158__ = ~new_new_n156__ & ~new_new_n157__;
  assign new_new_n159__ = ~new_new_n115__ & ~new_new_n158__;
  assign new_new_n160__ = new_new_n115__ & ~new_new_n157__;
  assign new_new_n161__ = ~new_new_n159__ & ~new_new_n160__;
  assign new_new_n162__ = new_new_n153__ & ~new_new_n161__;
  assign new_new_n163__ = ~new_new_n153__ & new_new_n161__;
  assign new_new_n164__ = ~new_new_n162__ & ~new_new_n163__;
  assign new_new_n165__ = ~new_new_n152__ & ~new_new_n164__;
  assign new_new_n166__ = new_new_n152__ & new_new_n164__;
  assign new_new_n167__ = ~new_new_n165__ & ~new_new_n166__;
  assign new_new_n168__ = new_new_n150__ & ~new_new_n167__;
  assign new_new_n169__ = ~new_new_n150__ & new_new_n167__;
  assign new_new_n170__ = ~new_new_n168__ & ~new_new_n169__;
  assign new_new_n171__ = ~new_new_n149__ & ~new_new_n170__;
  assign new_new_n172__ = new_new_n149__ & new_new_n170__;
  assign new_new_n173__ = ~new_new_n171__ & ~new_new_n172__;
  assign new_new_n174__ = new_new_n147__ & new_new_n173__;
  assign new_new_n175__ = ~new_new_n147__ & ~new_new_n173__;
  assign new_new_n176__ = ~new_new_n174__ & ~new_new_n175__;
  assign new_new_n177__ = ~new_new_n146__ & new_new_n176__;
  assign new_new_n178__ = new_new_n146__ & ~new_new_n176__;
  assign new_new_n179__ = ~new_new_n177__ & ~new_new_n178__;
  assign new_new_n180__ = new_new_n144__ & ~new_new_n179__;
  assign new_new_n181__ = ~new_new_n144__ & new_new_n179__;
  assign new_new_n182__ = ~new_new_n180__ & ~new_new_n181__;
  assign new_new_n183__ = ~new_new_n143__ & ~new_new_n182__;
  assign new_new_n184__ = new_new_n143__ & new_new_n182__;
  assign new_new_n185__ = ~new_new_n183__ & ~new_new_n184__;
  assign new_new_n186__ = new_new_n141__ & new_new_n185__;
  assign new_new_n187__ = ~new_new_n141__ & ~new_new_n185__;
  assign \O[6]  = ~new_new_n186__ & ~new_new_n187__;
  assign new_new_n189__ = \A[0]  & \B[7] ;
  assign new_new_n190__ = new_new_n141__ & ~new_new_n184__;
  assign new_new_n191__ = ~new_new_n183__ & ~new_new_n190__;
  assign new_new_n192__ = \A[1]  & \B[6] ;
  assign new_new_n193__ = new_new_n144__ & ~new_new_n178__;
  assign new_new_n194__ = ~new_new_n177__ & ~new_new_n193__;
  assign new_new_n195__ = \A[2]  & \B[5] ;
  assign new_new_n196__ = new_new_n147__ & ~new_new_n172__;
  assign new_new_n197__ = ~new_new_n171__ & ~new_new_n196__;
  assign new_new_n198__ = \A[3]  & \B[4] ;
  assign new_new_n199__ = new_new_n150__ & ~new_new_n166__;
  assign new_new_n200__ = ~new_new_n165__ & ~new_new_n199__;
  assign new_new_n201__ = \A[4]  & \B[3] ;
  assign new_new_n202__ = new_new_n153__ & ~new_new_n159__;
  assign new_new_n203__ = ~new_new_n160__ & ~new_new_n202__;
  assign new_new_n204__ = \A[5]  & \B[2] ;
  assign new_new_n205__ = \A[6]  & \B[1] ;
  assign new_new_n206__ = \A[7]  & \B[0] ;
  assign new_new_n207__ = ~new_new_n205__ & ~new_new_n206__;
  assign new_new_n208__ = new_new_n205__ & new_new_n206__;
  assign new_new_n209__ = ~new_new_n207__ & ~new_new_n208__;
  assign new_new_n210__ = ~new_new_n157__ & ~new_new_n209__;
  assign new_new_n211__ = new_new_n157__ & ~new_new_n208__;
  assign new_new_n212__ = ~new_new_n210__ & ~new_new_n211__;
  assign new_new_n213__ = new_new_n204__ & ~new_new_n212__;
  assign new_new_n214__ = ~new_new_n204__ & new_new_n212__;
  assign new_new_n215__ = ~new_new_n213__ & ~new_new_n214__;
  assign new_new_n216__ = ~new_new_n203__ & ~new_new_n215__;
  assign new_new_n217__ = new_new_n203__ & new_new_n215__;
  assign new_new_n218__ = ~new_new_n216__ & ~new_new_n217__;
  assign new_new_n219__ = new_new_n201__ & ~new_new_n218__;
  assign new_new_n220__ = ~new_new_n201__ & new_new_n218__;
  assign new_new_n221__ = ~new_new_n219__ & ~new_new_n220__;
  assign new_new_n222__ = ~new_new_n200__ & ~new_new_n221__;
  assign new_new_n223__ = new_new_n200__ & new_new_n221__;
  assign new_new_n224__ = ~new_new_n222__ & ~new_new_n223__;
  assign new_new_n225__ = new_new_n198__ & new_new_n224__;
  assign new_new_n226__ = ~new_new_n198__ & ~new_new_n224__;
  assign new_new_n227__ = ~new_new_n225__ & ~new_new_n226__;
  assign new_new_n228__ = ~new_new_n197__ & new_new_n227__;
  assign new_new_n229__ = new_new_n197__ & ~new_new_n227__;
  assign new_new_n230__ = ~new_new_n228__ & ~new_new_n229__;
  assign new_new_n231__ = new_new_n195__ & ~new_new_n230__;
  assign new_new_n232__ = ~new_new_n195__ & new_new_n230__;
  assign new_new_n233__ = ~new_new_n231__ & ~new_new_n232__;
  assign new_new_n234__ = ~new_new_n194__ & ~new_new_n233__;
  assign new_new_n235__ = new_new_n194__ & new_new_n233__;
  assign new_new_n236__ = ~new_new_n234__ & ~new_new_n235__;
  assign new_new_n237__ = new_new_n192__ & new_new_n236__;
  assign new_new_n238__ = ~new_new_n192__ & ~new_new_n236__;
  assign new_new_n239__ = ~new_new_n237__ & ~new_new_n238__;
  assign new_new_n240__ = ~new_new_n191__ & new_new_n239__;
  assign new_new_n241__ = new_new_n191__ & ~new_new_n239__;
  assign new_new_n242__ = ~new_new_n240__ & ~new_new_n241__;
  assign new_new_n243__ = new_new_n189__ & ~new_new_n242__;
  assign new_new_n244__ = ~new_new_n189__ & new_new_n242__;
  assign \O[7]  = new_new_n243__ | new_new_n244__;
  assign new_new_n246__ = new_new_n189__ & ~new_new_n241__;
  assign new_new_n247__ = ~new_new_n240__ & ~new_new_n246__;
  assign new_new_n248__ = \A[1]  & \B[7] ;
  assign new_new_n249__ = new_new_n192__ & ~new_new_n235__;
  assign new_new_n250__ = ~new_new_n234__ & ~new_new_n249__;
  assign new_new_n251__ = \A[2]  & \B[6] ;
  assign new_new_n252__ = new_new_n195__ & ~new_new_n229__;
  assign new_new_n253__ = ~new_new_n228__ & ~new_new_n252__;
  assign new_new_n254__ = \A[3]  & \B[5] ;
  assign new_new_n255__ = new_new_n198__ & ~new_new_n223__;
  assign new_new_n256__ = ~new_new_n222__ & ~new_new_n255__;
  assign new_new_n257__ = \A[4]  & \B[4] ;
  assign new_new_n258__ = new_new_n201__ & ~new_new_n217__;
  assign new_new_n259__ = ~new_new_n216__ & ~new_new_n258__;
  assign new_new_n260__ = \A[5]  & \B[3] ;
  assign new_new_n261__ = \A[7]  & \B[1] ;
  assign new_new_n262__ = \A[6]  & \B[2] ;
  assign new_new_n263__ = ~new_new_n261__ & ~new_new_n262__;
  assign new_new_n264__ = new_new_n261__ & new_new_n262__;
  assign new_new_n265__ = ~new_new_n208__ & ~new_new_n264__;
  assign new_new_n266__ = ~new_new_n263__ & new_new_n265__;
  assign new_new_n267__ = new_new_n208__ & new_new_n264__;
  assign new_new_n268__ = ~new_new_n266__ & ~new_new_n267__;
  assign new_new_n269__ = new_new_n204__ & ~new_new_n210__;
  assign new_new_n270__ = ~new_new_n211__ & ~new_new_n269__;
  assign new_new_n271__ = ~new_new_n268__ & ~new_new_n270__;
  assign new_new_n272__ = new_new_n268__ & new_new_n270__;
  assign new_new_n273__ = ~new_new_n271__ & ~new_new_n272__;
  assign new_new_n274__ = new_new_n260__ & ~new_new_n273__;
  assign new_new_n275__ = ~new_new_n260__ & new_new_n273__;
  assign new_new_n276__ = ~new_new_n274__ & ~new_new_n275__;
  assign new_new_n277__ = ~new_new_n259__ & ~new_new_n276__;
  assign new_new_n278__ = new_new_n259__ & new_new_n276__;
  assign new_new_n279__ = ~new_new_n277__ & ~new_new_n278__;
  assign new_new_n280__ = new_new_n257__ & new_new_n279__;
  assign new_new_n281__ = ~new_new_n257__ & ~new_new_n279__;
  assign new_new_n282__ = ~new_new_n280__ & ~new_new_n281__;
  assign new_new_n283__ = ~new_new_n256__ & new_new_n282__;
  assign new_new_n284__ = new_new_n256__ & ~new_new_n282__;
  assign new_new_n285__ = ~new_new_n283__ & ~new_new_n284__;
  assign new_new_n286__ = new_new_n254__ & ~new_new_n285__;
  assign new_new_n287__ = ~new_new_n254__ & new_new_n285__;
  assign new_new_n288__ = ~new_new_n286__ & ~new_new_n287__;
  assign new_new_n289__ = ~new_new_n253__ & ~new_new_n288__;
  assign new_new_n290__ = new_new_n253__ & new_new_n288__;
  assign new_new_n291__ = ~new_new_n289__ & ~new_new_n290__;
  assign new_new_n292__ = new_new_n251__ & new_new_n291__;
  assign new_new_n293__ = ~new_new_n251__ & ~new_new_n291__;
  assign new_new_n294__ = ~new_new_n292__ & ~new_new_n293__;
  assign new_new_n295__ = ~new_new_n250__ & new_new_n294__;
  assign new_new_n296__ = new_new_n250__ & ~new_new_n294__;
  assign new_new_n297__ = ~new_new_n295__ & ~new_new_n296__;
  assign new_new_n298__ = new_new_n248__ & ~new_new_n297__;
  assign new_new_n299__ = ~new_new_n248__ & new_new_n297__;
  assign new_new_n300__ = ~new_new_n298__ & ~new_new_n299__;
  assign new_new_n301__ = ~new_new_n247__ & ~new_new_n300__;
  assign new_new_n302__ = new_new_n247__ & new_new_n300__;
  assign \O[8]  = ~new_new_n301__ & ~new_new_n302__;
  assign new_new_n304__ = \A[2]  & \B[7] ;
  assign new_new_n305__ = new_new_n251__ & ~new_new_n290__;
  assign new_new_n306__ = ~new_new_n289__ & ~new_new_n305__;
  assign new_new_n307__ = \A[3]  & \B[6] ;
  assign new_new_n308__ = new_new_n254__ & ~new_new_n284__;
  assign new_new_n309__ = ~new_new_n283__ & ~new_new_n308__;
  assign new_new_n310__ = \A[4]  & \B[5] ;
  assign new_new_n311__ = new_new_n257__ & ~new_new_n278__;
  assign new_new_n312__ = ~new_new_n277__ & ~new_new_n311__;
  assign new_new_n313__ = \A[5]  & \B[4] ;
  assign new_new_n314__ = \A[6]  & \B[3] ;
  assign new_new_n315__ = \A[7]  & \B[2] ;
  assign new_new_n316__ = ~new_new_n265__ & new_new_n315__;
  assign new_new_n317__ = ~new_new_n208__ & ~new_new_n315__;
  assign new_new_n318__ = ~new_new_n316__ & ~new_new_n317__;
  assign new_new_n319__ = new_new_n314__ & ~new_new_n318__;
  assign new_new_n320__ = ~new_new_n314__ & new_new_n318__;
  assign new_new_n321__ = ~new_new_n319__ & ~new_new_n320__;
  assign new_new_n322__ = new_new_n260__ & ~new_new_n272__;
  assign new_new_n323__ = ~new_new_n271__ & ~new_new_n322__;
  assign new_new_n324__ = ~new_new_n321__ & ~new_new_n323__;
  assign new_new_n325__ = new_new_n321__ & new_new_n323__;
  assign new_new_n326__ = ~new_new_n324__ & ~new_new_n325__;
  assign new_new_n327__ = new_new_n313__ & ~new_new_n326__;
  assign new_new_n328__ = ~new_new_n313__ & new_new_n326__;
  assign new_new_n329__ = ~new_new_n327__ & ~new_new_n328__;
  assign new_new_n330__ = ~new_new_n312__ & ~new_new_n329__;
  assign new_new_n331__ = new_new_n312__ & new_new_n329__;
  assign new_new_n332__ = ~new_new_n330__ & ~new_new_n331__;
  assign new_new_n333__ = new_new_n310__ & new_new_n332__;
  assign new_new_n334__ = ~new_new_n310__ & ~new_new_n332__;
  assign new_new_n335__ = ~new_new_n333__ & ~new_new_n334__;
  assign new_new_n336__ = ~new_new_n309__ & new_new_n335__;
  assign new_new_n337__ = new_new_n309__ & ~new_new_n335__;
  assign new_new_n338__ = ~new_new_n336__ & ~new_new_n337__;
  assign new_new_n339__ = new_new_n307__ & ~new_new_n338__;
  assign new_new_n340__ = ~new_new_n307__ & new_new_n338__;
  assign new_new_n341__ = ~new_new_n339__ & ~new_new_n340__;
  assign new_new_n342__ = ~new_new_n306__ & ~new_new_n341__;
  assign new_new_n343__ = new_new_n306__ & new_new_n341__;
  assign new_new_n344__ = ~new_new_n342__ & ~new_new_n343__;
  assign new_new_n345__ = new_new_n304__ & new_new_n344__;
  assign new_new_n346__ = ~new_new_n304__ & ~new_new_n344__;
  assign new_new_n347__ = ~new_new_n345__ & ~new_new_n346__;
  assign new_new_n348__ = new_new_n301__ & new_new_n347__;
  assign new_new_n349__ = ~new_new_n301__ & ~new_new_n347__;
  assign new_new_n350__ = ~new_new_n348__ & ~new_new_n349__;
  assign new_new_n351__ = new_new_n248__ & ~new_new_n296__;
  assign new_new_n352__ = ~new_new_n295__ & ~new_new_n351__;
  assign new_new_n353__ = new_new_n350__ & ~new_new_n352__;
  assign new_new_n354__ = ~new_new_n350__ & new_new_n352__;
  assign \O[9]  = ~new_new_n353__ & ~new_new_n354__;
  assign new_new_n356__ = ~new_new_n349__ & ~new_new_n352__;
  assign new_new_n357__ = ~new_new_n348__ & ~new_new_n356__;
  assign new_new_n358__ = \A[3]  & \B[7] ;
  assign new_new_n359__ = new_new_n307__ & ~new_new_n337__;
  assign new_new_n360__ = ~new_new_n336__ & ~new_new_n359__;
  assign new_new_n361__ = \A[4]  & \B[6] ;
  assign new_new_n362__ = new_new_n310__ & ~new_new_n331__;
  assign new_new_n363__ = ~new_new_n330__ & ~new_new_n362__;
  assign new_new_n364__ = \A[5]  & \B[5] ;
  assign new_new_n365__ = new_new_n313__ & ~new_new_n325__;
  assign new_new_n366__ = ~new_new_n324__ & ~new_new_n365__;
  assign new_new_n367__ = \A[6]  & \B[4] ;
  assign new_new_n368__ = \A[7]  & \B[3] ;
  assign new_new_n369__ = new_new_n314__ & ~new_new_n317__;
  assign new_new_n370__ = ~new_new_n316__ & ~new_new_n369__;
  assign new_new_n371__ = new_new_n368__ & ~new_new_n370__;
  assign new_new_n372__ = ~new_new_n368__ & new_new_n370__;
  assign new_new_n373__ = ~new_new_n371__ & ~new_new_n372__;
  assign new_new_n374__ = new_new_n367__ & ~new_new_n373__;
  assign new_new_n375__ = ~new_new_n367__ & new_new_n373__;
  assign new_new_n376__ = ~new_new_n374__ & ~new_new_n375__;
  assign new_new_n377__ = ~new_new_n366__ & ~new_new_n376__;
  assign new_new_n378__ = new_new_n366__ & new_new_n376__;
  assign new_new_n379__ = ~new_new_n377__ & ~new_new_n378__;
  assign new_new_n380__ = new_new_n364__ & new_new_n379__;
  assign new_new_n381__ = ~new_new_n364__ & ~new_new_n379__;
  assign new_new_n382__ = ~new_new_n380__ & ~new_new_n381__;
  assign new_new_n383__ = ~new_new_n363__ & new_new_n382__;
  assign new_new_n384__ = new_new_n363__ & ~new_new_n382__;
  assign new_new_n385__ = ~new_new_n383__ & ~new_new_n384__;
  assign new_new_n386__ = new_new_n361__ & ~new_new_n385__;
  assign new_new_n387__ = ~new_new_n361__ & new_new_n385__;
  assign new_new_n388__ = ~new_new_n386__ & ~new_new_n387__;
  assign new_new_n389__ = ~new_new_n360__ & ~new_new_n388__;
  assign new_new_n390__ = new_new_n360__ & new_new_n388__;
  assign new_new_n391__ = ~new_new_n389__ & ~new_new_n390__;
  assign new_new_n392__ = new_new_n358__ & new_new_n391__;
  assign new_new_n393__ = ~new_new_n358__ & ~new_new_n391__;
  assign new_new_n394__ = ~new_new_n392__ & ~new_new_n393__;
  assign new_new_n395__ = ~new_new_n357__ & new_new_n394__;
  assign new_new_n396__ = new_new_n357__ & ~new_new_n394__;
  assign new_new_n397__ = ~new_new_n395__ & ~new_new_n396__;
  assign new_new_n398__ = new_new_n304__ & ~new_new_n343__;
  assign new_new_n399__ = ~new_new_n342__ & ~new_new_n398__;
  assign new_new_n400__ = new_new_n397__ & new_new_n399__;
  assign new_new_n401__ = ~new_new_n397__ & ~new_new_n399__;
  assign \O[10]  = new_new_n400__ | new_new_n401__;
  assign new_new_n403__ = ~new_new_n396__ & ~new_new_n399__;
  assign new_new_n404__ = ~new_new_n395__ & ~new_new_n403__;
  assign new_new_n405__ = \A[4]  & \B[7] ;
  assign new_new_n406__ = new_new_n361__ & ~new_new_n384__;
  assign new_new_n407__ = ~new_new_n383__ & ~new_new_n406__;
  assign new_new_n408__ = \A[5]  & \B[6] ;
  assign new_new_n409__ = new_new_n364__ & ~new_new_n378__;
  assign new_new_n410__ = ~new_new_n377__ & ~new_new_n409__;
  assign new_new_n411__ = \A[6]  & \B[5] ;
  assign new_new_n412__ = \A[7]  & \B[4] ;
  assign new_new_n413__ = new_new_n367__ & ~new_new_n372__;
  assign new_new_n414__ = ~new_new_n371__ & ~new_new_n413__;
  assign new_new_n415__ = new_new_n412__ & ~new_new_n414__;
  assign new_new_n416__ = ~new_new_n412__ & new_new_n414__;
  assign new_new_n417__ = ~new_new_n415__ & ~new_new_n416__;
  assign new_new_n418__ = new_new_n411__ & new_new_n417__;
  assign new_new_n419__ = ~new_new_n411__ & ~new_new_n417__;
  assign new_new_n420__ = ~new_new_n418__ & ~new_new_n419__;
  assign new_new_n421__ = ~new_new_n410__ & new_new_n420__;
  assign new_new_n422__ = new_new_n410__ & ~new_new_n420__;
  assign new_new_n423__ = ~new_new_n421__ & ~new_new_n422__;
  assign new_new_n424__ = new_new_n408__ & ~new_new_n423__;
  assign new_new_n425__ = ~new_new_n408__ & new_new_n423__;
  assign new_new_n426__ = ~new_new_n424__ & ~new_new_n425__;
  assign new_new_n427__ = ~new_new_n407__ & ~new_new_n426__;
  assign new_new_n428__ = new_new_n407__ & new_new_n426__;
  assign new_new_n429__ = ~new_new_n427__ & ~new_new_n428__;
  assign new_new_n430__ = new_new_n405__ & new_new_n429__;
  assign new_new_n431__ = ~new_new_n405__ & ~new_new_n429__;
  assign new_new_n432__ = ~new_new_n430__ & ~new_new_n431__;
  assign new_new_n433__ = ~new_new_n404__ & new_new_n432__;
  assign new_new_n434__ = new_new_n404__ & ~new_new_n432__;
  assign new_new_n435__ = ~new_new_n433__ & ~new_new_n434__;
  assign new_new_n436__ = new_new_n358__ & ~new_new_n390__;
  assign new_new_n437__ = ~new_new_n389__ & ~new_new_n436__;
  assign new_new_n438__ = new_new_n435__ & new_new_n437__;
  assign new_new_n439__ = ~new_new_n435__ & ~new_new_n437__;
  assign \O[11]  = new_new_n438__ | new_new_n439__;
  assign new_new_n441__ = ~new_new_n434__ & ~new_new_n437__;
  assign new_new_n442__ = ~new_new_n433__ & ~new_new_n441__;
  assign new_new_n443__ = \A[5]  & \B[7] ;
  assign new_new_n444__ = new_new_n408__ & ~new_new_n422__;
  assign new_new_n445__ = ~new_new_n421__ & ~new_new_n444__;
  assign new_new_n446__ = \A[6]  & \B[6] ;
  assign new_new_n447__ = \A[7]  & \B[5] ;
  assign new_new_n448__ = new_new_n411__ & ~new_new_n416__;
  assign new_new_n449__ = ~new_new_n415__ & ~new_new_n448__;
  assign new_new_n450__ = new_new_n447__ & ~new_new_n449__;
  assign new_new_n451__ = ~new_new_n447__ & new_new_n449__;
  assign new_new_n452__ = ~new_new_n450__ & ~new_new_n451__;
  assign new_new_n453__ = new_new_n446__ & new_new_n452__;
  assign new_new_n454__ = ~new_new_n446__ & ~new_new_n452__;
  assign new_new_n455__ = ~new_new_n453__ & ~new_new_n454__;
  assign new_new_n456__ = ~new_new_n445__ & new_new_n455__;
  assign new_new_n457__ = new_new_n445__ & ~new_new_n455__;
  assign new_new_n458__ = ~new_new_n456__ & ~new_new_n457__;
  assign new_new_n459__ = new_new_n443__ & ~new_new_n458__;
  assign new_new_n460__ = ~new_new_n443__ & new_new_n458__;
  assign new_new_n461__ = ~new_new_n459__ & ~new_new_n460__;
  assign new_new_n462__ = ~new_new_n442__ & ~new_new_n461__;
  assign new_new_n463__ = new_new_n442__ & new_new_n461__;
  assign new_new_n464__ = ~new_new_n462__ & ~new_new_n463__;
  assign new_new_n465__ = new_new_n405__ & ~new_new_n428__;
  assign new_new_n466__ = ~new_new_n427__ & ~new_new_n465__;
  assign new_new_n467__ = new_new_n464__ & ~new_new_n466__;
  assign new_new_n468__ = ~new_new_n464__ & new_new_n466__;
  assign \O[12]  = ~new_new_n467__ & ~new_new_n468__;
  assign new_new_n470__ = ~new_new_n463__ & ~new_new_n466__;
  assign new_new_n471__ = ~new_new_n462__ & ~new_new_n470__;
  assign new_new_n472__ = \A[6]  & \B[7] ;
  assign new_new_n473__ = \A[7]  & \B[6] ;
  assign new_new_n474__ = new_new_n446__ & ~new_new_n451__;
  assign new_new_n475__ = ~new_new_n450__ & ~new_new_n474__;
  assign new_new_n476__ = new_new_n473__ & ~new_new_n475__;
  assign new_new_n477__ = ~new_new_n473__ & new_new_n475__;
  assign new_new_n478__ = ~new_new_n476__ & ~new_new_n477__;
  assign new_new_n479__ = new_new_n472__ & new_new_n478__;
  assign new_new_n480__ = ~new_new_n472__ & ~new_new_n478__;
  assign new_new_n481__ = ~new_new_n479__ & ~new_new_n480__;
  assign new_new_n482__ = ~new_new_n471__ & new_new_n481__;
  assign new_new_n483__ = new_new_n471__ & ~new_new_n481__;
  assign new_new_n484__ = ~new_new_n482__ & ~new_new_n483__;
  assign new_new_n485__ = new_new_n443__ & ~new_new_n457__;
  assign new_new_n486__ = ~new_new_n456__ & ~new_new_n485__;
  assign new_new_n487__ = new_new_n484__ & new_new_n486__;
  assign new_new_n488__ = ~new_new_n484__ & ~new_new_n486__;
  assign \O[13]  = new_new_n487__ | new_new_n488__;
  assign new_new_n490__ = \A[7]  & \B[7] ;
  assign new_new_n491__ = new_new_n472__ & ~new_new_n477__;
  assign new_new_n492__ = ~new_new_n476__ & ~new_new_n491__;
  assign new_new_n493__ = ~new_new_n490__ & new_new_n492__;
  assign new_new_n494__ = new_new_n490__ & ~new_new_n492__;
  assign new_new_n495__ = ~new_new_n493__ & ~new_new_n494__;
  assign new_new_n496__ = ~new_new_n483__ & ~new_new_n486__;
  assign new_new_n497__ = ~new_new_n482__ & ~new_new_n496__;
  assign new_new_n498__ = new_new_n495__ & new_new_n497__;
  assign new_new_n499__ = ~new_new_n495__ & ~new_new_n497__;
  assign \O[14]  = new_new_n498__ | new_new_n499__;
  assign new_new_n501__ = ~new_new_n493__ & ~new_new_n497__;
  assign \O[15]  = new_new_n494__ | new_new_n501__;
endmodule


