module max_57_1(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 , po0 , po1 , po2 , po3 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ;
  output po0 , po1 , po2 , po3 ;
  wire new_n10, new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31;
  assign new_n10 = pi1 & ~pi4 ;
  assign new_n11 = pi0 & ~pi3 ;
  assign new_n12 = ~pi6 & ~new_n11 ;
  assign new_n13 = ~pi1 & pi4 ;
  assign new_n14 = ~pi0 & pi3 ;
  assign new_n15 = ~new_n13 & ~new_n14 ;
  assign new_n16 = ~new_n12 & new_n15 ;
  assign new_n17 = ~new_n10 & ~new_n16 ;
  assign new_n18 = ~pi2 & pi5 ;
  assign new_n19 = ~new_n17 & ~new_n18 ;
  assign new_n20 = pi2 & ~pi5 ;
  assign new_n21 = ~pi7 & ~new_n20 ;
  assign new_n22 = ~new_n19 & new_n21 ;
  assign new_n23 = pi2 & pi8 ;
  assign new_n24 = pi5 & ~pi8 ;
  assign new_n25 = ~new_n23 & ~new_n24 ;
  assign new_n26 = pi0 & pi8 ;
  assign new_n27 = pi3 & ~pi8 ;
  assign new_n28 = ~new_n26 & ~new_n27 ;
  assign new_n29 = pi1 & pi8 ;
  assign new_n30 = pi4 & ~pi8 ;
  assign new_n31 = ~new_n29 & ~new_n30 ;
  assign po0 = new_n22 ;
  assign po1 = new_n25 ;
  assign po2 = new_n28 ;
  assign po3 = new_n31 ;
endmodule
