// Benchmark "c5315" written by ABC on Thu Jul 14 21:14:28 2022

module c5315 ( 
    G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37,
    G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79,
    G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106,
    G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140,
    G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173,
    G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209,
    G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251,
    G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293,
    G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338,
    G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389,
    G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523,
    G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691,
    G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717,
    G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115,
    // G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612,
    G594, G599, G600, G601, G602, G611, G612,
    // G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921,
    G810, G848, G849, G850, G851, G634, G815, G845, G847,
    // G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636,
    G656, G809, G593, G636,
    // G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626,
    G704, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    // G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623,
    G1002, G1004, G591, G618, G822, G838, G861, G623,
    G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000,
    G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802,
    G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826,
    G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742,
    G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843,
    G882, G767, G807, G658, G690  );
  input  G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34,
    G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76,
    G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103,
    G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121,
    G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137,
    G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170,
    G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206,
    G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248,
    G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292,
    G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335,
    G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386,
    G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514,
    G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690,
    G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552,
    G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115;
  // output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
  output G594, G599, G600, G601, G602, G611,
    // G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923,
    G612, G810, G848, G849, G850, G851, G634, G815, G845, G847,
    // G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593,
    G656, G809, G593,
    // G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    G636, G704, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    // G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861,
    G1002, G1004, G591, G618, G822, G838, G861,
    G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998,
    G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792,
    G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813,
    G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732,
    G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685,
    G688, G843, G882, G767, G807, G658, G690;
  wire new_new_n310__, new_new_n311__, new_new_n312__, new_new_n314__,
    new_new_n315__, new_new_n316__, new_new_n319__, new_new_n320__,
    new_new_n321__, new_new_n322__, new_new_n324__, new_new_n325__,
    new_new_n326__, new_new_n327__, new_new_n329__, new_new_n330__,
    new_new_n331__, new_new_n332__, new_new_n334__, new_new_n335__,
    new_new_n336__, new_new_n337__, new_new_n339__, new_new_n340__,
    new_new_n341__, new_new_n342__, new_new_n343__, new_new_n344__,
    new_new_n345__, new_new_n346__, new_new_n347__, new_new_n348__,
    new_new_n349__, new_new_n350__, new_new_n351__, new_new_n352__,
    new_new_n353__, new_new_n354__, new_new_n355__, new_new_n356__,
    new_new_n357__, new_new_n358__, new_new_n359__, new_new_n360__,
    new_new_n361__, new_new_n362__, new_new_n363__, new_new_n364__,
    new_new_n365__, new_new_n366__, new_new_n367__, new_new_n368__,
    new_new_n369__, new_new_n370__, new_new_n371__, new_new_n372__,
    new_new_n373__, new_new_n374__, new_new_n375__, new_new_n376__,
    new_new_n377__, new_new_n378__, new_new_n379__, new_new_n380__,
    new_new_n381__, new_new_n382__, new_new_n383__, new_new_n384__,
    new_new_n385__, new_new_n386__, new_new_n387__, new_new_n388__,
    new_new_n389__, new_new_n390__, new_new_n391__, new_new_n392__,
    new_new_n393__, new_new_n394__, new_new_n395__, new_new_n396__,
    new_new_n397__, new_new_n398__, new_new_n399__, new_new_n400__,
    new_new_n401__, new_new_n402__, new_new_n404__, new_new_n405__,
    new_new_n406__, new_new_n407__, new_new_n408__, new_new_n409__,
    new_new_n410__, new_new_n411__, new_new_n412__, new_new_n413__,
    new_new_n414__, new_new_n415__, new_new_n416__, new_new_n417__,
    new_new_n418__, new_new_n419__, new_new_n420__, new_new_n421__,
    new_new_n422__, new_new_n423__, new_new_n424__, new_new_n425__,
    new_new_n426__, new_new_n427__, new_new_n428__, new_new_n429__,
    new_new_n430__, new_new_n431__, new_new_n432__, new_new_n433__,
    new_new_n434__, new_new_n435__, new_new_n436__, new_new_n437__,
    new_new_n438__, new_new_n439__, new_new_n440__, new_new_n441__,
    new_new_n442__, new_new_n443__, new_new_n444__, new_new_n445__,
    new_new_n446__, new_new_n447__, new_new_n448__, new_new_n449__,
    new_new_n450__, new_new_n451__, new_new_n452__, new_new_n453__,
    new_new_n454__, new_new_n455__, new_new_n456__, new_new_n457__,
    new_new_n458__, new_new_n459__, new_new_n460__, new_new_n461__,
    new_new_n462__, new_new_n463__, new_new_n464__, new_new_n465__,
    new_new_n466__, new_new_n467__, new_new_n468__, new_new_n469__,
    new_new_n470__, new_new_n471__, new_new_n472__, new_new_n473__,
    new_new_n474__, new_new_n475__, new_new_n476__, new_new_n477__,
    new_new_n478__, new_new_n479__, new_new_n480__, new_new_n481__,
    new_new_n482__, new_new_n483__, new_new_n484__, new_new_n485__,
    new_new_n486__, new_new_n487__, new_new_n488__, new_new_n489__,
    new_new_n490__, new_new_n491__, new_new_n492__, new_new_n493__,
    new_new_n494__, new_new_n495__, new_new_n497__, new_new_n498__,
    new_new_n499__, new_new_n500__, new_new_n501__, new_new_n502__,
    new_new_n503__, new_new_n504__, new_new_n505__, new_new_n506__,
    new_new_n507__, new_new_n508__, new_new_n509__, new_new_n510__,
    new_new_n511__, new_new_n512__, new_new_n513__, new_new_n514__,
    new_new_n515__, new_new_n516__, new_new_n517__, new_new_n518__,
    new_new_n519__, new_new_n520__, new_new_n521__, new_new_n522__,
    new_new_n523__, new_new_n524__, new_new_n525__, new_new_n526__,
    new_new_n527__, new_new_n528__, new_new_n529__, new_new_n530__,
    new_new_n531__, new_new_n532__, new_new_n533__, new_new_n534__,
    new_new_n535__, new_new_n536__, new_new_n537__, new_new_n538__,
    new_new_n539__, new_new_n540__, new_new_n541__, new_new_n542__,
    new_new_n543__, new_new_n544__, new_new_n545__, new_new_n546__,
    new_new_n547__, new_new_n548__, new_new_n549__, new_new_n550__,
    new_new_n551__, new_new_n552__, new_new_n553__, new_new_n554__,
    new_new_n555__, new_new_n556__, new_new_n557__, new_new_n559__,
    new_new_n560__, new_new_n561__, new_new_n562__, new_new_n563__,
    new_new_n564__, new_new_n565__, new_new_n566__, new_new_n567__,
    new_new_n568__, new_new_n569__, new_new_n570__, new_new_n571__,
    new_new_n572__, new_new_n573__, new_new_n574__, new_new_n575__,
    new_new_n576__, new_new_n577__, new_new_n578__, new_new_n579__,
    new_new_n580__, new_new_n581__, new_new_n582__, new_new_n583__,
    new_new_n584__, new_new_n585__, new_new_n586__, new_new_n587__,
    new_new_n588__, new_new_n589__, new_new_n590__, new_new_n591__,
    new_new_n592__, new_new_n593__, new_new_n594__, new_new_n595__,
    new_new_n596__, new_new_n597__, new_new_n598__, new_new_n599__,
    new_new_n600__, new_new_n601__, new_new_n602__, new_new_n603__,
    new_new_n604__, new_new_n605__, new_new_n606__, new_new_n607__,
    new_new_n608__, new_new_n610__, new_new_n611__, new_new_n612__,
    new_new_n613__, new_new_n614__, new_new_n615__, new_new_n616__,
    new_new_n617__, new_new_n618__, new_new_n619__, new_new_n620__,
    new_new_n621__, new_new_n622__, new_new_n623__, new_new_n624__,
    new_new_n625__, new_new_n626__, new_new_n627__, new_new_n628__,
    new_new_n629__, new_new_n630__, new_new_n631__, new_new_n632__,
    new_new_n634__, new_new_n635__, new_new_n636__, new_new_n637__,
    new_new_n638__, new_new_n639__, new_new_n640__, new_new_n641__,
    new_new_n642__, new_new_n643__, new_new_n644__, new_new_n645__,
    new_new_n646__, new_new_n647__, new_new_n648__, new_new_n649__,
    new_new_n650__, new_new_n651__, new_new_n652__, new_new_n653__,
    new_new_n654__, new_new_n655__, new_new_n656__, new_new_n657__,
    new_new_n658__, new_new_n659__, new_new_n661__, new_new_n662__,
    new_new_n663__, new_new_n664__, new_new_n665__, new_new_n666__,
    new_new_n667__, new_new_n668__, new_new_n669__, new_new_n670__,
    new_new_n671__, new_new_n672__, new_new_n673__, new_new_n674__,
    new_new_n675__, new_new_n677__, new_new_n678__, new_new_n679__,
    new_new_n680__, new_new_n681__, new_new_n682__, new_new_n683__,
    new_new_n684__, new_new_n685__, new_new_n686__, new_new_n687__,
    new_new_n688__, new_new_n690__, new_new_n691__, new_new_n692__,
    new_new_n693__, new_new_n694__, new_new_n695__, new_new_n696__,
    new_new_n697__, new_new_n698__, new_new_n699__, new_new_n701__,
    new_new_n702__, new_new_n703__, new_new_n704__, new_new_n705__,
    new_new_n706__, new_new_n707__, new_new_n709__, new_new_n710__,
    new_new_n711__, new_new_n712__, new_new_n713__, new_new_n714__,
    new_new_n715__, new_new_n717__, new_new_n718__, new_new_n719__,
    new_new_n720__, new_new_n721__, new_new_n722__, new_new_n723__,
    new_new_n724__, new_new_n726__, new_new_n727__, new_new_n728__,
    new_new_n729__, new_new_n730__, new_new_n731__, new_new_n732__,
    new_new_n733__, new_new_n734__, new_new_n736__, new_new_n737__,
    new_new_n738__, new_new_n739__, new_new_n740__, new_new_n741__,
    new_new_n742__, new_new_n743__, new_new_n744__, new_new_n745__,
    new_new_n747__, new_new_n748__, new_new_n749__, new_new_n750__,
    new_new_n751__, new_new_n752__, new_new_n753__, new_new_n754__,
    new_new_n755__, new_new_n756__, new_new_n757__, new_new_n759__,
    new_new_n760__, new_new_n761__, new_new_n762__, new_new_n763__,
    new_new_n764__, new_new_n765__, new_new_n766__, new_new_n767__,
    new_new_n769__, new_new_n770__, new_new_n771__, new_new_n772__,
    new_new_n773__, new_new_n774__, new_new_n775__, new_new_n776__,
    new_new_n777__, new_new_n779__, new_new_n780__, new_new_n781__,
    new_new_n782__, new_new_n783__, new_new_n784__, new_new_n785__,
    new_new_n786__, new_new_n787__, new_new_n788__, new_new_n789__,
    new_new_n790__, new_new_n791__, new_new_n793__, new_new_n794__,
    new_new_n795__, new_new_n796__, new_new_n797__, new_new_n798__,
    new_new_n799__, new_new_n801__, new_new_n802__, new_new_n803__,
    new_new_n804__, new_new_n805__, new_new_n806__, new_new_n807__,
    new_new_n808__, new_new_n809__, new_new_n810__, new_new_n812__,
    new_new_n813__, new_new_n814__, new_new_n815__, new_new_n816__,
    new_new_n817__, new_new_n818__, new_new_n820__, new_new_n821__,
    new_new_n822__, new_new_n823__, new_new_n824__, new_new_n825__,
    new_new_n826__, new_new_n827__, new_new_n828__, new_new_n829__,
    new_new_n830__, new_new_n831__, new_new_n832__, new_new_n833__,
    new_new_n834__, new_new_n835__, new_new_n836__, new_new_n837__,
    new_new_n838__, new_new_n839__, new_new_n840__, new_new_n841__,
    new_new_n842__, new_new_n843__, new_new_n844__, new_new_n845__,
    new_new_n847__, new_new_n848__, new_new_n849__, new_new_n850__,
    new_new_n851__, new_new_n852__, new_new_n853__, new_new_n854__,
    new_new_n855__, new_new_n856__, new_new_n857__, new_new_n858__,
    new_new_n859__, new_new_n860__, new_new_n861__, new_new_n862__,
    new_new_n863__, new_new_n864__, new_new_n865__, new_new_n866__,
    new_new_n867__, new_new_n868__, new_new_n869__, new_new_n870__,
    new_new_n871__, new_new_n872__, new_new_n873__, new_new_n874__,
    new_new_n875__, new_new_n877__, new_new_n878__, new_new_n879__,
    new_new_n880__, new_new_n881__, new_new_n882__, new_new_n883__,
    new_new_n884__, new_new_n885__, new_new_n886__, new_new_n887__,
    new_new_n888__, new_new_n889__, new_new_n890__, new_new_n891__,
    new_new_n892__, new_new_n893__, new_new_n894__, new_new_n895__,
    new_new_n896__, new_new_n897__, new_new_n898__, new_new_n899__,
    new_new_n900__, new_new_n901__, new_new_n902__, new_new_n903__,
    new_new_n904__, new_new_n905__, new_new_n907__, new_new_n908__,
    new_new_n909__, new_new_n910__, new_new_n911__, new_new_n912__,
    new_new_n913__, new_new_n914__, new_new_n915__, new_new_n916__,
    new_new_n917__, new_new_n918__, new_new_n919__, new_new_n920__,
    new_new_n921__, new_new_n922__, new_new_n923__, new_new_n924__,
    new_new_n926__, new_new_n927__, new_new_n928__, new_new_n929__,
    new_new_n930__, new_new_n931__, new_new_n932__, new_new_n933__,
    new_new_n934__, new_new_n935__, new_new_n937__, new_new_n938__,
    new_new_n939__, new_new_n940__, new_new_n941__, new_new_n942__,
    new_new_n943__, new_new_n944__, new_new_n945__, new_new_n946__,
    new_new_n948__, new_new_n949__, new_new_n950__, new_new_n951__,
    new_new_n952__, new_new_n953__, new_new_n954__, new_new_n956__,
    new_new_n957__, new_new_n958__, new_new_n959__, new_new_n960__,
    new_new_n961__, new_new_n962__, new_new_n964__, new_new_n965__,
    new_new_n966__, new_new_n967__, new_new_n968__, new_new_n969__,
    new_new_n970__, new_new_n972__, new_new_n973__, new_new_n974__,
    new_new_n975__, new_new_n976__, new_new_n977__, new_new_n978__,
    new_new_n980__, new_new_n981__, new_new_n982__, new_new_n983__,
    new_new_n984__, new_new_n985__, new_new_n986__, new_new_n988__,
    new_new_n989__, new_new_n990__, new_new_n991__, new_new_n992__,
    new_new_n993__, new_new_n994__, new_new_n996__, new_new_n997__,
    new_new_n998__, new_new_n999__, new_new_n1000__, new_new_n1001__,
    new_new_n1002__, new_new_n1004__, new_new_n1005__, new_new_n1006__,
    new_new_n1007__, new_new_n1008__, new_new_n1009__, new_new_n1010__,
    new_new_n1012__, new_new_n1013__, new_new_n1014__, new_new_n1015__,
    new_new_n1016__, new_new_n1017__, new_new_n1018__, new_new_n1019__,
    new_new_n1021__, new_new_n1022__, new_new_n1023__, new_new_n1024__,
    new_new_n1025__, new_new_n1026__, new_new_n1027__, new_new_n1028__,
    new_new_n1030__, new_new_n1031__, new_new_n1032__, new_new_n1033__,
    new_new_n1034__, new_new_n1035__, new_new_n1036__, new_new_n1037__,
    new_new_n1039__, new_new_n1040__, new_new_n1041__, new_new_n1042__,
    new_new_n1043__, new_new_n1044__, new_new_n1045__, new_new_n1046__,
    new_new_n1048__, new_new_n1049__, new_new_n1050__, new_new_n1051__,
    new_new_n1052__, new_new_n1053__, new_new_n1054__, new_new_n1055__,
    new_new_n1057__, new_new_n1058__, new_new_n1059__, new_new_n1060__,
    new_new_n1061__, new_new_n1062__, new_new_n1063__, new_new_n1064__,
    new_new_n1066__, new_new_n1067__, new_new_n1068__, new_new_n1069__,
    new_new_n1070__, new_new_n1071__, new_new_n1072__, new_new_n1073__,
    new_new_n1075__, new_new_n1076__, new_new_n1077__, new_new_n1078__,
    new_new_n1079__, new_new_n1080__, new_new_n1081__, new_new_n1082__,
    new_new_n1084__, new_new_n1085__, new_new_n1086__, new_new_n1087__,
    new_new_n1088__, new_new_n1089__, new_new_n1090__, new_new_n1091__,
    new_new_n1092__, new_new_n1093__, new_new_n1094__, new_new_n1095__,
    new_new_n1096__, new_new_n1098__, new_new_n1099__, new_new_n1101__,
    new_new_n1102__, new_new_n1103__, new_new_n1104__, new_new_n1106__,
    new_new_n1107__, new_new_n1108__, new_new_n1109__, new_new_n1111__,
    new_new_n1112__, new_new_n1113__, new_new_n1114__, new_new_n1116__,
    new_new_n1117__, new_new_n1118__, new_new_n1119__, new_new_n1121__,
    new_new_n1122__, new_new_n1123__, new_new_n1124__, new_new_n1125__,
    new_new_n1126__, new_new_n1128__, new_new_n1129__, new_new_n1130__,
    new_new_n1131__, new_new_n1133__, new_new_n1134__, new_new_n1135__,
    new_new_n1136__, new_new_n1138__, new_new_n1139__, new_new_n1140__,
    new_new_n1141__, new_new_n1143__, new_new_n1144__, new_new_n1145__,
    new_new_n1146__, new_new_n1148__, new_new_n1149__, new_new_n1150__,
    new_new_n1151__, new_new_n1152__, new_new_n1153__, new_new_n1154__,
    new_new_n1156__, new_new_n1157__, new_new_n1158__, new_new_n1159__,
    new_new_n1160__, new_new_n1161__, new_new_n1162__, new_new_n1164__,
    new_new_n1165__, new_new_n1166__, new_new_n1167__, new_new_n1168__,
    new_new_n1169__, new_new_n1170__, new_new_n1172__, new_new_n1173__,
    new_new_n1174__, new_new_n1175__, new_new_n1176__, new_new_n1177__,
    new_new_n1178__, new_new_n1180__, new_new_n1181__, new_new_n1182__,
    new_new_n1183__, new_new_n1184__, new_new_n1185__, new_new_n1186__,
    new_new_n1188__, new_new_n1189__, new_new_n1190__, new_new_n1191__,
    new_new_n1192__, new_new_n1193__, new_new_n1194__, new_new_n1196__,
    new_new_n1197__, new_new_n1198__, new_new_n1199__, new_new_n1200__,
    new_new_n1201__, new_new_n1202__, new_new_n1204__, new_new_n1205__,
    new_new_n1206__, new_new_n1207__, new_new_n1208__, new_new_n1209__,
    new_new_n1210__, new_new_n1212__, new_new_n1213__, new_new_n1214__,
    new_new_n1215__, new_new_n1216__, new_new_n1217__, new_new_n1218__,
    new_new_n1219__, new_new_n1221__, new_new_n1222__, new_new_n1223__,
    new_new_n1224__, new_new_n1225__, new_new_n1226__, new_new_n1227__,
    new_new_n1228__, new_new_n1230__, new_new_n1231__, new_new_n1232__,
    new_new_n1233__, new_new_n1234__, new_new_n1235__, new_new_n1236__,
    new_new_n1237__, new_new_n1239__, new_new_n1240__, new_new_n1241__,
    new_new_n1242__, new_new_n1243__, new_new_n1244__, new_new_n1245__,
    new_new_n1246__, new_new_n1248__, new_new_n1249__, new_new_n1250__,
    new_new_n1251__, new_new_n1252__, new_new_n1253__, new_new_n1254__,
    new_new_n1255__, new_new_n1257__, new_new_n1258__, new_new_n1259__,
    new_new_n1260__, new_new_n1261__, new_new_n1262__, new_new_n1263__,
    new_new_n1264__, new_new_n1266__, new_new_n1267__, new_new_n1268__,
    new_new_n1269__, new_new_n1270__, new_new_n1271__, new_new_n1272__,
    new_new_n1273__, new_new_n1275__, new_new_n1276__, new_new_n1277__,
    new_new_n1278__, new_new_n1279__, new_new_n1280__, new_new_n1281__,
    new_new_n1282__, new_new_n1284__, new_new_n1285__, new_new_n1286__,
    new_new_n1287__, new_new_n1288__, new_new_n1289__, new_new_n1290__,
    new_new_n1291__, new_new_n1292__, new_new_n1293__, new_new_n1294__,
    new_new_n1295__, new_new_n1296__, new_new_n1297__, new_new_n1298__,
    new_new_n1299__, new_new_n1300__, new_new_n1301__, new_new_n1302__,
    new_new_n1303__, new_new_n1304__, new_new_n1305__, new_new_n1306__,
    new_new_n1307__, new_new_n1308__, new_new_n1309__, new_new_n1310__,
    new_new_n1311__, new_new_n1312__, new_new_n1313__, new_new_n1314__,
    new_new_n1315__, new_new_n1316__, new_new_n1317__, new_new_n1318__,
    new_new_n1319__, new_new_n1320__, new_new_n1321__, new_new_n1322__,
    new_new_n1323__, new_new_n1324__, new_new_n1325__, new_new_n1326__,
    new_new_n1327__, new_new_n1328__, new_new_n1329__, new_new_n1330__,
    new_new_n1331__, new_new_n1332__, new_new_n1333__, new_new_n1334__,
    new_new_n1335__, new_new_n1336__, new_new_n1337__, new_new_n1338__,
    new_new_n1339__, new_new_n1340__, new_new_n1341__, new_new_n1342__,
    new_new_n1343__, new_new_n1344__, new_new_n1345__, new_new_n1346__,
    new_new_n1347__, new_new_n1348__, new_new_n1349__, new_new_n1350__,
    new_new_n1351__, new_new_n1352__, new_new_n1353__, new_new_n1354__,
    new_new_n1355__, new_new_n1356__, new_new_n1357__, new_new_n1358__,
    new_new_n1359__, new_new_n1360__, new_new_n1361__, new_new_n1362__,
    new_new_n1363__, new_new_n1364__, new_new_n1365__, new_new_n1366__,
    new_new_n1367__, new_new_n1368__, new_new_n1369__, new_new_n1370__,
    new_new_n1371__, new_new_n1372__, new_new_n1373__, new_new_n1374__,
    new_new_n1375__, new_new_n1376__, new_new_n1377__, new_new_n1378__,
    new_new_n1379__, new_new_n1380__, new_new_n1381__, new_new_n1382__,
    new_new_n1383__, new_new_n1384__, new_new_n1385__, new_new_n1386__,
    new_new_n1387__, new_new_n1388__, new_new_n1389__, new_new_n1390__,
    new_new_n1391__, new_new_n1392__, new_new_n1393__, new_new_n1395__,
    new_new_n1396__, new_new_n1397__, new_new_n1398__, new_new_n1399__,
    new_new_n1400__, new_new_n1401__, new_new_n1402__, new_new_n1403__,
    new_new_n1404__, new_new_n1405__, new_new_n1406__, new_new_n1407__,
    new_new_n1408__, new_new_n1409__, new_new_n1410__, new_new_n1411__,
    new_new_n1412__, new_new_n1413__, new_new_n1414__, new_new_n1415__,
    new_new_n1416__, new_new_n1417__, new_new_n1418__, new_new_n1419__,
    new_new_n1420__, new_new_n1421__, new_new_n1422__, new_new_n1423__,
    new_new_n1424__, new_new_n1425__, new_new_n1426__, new_new_n1427__,
    new_new_n1428__, new_new_n1429__, new_new_n1430__, new_new_n1431__,
    new_new_n1432__, new_new_n1433__, new_new_n1434__, new_new_n1435__,
    new_new_n1436__, new_new_n1437__, new_new_n1438__, new_new_n1439__,
    new_new_n1440__, new_new_n1441__, new_new_n1442__, new_new_n1443__,
    new_new_n1444__, new_new_n1445__, new_new_n1446__, new_new_n1447__,
    new_new_n1448__, new_new_n1449__, new_new_n1450__, new_new_n1451__,
    new_new_n1452__, new_new_n1453__, new_new_n1454__, new_new_n1455__,
    new_new_n1456__, new_new_n1457__, new_new_n1458__, new_new_n1459__,
    new_new_n1460__, new_new_n1461__, new_new_n1462__, new_new_n1463__,
    new_new_n1464__, new_new_n1465__, new_new_n1466__, new_new_n1467__,
    new_new_n1468__, new_new_n1469__, new_new_n1470__, new_new_n1471__,
    new_new_n1472__, new_new_n1473__, new_new_n1474__, new_new_n1475__,
    new_new_n1476__, new_new_n1477__, new_new_n1478__, new_new_n1479__,
    new_new_n1480__, new_new_n1481__, new_new_n1482__, new_new_n1483__,
    new_new_n1484__, new_new_n1485__, new_new_n1486__, new_new_n1487__,
    new_new_n1488__, new_new_n1489__, new_new_n1490__, new_new_n1491__,
    new_new_n1492__, new_new_n1493__, new_new_n1494__, new_new_n1495__,
    new_new_n1496__, new_new_n1497__, new_new_n1498__, new_new_n1499__,
    new_new_n1500__, new_new_n1501__, new_new_n1502__, new_new_n1503__,
    new_new_n1504__, new_new_n1505__, new_new_n1506__, new_new_n1507__,
    new_new_n1508__, new_new_n1509__, new_new_n1510__, new_new_n1511__,
    new_new_n1512__, new_new_n1513__, new_new_n1514__, new_new_n1515__,
    new_new_n1516__, new_new_n1517__, new_new_n1518__, new_new_n1519__,
    new_new_n1520__, new_new_n1521__, new_new_n1522__, new_new_n1523__,
    new_new_n1524__, new_new_n1525__, new_new_n1526__, new_new_n1527__,
    new_new_n1528__, new_new_n1529__, new_new_n1530__, new_new_n1531__,
    new_new_n1532__, new_new_n1533__, new_new_n1534__, new_new_n1535__,
    new_new_n1536__, new_new_n1537__, new_new_n1538__, new_new_n1539__,
    new_new_n1540__, new_new_n1541__, new_new_n1542__, new_new_n1543__,
    new_new_n1544__, new_new_n1545__, new_new_n1546__, new_new_n1547__,
    new_new_n1548__, new_new_n1549__, new_new_n1550__, new_new_n1551__,
    new_new_n1552__, new_new_n1553__, new_new_n1554__, new_new_n1555__,
    new_new_n1556__, new_new_n1557__, new_new_n1558__, new_new_n1559__,
    new_new_n1560__, new_new_n1561__, new_new_n1562__, new_new_n1563__,
    new_new_n1564__, new_new_n1565__, new_new_n1566__, new_new_n1567__,
    new_new_n1568__, new_new_n1570__, new_new_n1571__, new_new_n1572__,
    new_new_n1573__, new_new_n1574__, new_new_n1575__, new_new_n1576__,
    new_new_n1577__, new_new_n1578__, new_new_n1579__, new_new_n1580__,
    new_new_n1582__, new_new_n1583__, new_new_n1584__, new_new_n1585__,
    new_new_n1586__, new_new_n1587__, new_new_n1588__, new_new_n1590__,
    new_new_n1591__, new_new_n1592__, new_new_n1593__, new_new_n1594__,
    new_new_n1595__, new_new_n1596__, new_new_n1597__, new_new_n1599__,
    new_new_n1600__, new_new_n1601__, new_new_n1602__, new_new_n1603__,
    new_new_n1604__, new_new_n1605__, new_new_n1606__;
  assign G601 = G552 & G562;
  assign G810 = G141 & G145;
  assign G634 = G1 & G373;
  assign G815 = G136 & ~G3173;
  assign G845 = ~G27 | G2824;
  assign G847 = ~G386 | ~G556;
  assign G809 = ~G27 | ~G31;
  assign G656 = ~G140 | G809;
  assign new_new_n310__ = ~G86 & ~G2358;
  assign new_new_n311__ = ~G87 & G2358;
  assign new_new_n312__ = ~G809 & ~new_new_n310__;
  assign G636 = new_new_n311__ | ~new_new_n312__;
  assign new_new_n314__ = ~G88 & ~G2358;
  assign new_new_n315__ = ~G34 & G2358;
  assign new_new_n316__ = ~G809 & ~new_new_n314__;
  assign G704 = new_new_n315__ | ~new_new_n316__;
  assign G820 = ~G83 | G809;
  assign new_new_n319__ = G24 & ~G2358;
  assign new_new_n320__ = G25 & G2358;
  assign new_new_n321__ = ~G809 & ~new_new_n319__;
  assign new_new_n322__ = ~new_new_n320__ & new_new_n321__;
  assign G639 = G141 & ~new_new_n322__;
  assign new_new_n324__ = G26 & ~G2358;
  assign new_new_n325__ = G81 & G2358;
  assign new_new_n326__ = ~G809 & ~new_new_n324__;
  assign new_new_n327__ = ~new_new_n325__ & new_new_n326__;
  assign G673 = G141 & ~new_new_n327__;
  assign new_new_n329__ = G79 & ~G2358;
  assign new_new_n330__ = G23 & G2358;
  assign new_new_n331__ = ~G809 & ~new_new_n329__;
  assign new_new_n332__ = ~new_new_n330__ & new_new_n331__;
  assign G707 = G141 & ~new_new_n332__;
  assign new_new_n334__ = G82 & ~G2358;
  assign new_new_n335__ = G80 & G2358;
  assign new_new_n336__ = ~G809 & ~new_new_n334__;
  assign new_new_n337__ = ~new_new_n335__ & new_new_n336__;
  assign G715 = G141 & ~new_new_n337__;
  assign new_new_n339__ = ~G324 & ~G3550;
  assign new_new_n340__ = G324 & ~G3552;
  assign new_new_n341__ = G503 & ~new_new_n339__;
  assign new_new_n342__ = ~new_new_n340__ & new_new_n341__;
  assign new_new_n343__ = ~G324 & G3548;
  assign new_new_n344__ = G324 & G3546;
  assign new_new_n345__ = ~G503 & ~new_new_n343__;
  assign new_new_n346__ = ~new_new_n344__ & new_new_n345__;
  assign new_new_n347__ = ~new_new_n342__ & ~new_new_n346__;
  assign new_new_n348__ = ~G251 & ~G302;
  assign new_new_n349__ = ~G248 & G302;
  assign new_new_n350__ = ~new_new_n348__ & ~new_new_n349__;
  assign new_new_n351__ = ~G254 & ~G293;
  assign new_new_n352__ = ~G242 & G293;
  assign new_new_n353__ = ~new_new_n351__ & ~new_new_n352__;
  assign new_new_n354__ = ~G251 & ~G361;
  assign new_new_n355__ = ~G248 & G361;
  assign new_new_n356__ = ~new_new_n354__ & ~new_new_n355__;
  assign new_new_n357__ = ~G514 & ~G3546;
  assign new_new_n358__ = G514 & G3552;
  assign new_new_n359__ = ~new_new_n357__ & ~new_new_n358__;
  assign new_new_n360__ = ~G351 & ~G3550;
  assign new_new_n361__ = G351 & ~G3552;
  assign new_new_n362__ = G534 & ~new_new_n360__;
  assign new_new_n363__ = ~new_new_n361__ & new_new_n362__;
  assign new_new_n364__ = ~G351 & G3548;
  assign new_new_n365__ = G351 & G3546;
  assign new_new_n366__ = ~G534 & ~new_new_n364__;
  assign new_new_n367__ = ~new_new_n365__ & new_new_n366__;
  assign new_new_n368__ = ~new_new_n363__ & ~new_new_n367__;
  assign new_new_n369__ = ~G341 & ~G3550;
  assign new_new_n370__ = G341 & ~G3552;
  assign new_new_n371__ = G523 & ~new_new_n369__;
  assign new_new_n372__ = ~new_new_n370__ & new_new_n371__;
  assign new_new_n373__ = ~G341 & G3548;
  assign new_new_n374__ = G341 & G3546;
  assign new_new_n375__ = ~G523 & ~new_new_n373__;
  assign new_new_n376__ = ~new_new_n374__ & new_new_n375__;
  assign new_new_n377__ = ~new_new_n372__ & ~new_new_n376__;
  assign new_new_n378__ = G251 & ~G316;
  assign new_new_n379__ = G248 & G316;
  assign new_new_n380__ = G490 & ~new_new_n378__;
  assign new_new_n381__ = ~new_new_n379__ & new_new_n380__;
  assign new_new_n382__ = ~G254 & ~G316;
  assign new_new_n383__ = ~G242 & G316;
  assign new_new_n384__ = ~G490 & ~new_new_n382__;
  assign new_new_n385__ = ~new_new_n383__ & new_new_n384__;
  assign new_new_n386__ = ~new_new_n381__ & ~new_new_n385__;
  assign new_new_n387__ = G251 & ~G308;
  assign new_new_n388__ = G248 & G308;
  assign new_new_n389__ = G479 & ~new_new_n387__;
  assign new_new_n390__ = ~new_new_n388__ & new_new_n389__;
  assign new_new_n391__ = ~G254 & ~G308;
  assign new_new_n392__ = ~G242 & G308;
  assign new_new_n393__ = ~G479 & ~new_new_n391__;
  assign new_new_n394__ = ~new_new_n392__ & new_new_n393__;
  assign new_new_n395__ = ~new_new_n390__ & ~new_new_n394__;
  assign new_new_n396__ = new_new_n386__ & new_new_n395__;
  assign new_new_n397__ = new_new_n350__ & ~new_new_n353__;
  assign new_new_n398__ = new_new_n356__ & new_new_n359__;
  assign new_new_n399__ = new_new_n397__ & new_new_n398__;
  assign new_new_n400__ = new_new_n347__ & new_new_n399__;
  assign new_new_n401__ = new_new_n368__ & new_new_n377__;
  assign new_new_n402__ = new_new_n400__ & new_new_n401__;
  assign G598 = new_new_n396__ & new_new_n402__;
  assign new_new_n404__ = ~G257 & ~G3550;
  assign new_new_n405__ = G257 & ~G3552;
  assign new_new_n406__ = G389 & ~new_new_n404__;
  assign new_new_n407__ = ~new_new_n405__ & new_new_n406__;
  assign new_new_n408__ = ~G257 & G3548;
  assign new_new_n409__ = G257 & G3546;
  assign new_new_n410__ = ~G389 & ~new_new_n408__;
  assign new_new_n411__ = ~new_new_n409__ & new_new_n410__;
  assign new_new_n412__ = ~new_new_n407__ & ~new_new_n411__;
  assign new_new_n413__ = G234 & G435;
  assign new_new_n414__ = ~G3552 & new_new_n413__;
  assign new_new_n415__ = ~G234 & G435;
  assign new_new_n416__ = ~G3550 & new_new_n415__;
  assign new_new_n417__ = ~G234 & ~G3548;
  assign new_new_n418__ = G234 & ~G3546;
  assign new_new_n419__ = ~G435 & ~new_new_n417__;
  assign new_new_n420__ = ~new_new_n418__ & new_new_n419__;
  assign new_new_n421__ = ~new_new_n414__ & ~new_new_n416__;
  assign new_new_n422__ = ~new_new_n420__ & new_new_n421__;
  assign new_new_n423__ = ~G206 & G251;
  assign new_new_n424__ = G206 & G248;
  assign new_new_n425__ = G446 & ~new_new_n423__;
  assign new_new_n426__ = ~new_new_n424__ & new_new_n425__;
  assign new_new_n427__ = ~G206 & ~G254;
  assign new_new_n428__ = G206 & ~G242;
  assign new_new_n429__ = ~G446 & ~new_new_n427__;
  assign new_new_n430__ = ~new_new_n428__ & new_new_n429__;
  assign new_new_n431__ = ~new_new_n426__ & ~new_new_n430__;
  assign new_new_n432__ = G226 & G422;
  assign new_new_n433__ = ~G3552 & new_new_n432__;
  assign new_new_n434__ = ~G226 & G422;
  assign new_new_n435__ = ~G3550 & new_new_n434__;
  assign new_new_n436__ = ~G226 & ~G3548;
  assign new_new_n437__ = G226 & ~G3546;
  assign new_new_n438__ = ~G422 & ~new_new_n436__;
  assign new_new_n439__ = ~new_new_n437__ & new_new_n438__;
  assign new_new_n440__ = ~new_new_n433__ & ~new_new_n435__;
  assign new_new_n441__ = ~new_new_n439__ & new_new_n440__;
  assign new_new_n442__ = ~G281 & ~G3550;
  assign new_new_n443__ = G281 & ~G3552;
  assign new_new_n444__ = G374 & ~new_new_n442__;
  assign new_new_n445__ = ~new_new_n443__ & new_new_n444__;
  assign new_new_n446__ = ~G281 & G3548;
  assign new_new_n447__ = G281 & G3546;
  assign new_new_n448__ = ~G374 & ~new_new_n446__;
  assign new_new_n449__ = ~new_new_n447__ & new_new_n448__;
  assign new_new_n450__ = ~new_new_n445__ & ~new_new_n449__;
  assign new_new_n451__ = ~G265 & ~G3550;
  assign new_new_n452__ = G265 & ~G3552;
  assign new_new_n453__ = G400 & ~new_new_n451__;
  assign new_new_n454__ = ~new_new_n452__ & new_new_n453__;
  assign new_new_n455__ = ~G265 & G3548;
  assign new_new_n456__ = G265 & G3546;
  assign new_new_n457__ = ~G400 & ~new_new_n455__;
  assign new_new_n458__ = ~new_new_n456__ & new_new_n457__;
  assign new_new_n459__ = ~new_new_n454__ & ~new_new_n458__;
  assign new_new_n460__ = G210 & G457;
  assign new_new_n461__ = ~G3552 & new_new_n460__;
  assign new_new_n462__ = ~G210 & G457;
  assign new_new_n463__ = ~G3550 & new_new_n462__;
  assign new_new_n464__ = ~G210 & ~G3548;
  assign new_new_n465__ = G210 & ~G3546;
  assign new_new_n466__ = ~G457 & ~new_new_n464__;
  assign new_new_n467__ = ~new_new_n465__ & new_new_n466__;
  assign new_new_n468__ = ~new_new_n461__ & ~new_new_n463__;
  assign new_new_n469__ = ~new_new_n467__ & new_new_n468__;
  assign new_new_n470__ = ~G273 & ~G3550;
  assign new_new_n471__ = G273 & ~G3552;
  assign new_new_n472__ = G411 & ~new_new_n470__;
  assign new_new_n473__ = ~new_new_n471__ & new_new_n472__;
  assign new_new_n474__ = ~G273 & G3548;
  assign new_new_n475__ = G273 & G3546;
  assign new_new_n476__ = ~G411 & ~new_new_n474__;
  assign new_new_n477__ = ~new_new_n475__ & new_new_n476__;
  assign new_new_n478__ = ~new_new_n473__ & ~new_new_n477__;
  assign new_new_n479__ = G218 & G468;
  assign new_new_n480__ = ~G3552 & new_new_n479__;
  assign new_new_n481__ = ~G218 & G468;
  assign new_new_n482__ = ~G3550 & new_new_n481__;
  assign new_new_n483__ = ~G218 & ~G3548;
  assign new_new_n484__ = G218 & ~G3546;
  assign new_new_n485__ = ~G468 & ~new_new_n483__;
  assign new_new_n486__ = ~new_new_n484__ & new_new_n485__;
  assign new_new_n487__ = ~new_new_n480__ & ~new_new_n482__;
  assign new_new_n488__ = ~new_new_n486__ & new_new_n487__;
  assign new_new_n489__ = new_new_n412__ & ~new_new_n422__;
  assign new_new_n490__ = new_new_n431__ & ~new_new_n441__;
  assign new_new_n491__ = new_new_n450__ & new_new_n459__;
  assign new_new_n492__ = ~new_new_n469__ & new_new_n478__;
  assign new_new_n493__ = ~new_new_n488__ & new_new_n492__;
  assign new_new_n494__ = new_new_n490__ & new_new_n491__;
  assign new_new_n495__ = new_new_n489__ & new_new_n494__;
  assign G610 = new_new_n493__ & new_new_n495__;
  assign new_new_n497__ = ~G233 & G335;
  assign new_new_n498__ = ~G226 & ~G335;
  assign new_new_n499__ = ~new_new_n497__ & ~new_new_n498__;
  assign new_new_n500__ = G422 & new_new_n499__;
  assign new_new_n501__ = ~G422 & ~new_new_n499__;
  assign new_new_n502__ = ~new_new_n500__ & ~new_new_n501__;
  assign new_new_n503__ = ~G225 & G335;
  assign new_new_n504__ = ~G218 & ~G335;
  assign new_new_n505__ = ~new_new_n503__ & ~new_new_n504__;
  assign new_new_n506__ = G468 & new_new_n505__;
  assign new_new_n507__ = ~G468 & ~new_new_n505__;
  assign new_new_n508__ = ~new_new_n506__ & ~new_new_n507__;
  assign new_new_n509__ = ~G217 & G335;
  assign new_new_n510__ = ~G210 & ~G335;
  assign new_new_n511__ = ~new_new_n509__ & ~new_new_n510__;
  assign new_new_n512__ = G457 & new_new_n511__;
  assign new_new_n513__ = ~G457 & ~new_new_n511__;
  assign new_new_n514__ = ~new_new_n512__ & ~new_new_n513__;
  assign new_new_n515__ = new_new_n502__ & new_new_n508__;
  assign new_new_n516__ = new_new_n514__ & new_new_n515__;
  assign new_new_n517__ = ~G209 & G335;
  assign new_new_n518__ = ~G206 & ~G335;
  assign new_new_n519__ = ~new_new_n517__ & ~new_new_n518__;
  assign new_new_n520__ = G446 & new_new_n519__;
  assign new_new_n521__ = ~G446 & ~new_new_n519__;
  assign new_new_n522__ = ~new_new_n520__ & ~new_new_n521__;
  assign new_new_n523__ = new_new_n516__ & new_new_n522__;
  assign new_new_n524__ = ~G241 & G335;
  assign new_new_n525__ = ~G234 & ~G335;
  assign new_new_n526__ = ~new_new_n524__ & ~new_new_n525__;
  assign new_new_n527__ = G435 & new_new_n526__;
  assign new_new_n528__ = ~G435 & ~new_new_n526__;
  assign new_new_n529__ = ~new_new_n527__ & ~new_new_n528__;
  assign new_new_n530__ = ~G288 & G335;
  assign new_new_n531__ = ~G281 & ~G335;
  assign new_new_n532__ = ~new_new_n530__ & ~new_new_n531__;
  assign new_new_n533__ = G374 & new_new_n532__;
  assign new_new_n534__ = ~G374 & ~new_new_n532__;
  assign new_new_n535__ = ~new_new_n533__ & ~new_new_n534__;
  assign new_new_n536__ = ~G280 & G335;
  assign new_new_n537__ = ~G273 & ~G335;
  assign new_new_n538__ = ~new_new_n536__ & ~new_new_n537__;
  assign new_new_n539__ = G411 & new_new_n538__;
  assign new_new_n540__ = ~G411 & ~new_new_n538__;
  assign new_new_n541__ = ~new_new_n539__ & ~new_new_n540__;
  assign new_new_n542__ = new_new_n535__ & new_new_n541__;
  assign new_new_n543__ = ~G264 & G335;
  assign new_new_n544__ = ~G257 & ~G335;
  assign new_new_n545__ = ~new_new_n543__ & ~new_new_n544__;
  assign new_new_n546__ = G389 & new_new_n545__;
  assign new_new_n547__ = ~G389 & ~new_new_n545__;
  assign new_new_n548__ = ~new_new_n546__ & ~new_new_n547__;
  assign new_new_n549__ = ~G272 & G335;
  assign new_new_n550__ = ~G265 & ~G335;
  assign new_new_n551__ = ~new_new_n549__ & ~new_new_n550__;
  assign new_new_n552__ = G400 & new_new_n551__;
  assign new_new_n553__ = ~G400 & ~new_new_n551__;
  assign new_new_n554__ = ~new_new_n552__ & ~new_new_n553__;
  assign new_new_n555__ = new_new_n548__ & new_new_n554__;
  assign new_new_n556__ = new_new_n542__ & new_new_n555__;
  assign new_new_n557__ = new_new_n529__ & new_new_n556__;
  assign G588 = new_new_n523__ & new_new_n557__;
  assign new_new_n559__ = ~G299 & G332;
  assign new_new_n560__ = ~G293 & ~G332;
  assign new_new_n561__ = ~new_new_n559__ & ~new_new_n560__;
  assign new_new_n562__ = ~G307 & G332;
  assign new_new_n563__ = ~G302 & ~G332;
  assign new_new_n564__ = ~new_new_n562__ & ~new_new_n563__;
  assign new_new_n565__ = ~new_new_n561__ & ~new_new_n564__;
  assign new_new_n566__ = ~G315 & G332;
  assign new_new_n567__ = ~G308 & ~G332;
  assign new_new_n568__ = ~new_new_n566__ & ~new_new_n567__;
  assign new_new_n569__ = G479 & new_new_n568__;
  assign new_new_n570__ = ~G479 & ~new_new_n568__;
  assign new_new_n571__ = ~new_new_n569__ & ~new_new_n570__;
  assign new_new_n572__ = ~G323 & G332;
  assign new_new_n573__ = ~G316 & ~G332;
  assign new_new_n574__ = ~new_new_n572__ & ~new_new_n573__;
  assign new_new_n575__ = G490 & new_new_n574__;
  assign new_new_n576__ = ~G490 & ~new_new_n574__;
  assign new_new_n577__ = ~new_new_n575__ & ~new_new_n576__;
  assign new_new_n578__ = new_new_n571__ & new_new_n577__;
  assign new_new_n579__ = ~G331 & G332;
  assign new_new_n580__ = ~G324 & ~G332;
  assign new_new_n581__ = ~new_new_n579__ & ~new_new_n580__;
  assign new_new_n582__ = G503 & new_new_n581__;
  assign new_new_n583__ = ~G503 & ~new_new_n581__;
  assign new_new_n584__ = ~new_new_n582__ & ~new_new_n583__;
  assign new_new_n585__ = G332 & ~G358;
  assign new_new_n586__ = ~G332 & ~G351;
  assign new_new_n587__ = ~new_new_n585__ & ~new_new_n586__;
  assign new_new_n588__ = G534 & new_new_n587__;
  assign new_new_n589__ = ~G534 & ~new_new_n587__;
  assign new_new_n590__ = ~new_new_n588__ & ~new_new_n589__;
  assign new_new_n591__ = G332 & ~G366;
  assign new_new_n592__ = ~G332 & ~G361;
  assign new_new_n593__ = ~new_new_n591__ & ~new_new_n592__;
  assign new_new_n594__ = new_new_n590__ & ~new_new_n593__;
  assign new_new_n595__ = G332 & ~G338;
  assign new_new_n596__ = G514 & ~new_new_n595__;
  assign new_new_n597__ = ~G514 & new_new_n595__;
  assign new_new_n598__ = ~new_new_n596__ & ~new_new_n597__;
  assign new_new_n599__ = G332 & ~G348;
  assign new_new_n600__ = ~G332 & ~G341;
  assign new_new_n601__ = ~new_new_n599__ & ~new_new_n600__;
  assign new_new_n602__ = G523 & new_new_n601__;
  assign new_new_n603__ = ~G523 & ~new_new_n601__;
  assign new_new_n604__ = ~new_new_n602__ & ~new_new_n603__;
  assign new_new_n605__ = new_new_n598__ & new_new_n604__;
  assign new_new_n606__ = new_new_n594__ & new_new_n605__;
  assign new_new_n607__ = new_new_n584__ & new_new_n606__;
  assign new_new_n608__ = new_new_n565__ & new_new_n578__;
  assign G615 = new_new_n607__ & new_new_n608__;
  assign new_new_n610__ = ~G308 & ~G316;
  assign new_new_n611__ = G308 & G316;
  assign new_new_n612__ = ~new_new_n610__ & ~new_new_n611__;
  assign new_new_n613__ = ~G361 & ~G369;
  assign new_new_n614__ = G361 & G369;
  assign new_new_n615__ = ~new_new_n613__ & ~new_new_n614__;
  assign new_new_n616__ = new_new_n612__ & ~new_new_n615__;
  assign new_new_n617__ = ~new_new_n612__ & new_new_n615__;
  assign new_new_n618__ = ~new_new_n616__ & ~new_new_n617__;
  assign new_new_n619__ = ~G341 & ~G351;
  assign new_new_n620__ = G341 & G351;
  assign new_new_n621__ = ~new_new_n619__ & ~new_new_n620__;
  assign new_new_n622__ = G324 & new_new_n621__;
  assign new_new_n623__ = ~G324 & ~new_new_n621__;
  assign new_new_n624__ = ~new_new_n622__ & ~new_new_n623__;
  assign new_new_n625__ = G293 & ~G302;
  assign new_new_n626__ = ~G293 & G302;
  assign new_new_n627__ = ~new_new_n625__ & ~new_new_n626__;
  assign new_new_n628__ = new_new_n624__ & ~new_new_n627__;
  assign new_new_n629__ = ~new_new_n624__ & new_new_n627__;
  assign new_new_n630__ = ~new_new_n628__ & ~new_new_n629__;
  assign new_new_n631__ = new_new_n618__ & new_new_n630__;
  assign new_new_n632__ = ~new_new_n618__ & ~new_new_n630__;
  assign G1002 = ~new_new_n631__ & ~new_new_n632__;
  assign new_new_n634__ = ~G218 & ~G226;
  assign new_new_n635__ = G218 & G226;
  assign new_new_n636__ = ~new_new_n634__ & ~new_new_n635__;
  assign new_new_n637__ = ~G234 & ~G257;
  assign new_new_n638__ = G234 & G257;
  assign new_new_n639__ = ~new_new_n637__ & ~new_new_n638__;
  assign new_new_n640__ = G281 & new_new_n639__;
  assign new_new_n641__ = ~G281 & ~new_new_n639__;
  assign new_new_n642__ = ~new_new_n640__ & ~new_new_n641__;
  assign new_new_n643__ = new_new_n636__ & ~new_new_n642__;
  assign new_new_n644__ = ~new_new_n636__ & new_new_n642__;
  assign new_new_n645__ = ~new_new_n643__ & ~new_new_n644__;
  assign new_new_n646__ = ~G265 & ~G273;
  assign new_new_n647__ = G265 & G273;
  assign new_new_n648__ = ~new_new_n646__ & ~new_new_n647__;
  assign new_new_n649__ = G289 & new_new_n648__;
  assign new_new_n650__ = ~G289 & ~new_new_n648__;
  assign new_new_n651__ = ~new_new_n649__ & ~new_new_n650__;
  assign new_new_n652__ = G206 & ~G210;
  assign new_new_n653__ = ~G206 & G210;
  assign new_new_n654__ = ~new_new_n652__ & ~new_new_n653__;
  assign new_new_n655__ = new_new_n651__ & ~new_new_n654__;
  assign new_new_n656__ = ~new_new_n651__ & new_new_n654__;
  assign new_new_n657__ = ~new_new_n655__ & ~new_new_n656__;
  assign new_new_n658__ = new_new_n645__ & new_new_n657__;
  assign new_new_n659__ = ~new_new_n645__ & ~new_new_n657__;
  assign G1004 = new_new_n658__ | new_new_n659__;
  assign new_new_n661__ = new_new_n500__ & new_new_n508__;
  assign new_new_n662__ = ~new_new_n506__ & ~new_new_n661__;
  assign new_new_n663__ = ~new_new_n512__ & new_new_n662__;
  assign new_new_n664__ = ~new_new_n513__ & ~new_new_n663__;
  assign new_new_n665__ = ~new_new_n521__ & new_new_n664__;
  assign new_new_n666__ = new_new_n533__ & new_new_n541__;
  assign new_new_n667__ = ~new_new_n539__ & ~new_new_n552__;
  assign new_new_n668__ = ~new_new_n666__ & new_new_n667__;
  assign new_new_n669__ = ~new_new_n553__ & ~new_new_n668__;
  assign new_new_n670__ = ~new_new_n546__ & ~new_new_n669__;
  assign new_new_n671__ = ~new_new_n547__ & ~new_new_n670__;
  assign new_new_n672__ = ~new_new_n527__ & ~new_new_n671__;
  assign new_new_n673__ = ~new_new_n528__ & ~new_new_n672__;
  assign new_new_n674__ = new_new_n523__ & new_new_n673__;
  assign new_new_n675__ = ~new_new_n520__ & ~new_new_n665__;
  assign G591 = new_new_n674__ | ~new_new_n675__;
  assign new_new_n677__ = ~new_new_n588__ & ~new_new_n593__;
  assign new_new_n678__ = ~new_new_n589__ & ~new_new_n603__;
  assign new_new_n679__ = ~new_new_n677__ & new_new_n678__;
  assign new_new_n680__ = ~new_new_n602__ & ~new_new_n679__;
  assign new_new_n681__ = ~new_new_n597__ & ~new_new_n680__;
  assign new_new_n682__ = ~new_new_n596__ & ~new_new_n681__;
  assign new_new_n683__ = new_new_n584__ & ~new_new_n682__;
  assign new_new_n684__ = ~new_new_n582__ & ~new_new_n683__;
  assign new_new_n685__ = new_new_n578__ & ~new_new_n684__;
  assign new_new_n686__ = ~new_new_n569__ & ~new_new_n575__;
  assign new_new_n687__ = ~new_new_n570__ & ~new_new_n686__;
  assign new_new_n688__ = new_new_n565__ & ~new_new_n687__;
  assign G618 = new_new_n685__ | ~new_new_n688__;
  assign new_new_n690__ = ~G4091 & ~G4092;
  assign new_new_n691__ = ~new_new_n356__ & new_new_n690__;
  assign new_new_n692__ = ~G54 & ~new_new_n593__;
  assign new_new_n693__ = G54 & new_new_n593__;
  assign new_new_n694__ = ~new_new_n692__ & ~new_new_n693__;
  assign new_new_n695__ = G4091 & ~G4092;
  assign new_new_n696__ = ~new_new_n694__ & new_new_n695__;
  assign new_new_n697__ = ~G4091 & G4092;
  assign new_new_n698__ = G131 & new_new_n697__;
  assign new_new_n699__ = ~new_new_n691__ & ~new_new_n698__;
  assign G822 = ~new_new_n696__ & new_new_n699__;
  assign new_new_n701__ = ~new_new_n368__ & new_new_n690__;
  assign new_new_n702__ = G129 & new_new_n697__;
  assign new_new_n703__ = new_new_n590__ & ~new_new_n692__;
  assign new_new_n704__ = ~new_new_n590__ & new_new_n692__;
  assign new_new_n705__ = new_new_n695__ & ~new_new_n703__;
  assign new_new_n706__ = ~new_new_n704__ & new_new_n705__;
  assign new_new_n707__ = ~new_new_n701__ & ~new_new_n702__;
  assign G838 = ~new_new_n706__ & new_new_n707__;
  assign new_new_n709__ = ~new_new_n450__ & new_new_n690__;
  assign new_new_n710__ = G4 & new_new_n535__;
  assign new_new_n711__ = ~G4 & ~new_new_n535__;
  assign new_new_n712__ = ~new_new_n710__ & ~new_new_n711__;
  assign new_new_n713__ = new_new_n695__ & new_new_n712__;
  assign new_new_n714__ = G117 & new_new_n697__;
  assign new_new_n715__ = ~new_new_n709__ & ~new_new_n714__;
  assign G861 = ~new_new_n713__ & new_new_n715__;
  assign new_new_n717__ = G54 & new_new_n607__;
  assign new_new_n718__ = new_new_n684__ & ~new_new_n717__;
  assign new_new_n719__ = new_new_n578__ & ~new_new_n718__;
  assign new_new_n720__ = ~new_new_n687__ & ~new_new_n719__;
  assign new_new_n721__ = ~new_new_n561__ & ~new_new_n720__;
  assign new_new_n722__ = new_new_n561__ & new_new_n564__;
  assign new_new_n723__ = ~new_new_n565__ & ~new_new_n722__;
  assign new_new_n724__ = new_new_n720__ & new_new_n723__;
  assign G623 = new_new_n721__ | new_new_n724__;
  assign new_new_n726__ = ~G4087 & ~G4088;
  assign new_new_n727__ = ~G822 & new_new_n726__;
  assign new_new_n728__ = ~G4087 & G4088;
  assign new_new_n729__ = ~G861 & new_new_n728__;
  assign new_new_n730__ = ~G11 & ~G4088;
  assign new_new_n731__ = ~G61 & G4088;
  assign new_new_n732__ = G4087 & ~new_new_n730__;
  assign new_new_n733__ = ~new_new_n731__ & new_new_n732__;
  assign new_new_n734__ = ~new_new_n727__ & ~new_new_n733__;
  assign G722 = new_new_n729__ | ~new_new_n734__;
  assign new_new_n736__ = ~new_new_n347__ & new_new_n690__;
  assign new_new_n737__ = ~new_new_n606__ & new_new_n682__;
  assign new_new_n738__ = ~G54 & new_new_n682__;
  assign new_new_n739__ = ~new_new_n737__ & ~new_new_n738__;
  assign new_new_n740__ = new_new_n584__ & ~new_new_n739__;
  assign new_new_n741__ = ~new_new_n584__ & new_new_n739__;
  assign new_new_n742__ = ~new_new_n740__ & ~new_new_n741__;
  assign new_new_n743__ = new_new_n695__ & ~new_new_n742__;
  assign new_new_n744__ = G52 & new_new_n697__;
  assign new_new_n745__ = ~new_new_n736__ & ~new_new_n744__;
  assign G832 = ~new_new_n743__ & new_new_n745__;
  assign new_new_n747__ = ~new_new_n359__ & new_new_n690__;
  assign new_new_n748__ = ~G54 & new_new_n680__;
  assign new_new_n749__ = new_new_n594__ & ~new_new_n603__;
  assign new_new_n750__ = new_new_n680__ & ~new_new_n749__;
  assign new_new_n751__ = ~new_new_n748__ & ~new_new_n750__;
  assign new_new_n752__ = new_new_n598__ & ~new_new_n751__;
  assign new_new_n753__ = ~new_new_n598__ & new_new_n751__;
  assign new_new_n754__ = ~new_new_n752__ & ~new_new_n753__;
  assign new_new_n755__ = new_new_n695__ & ~new_new_n754__;
  assign new_new_n756__ = G130 & new_new_n697__;
  assign new_new_n757__ = ~new_new_n747__ & ~new_new_n756__;
  assign G834 = ~new_new_n755__ & new_new_n757__;
  assign new_new_n759__ = ~new_new_n377__ & new_new_n690__;
  assign new_new_n760__ = ~new_new_n588__ & new_new_n692__;
  assign new_new_n761__ = ~new_new_n589__ & ~new_new_n760__;
  assign new_new_n762__ = new_new_n604__ & ~new_new_n761__;
  assign new_new_n763__ = ~new_new_n604__ & new_new_n761__;
  assign new_new_n764__ = ~new_new_n762__ & ~new_new_n763__;
  assign new_new_n765__ = new_new_n695__ & ~new_new_n764__;
  assign new_new_n766__ = G119 & new_new_n697__;
  assign new_new_n767__ = ~new_new_n759__ & ~new_new_n766__;
  assign G836 = ~new_new_n765__ & new_new_n767__;
  assign new_new_n769__ = ~G4089 & ~G4090;
  assign new_new_n770__ = ~G822 & new_new_n769__;
  assign new_new_n771__ = G4089 & ~G4090;
  assign new_new_n772__ = ~G861 & new_new_n771__;
  assign new_new_n773__ = ~G11 & ~G4089;
  assign new_new_n774__ = ~G61 & G4089;
  assign new_new_n775__ = G4090 & ~new_new_n773__;
  assign new_new_n776__ = ~new_new_n774__ & new_new_n775__;
  assign new_new_n777__ = ~new_new_n770__ & ~new_new_n776__;
  assign G859 = new_new_n772__ | ~new_new_n777__;
  assign new_new_n779__ = new_new_n422__ & new_new_n690__;
  assign new_new_n780__ = new_new_n542__ & new_new_n554__;
  assign new_new_n781__ = ~new_new_n669__ & ~new_new_n780__;
  assign new_new_n782__ = ~G4 & ~new_new_n669__;
  assign new_new_n783__ = ~new_new_n781__ & ~new_new_n782__;
  assign new_new_n784__ = ~new_new_n546__ & ~new_new_n783__;
  assign new_new_n785__ = ~new_new_n547__ & ~new_new_n784__;
  assign new_new_n786__ = new_new_n529__ & ~new_new_n785__;
  assign new_new_n787__ = ~new_new_n529__ & new_new_n785__;
  assign new_new_n788__ = ~new_new_n786__ & ~new_new_n787__;
  assign new_new_n789__ = new_new_n695__ & ~new_new_n788__;
  assign new_new_n790__ = G122 & new_new_n697__;
  assign new_new_n791__ = ~new_new_n779__ & ~new_new_n790__;
  assign G871 = ~new_new_n789__ & new_new_n791__;
  assign new_new_n793__ = ~new_new_n412__ & new_new_n690__;
  assign new_new_n794__ = ~new_new_n548__ & new_new_n783__;
  assign new_new_n795__ = new_new_n548__ & ~new_new_n783__;
  assign new_new_n796__ = ~new_new_n794__ & ~new_new_n795__;
  assign new_new_n797__ = new_new_n695__ & ~new_new_n796__;
  assign new_new_n798__ = G128 & new_new_n697__;
  assign new_new_n799__ = ~new_new_n793__ & ~new_new_n798__;
  assign G873 = ~new_new_n797__ & new_new_n799__;
  assign new_new_n801__ = ~new_new_n459__ & new_new_n690__;
  assign new_new_n802__ = ~new_new_n533__ & ~new_new_n710__;
  assign new_new_n803__ = new_new_n541__ & ~new_new_n802__;
  assign new_new_n804__ = ~new_new_n539__ & ~new_new_n803__;
  assign new_new_n805__ = new_new_n554__ & ~new_new_n804__;
  assign new_new_n806__ = ~new_new_n554__ & new_new_n804__;
  assign new_new_n807__ = ~new_new_n805__ & ~new_new_n806__;
  assign new_new_n808__ = new_new_n695__ & new_new_n807__;
  assign new_new_n809__ = G127 & new_new_n697__;
  assign new_new_n810__ = ~new_new_n801__ & ~new_new_n809__;
  assign G875 = ~new_new_n808__ & new_new_n810__;
  assign new_new_n812__ = ~new_new_n478__ & new_new_n690__;
  assign new_new_n813__ = ~new_new_n533__ & ~new_new_n541__;
  assign new_new_n814__ = ~new_new_n710__ & new_new_n813__;
  assign new_new_n815__ = ~new_new_n803__ & ~new_new_n814__;
  assign new_new_n816__ = new_new_n695__ & new_new_n815__;
  assign new_new_n817__ = G126 & new_new_n697__;
  assign new_new_n818__ = ~new_new_n812__ & ~new_new_n817__;
  assign G877 = ~new_new_n816__ & new_new_n818__;
  assign new_new_n820__ = new_new_n568__ & ~new_new_n574__;
  assign new_new_n821__ = ~new_new_n568__ & new_new_n574__;
  assign new_new_n822__ = ~new_new_n820__ & ~new_new_n821__;
  assign new_new_n823__ = new_new_n723__ & ~new_new_n822__;
  assign new_new_n824__ = ~new_new_n723__ & new_new_n822__;
  assign new_new_n825__ = ~new_new_n823__ & ~new_new_n824__;
  assign new_new_n826__ = G332 & ~G372;
  assign new_new_n827__ = ~G332 & ~G369;
  assign new_new_n828__ = ~new_new_n826__ & ~new_new_n827__;
  assign new_new_n829__ = new_new_n593__ & ~new_new_n828__;
  assign new_new_n830__ = ~new_new_n593__ & new_new_n828__;
  assign new_new_n831__ = ~new_new_n829__ & ~new_new_n830__;
  assign new_new_n832__ = new_new_n587__ & ~new_new_n831__;
  assign new_new_n833__ = ~new_new_n587__ & new_new_n831__;
  assign new_new_n834__ = ~new_new_n832__ & ~new_new_n833__;
  assign new_new_n835__ = new_new_n601__ & new_new_n834__;
  assign new_new_n836__ = ~new_new_n601__ & ~new_new_n834__;
  assign new_new_n837__ = ~new_new_n835__ & ~new_new_n836__;
  assign new_new_n838__ = new_new_n581__ & ~new_new_n595__;
  assign new_new_n839__ = ~G331 & new_new_n595__;
  assign new_new_n840__ = ~new_new_n838__ & ~new_new_n839__;
  assign new_new_n841__ = new_new_n837__ & ~new_new_n840__;
  assign new_new_n842__ = ~new_new_n837__ & new_new_n840__;
  assign new_new_n843__ = ~new_new_n841__ & ~new_new_n842__;
  assign new_new_n844__ = new_new_n825__ & new_new_n843__;
  assign new_new_n845__ = ~new_new_n825__ & ~new_new_n843__;
  assign G998 = new_new_n844__ | new_new_n845__;
  assign new_new_n847__ = ~new_new_n532__ & new_new_n545__;
  assign new_new_n848__ = new_new_n532__ & ~new_new_n545__;
  assign new_new_n849__ = ~new_new_n847__ & ~new_new_n848__;
  assign new_new_n850__ = ~new_new_n538__ & new_new_n551__;
  assign new_new_n851__ = new_new_n538__ & ~new_new_n551__;
  assign new_new_n852__ = ~new_new_n850__ & ~new_new_n851__;
  assign new_new_n853__ = new_new_n849__ & new_new_n852__;
  assign new_new_n854__ = ~new_new_n849__ & ~new_new_n852__;
  assign new_new_n855__ = ~new_new_n853__ & ~new_new_n854__;
  assign new_new_n856__ = new_new_n526__ & ~new_new_n855__;
  assign new_new_n857__ = ~new_new_n526__ & new_new_n855__;
  assign new_new_n858__ = ~new_new_n856__ & ~new_new_n857__;
  assign new_new_n859__ = G289 & ~G335;
  assign new_new_n860__ = G292 & G335;
  assign new_new_n861__ = ~new_new_n859__ & ~new_new_n860__;
  assign new_new_n862__ = new_new_n505__ & ~new_new_n861__;
  assign new_new_n863__ = ~new_new_n505__ & new_new_n861__;
  assign new_new_n864__ = ~new_new_n862__ & ~new_new_n863__;
  assign new_new_n865__ = new_new_n511__ & new_new_n864__;
  assign new_new_n866__ = ~new_new_n511__ & ~new_new_n864__;
  assign new_new_n867__ = ~new_new_n865__ & ~new_new_n866__;
  assign new_new_n868__ = new_new_n499__ & ~new_new_n519__;
  assign new_new_n869__ = ~new_new_n499__ & new_new_n519__;
  assign new_new_n870__ = ~new_new_n868__ & ~new_new_n869__;
  assign new_new_n871__ = new_new_n867__ & ~new_new_n870__;
  assign new_new_n872__ = ~new_new_n867__ & new_new_n870__;
  assign new_new_n873__ = ~new_new_n871__ & ~new_new_n872__;
  assign new_new_n874__ = new_new_n858__ & new_new_n873__;
  assign new_new_n875__ = ~new_new_n858__ & ~new_new_n873__;
  assign G1000 = new_new_n874__ | new_new_n875__;
  assign new_new_n877__ = G4 & new_new_n557__;
  assign new_new_n878__ = ~new_new_n673__ & ~new_new_n877__;
  assign new_new_n879__ = ~new_new_n500__ & new_new_n878__;
  assign new_new_n880__ = ~new_new_n501__ & ~new_new_n879__;
  assign new_new_n881__ = new_new_n508__ & ~new_new_n880__;
  assign new_new_n882__ = ~new_new_n508__ & new_new_n880__;
  assign new_new_n883__ = ~new_new_n881__ & ~new_new_n882__;
  assign new_new_n884__ = new_new_n516__ & ~new_new_n878__;
  assign new_new_n885__ = ~new_new_n664__ & ~new_new_n884__;
  assign new_new_n886__ = new_new_n522__ & ~new_new_n885__;
  assign new_new_n887__ = ~new_new_n522__ & new_new_n885__;
  assign new_new_n888__ = ~new_new_n886__ & ~new_new_n887__;
  assign new_new_n889__ = new_new_n502__ & ~new_new_n878__;
  assign new_new_n890__ = ~new_new_n502__ & new_new_n878__;
  assign new_new_n891__ = ~new_new_n889__ & ~new_new_n890__;
  assign new_new_n892__ = new_new_n662__ & new_new_n878__;
  assign new_new_n893__ = ~new_new_n501__ & new_new_n508__;
  assign new_new_n894__ = ~new_new_n506__ & ~new_new_n893__;
  assign new_new_n895__ = ~new_new_n892__ & ~new_new_n894__;
  assign new_new_n896__ = new_new_n514__ & ~new_new_n895__;
  assign new_new_n897__ = ~new_new_n514__ & new_new_n895__;
  assign new_new_n898__ = ~new_new_n896__ & ~new_new_n897__;
  assign new_new_n899__ = ~new_new_n712__ & ~new_new_n815__;
  assign new_new_n900__ = ~new_new_n807__ & new_new_n899__;
  assign new_new_n901__ = new_new_n796__ & new_new_n900__;
  assign new_new_n902__ = new_new_n788__ & new_new_n901__;
  assign new_new_n903__ = ~new_new_n891__ & new_new_n902__;
  assign new_new_n904__ = new_new_n883__ & new_new_n903__;
  assign new_new_n905__ = ~new_new_n888__ & new_new_n898__;
  assign G575 = new_new_n904__ & new_new_n905__;
  assign new_new_n907__ = new_new_n577__ & ~new_new_n718__;
  assign new_new_n908__ = ~new_new_n577__ & new_new_n718__;
  assign new_new_n909__ = ~new_new_n907__ & ~new_new_n908__;
  assign new_new_n910__ = ~new_new_n575__ & new_new_n718__;
  assign new_new_n911__ = ~new_new_n576__ & ~new_new_n910__;
  assign new_new_n912__ = new_new_n571__ & ~new_new_n911__;
  assign new_new_n913__ = ~new_new_n571__ & new_new_n911__;
  assign new_new_n914__ = ~new_new_n912__ & ~new_new_n913__;
  assign new_new_n915__ = ~new_new_n564__ & new_new_n720__;
  assign new_new_n916__ = new_new_n564__ & ~new_new_n720__;
  assign new_new_n917__ = ~new_new_n915__ & ~new_new_n916__;
  assign new_new_n918__ = ~new_new_n693__ & new_new_n703__;
  assign new_new_n919__ = new_new_n764__ & new_new_n918__;
  assign new_new_n920__ = new_new_n754__ & new_new_n919__;
  assign new_new_n921__ = new_new_n742__ & new_new_n920__;
  assign new_new_n922__ = ~new_new_n909__ & new_new_n921__;
  assign new_new_n923__ = G623 & new_new_n922__;
  assign new_new_n924__ = new_new_n914__ & new_new_n917__;
  assign G585 = new_new_n923__ & new_new_n924__;
  assign new_new_n926__ = ~G1689 & ~G1690;
  assign new_new_n927__ = ~G822 & new_new_n926__;
  assign new_new_n928__ = G1689 & ~G1690;
  assign new_new_n929__ = ~G861 & new_new_n928__;
  assign new_new_n930__ = ~G182 & ~G1689;
  assign new_new_n931__ = ~G185 & G1689;
  assign new_new_n932__ = G1690 & ~new_new_n930__;
  assign new_new_n933__ = ~new_new_n931__ & new_new_n932__;
  assign new_new_n934__ = ~new_new_n927__ & ~new_new_n933__;
  assign new_new_n935__ = ~new_new_n929__ & new_new_n934__;
  assign G661 = G137 & ~new_new_n935__;
  assign new_new_n937__ = ~G1691 & ~G1694;
  assign new_new_n938__ = ~G822 & new_new_n937__;
  assign new_new_n939__ = G1691 & ~G1694;
  assign new_new_n940__ = ~G861 & new_new_n939__;
  assign new_new_n941__ = ~G182 & ~G1691;
  assign new_new_n942__ = ~G185 & G1691;
  assign new_new_n943__ = G1694 & ~new_new_n941__;
  assign new_new_n944__ = ~new_new_n942__ & new_new_n943__;
  assign new_new_n945__ = ~new_new_n938__ & ~new_new_n944__;
  assign new_new_n946__ = ~new_new_n940__ & new_new_n945__;
  assign G693 = G137 & ~new_new_n946__;
  assign new_new_n948__ = new_new_n728__ & ~G871;
  assign new_new_n949__ = new_new_n726__ & ~G832;
  assign new_new_n950__ = ~G43 & ~G4088;
  assign new_new_n951__ = ~G37 & G4088;
  assign new_new_n952__ = G4087 & ~new_new_n950__;
  assign new_new_n953__ = ~new_new_n951__ & new_new_n952__;
  assign new_new_n954__ = ~new_new_n949__ & ~new_new_n953__;
  assign G747 = new_new_n948__ | ~new_new_n954__;
  assign new_new_n956__ = new_new_n728__ & ~G873;
  assign new_new_n957__ = new_new_n726__ & ~G834;
  assign new_new_n958__ = ~G76 & ~G4088;
  assign new_new_n959__ = ~G20 & G4088;
  assign new_new_n960__ = G4087 & ~new_new_n958__;
  assign new_new_n961__ = ~new_new_n959__ & new_new_n960__;
  assign new_new_n962__ = ~new_new_n957__ & ~new_new_n961__;
  assign G752 = new_new_n956__ | ~new_new_n962__;
  assign new_new_n964__ = new_new_n726__ & ~G836;
  assign new_new_n965__ = new_new_n728__ & ~G875;
  assign new_new_n966__ = ~G73 & ~G4088;
  assign new_new_n967__ = ~G17 & G4088;
  assign new_new_n968__ = G4087 & ~new_new_n966__;
  assign new_new_n969__ = ~new_new_n967__ & new_new_n968__;
  assign new_new_n970__ = ~new_new_n964__ & ~new_new_n969__;
  assign G757 = new_new_n965__ | ~new_new_n970__;
  assign new_new_n972__ = ~G838 & new_new_n726__;
  assign new_new_n973__ = new_new_n728__ & ~G877;
  assign new_new_n974__ = ~G67 & ~G4088;
  assign new_new_n975__ = ~G70 & G4088;
  assign new_new_n976__ = G4087 & ~new_new_n974__;
  assign new_new_n977__ = ~new_new_n975__ & new_new_n976__;
  assign new_new_n978__ = ~new_new_n972__ & ~new_new_n977__;
  assign G762 = new_new_n973__ | ~new_new_n978__;
  assign new_new_n980__ = new_new_n771__ & ~G871;
  assign new_new_n981__ = ~G832 & new_new_n769__;
  assign new_new_n982__ = ~G43 & ~G4089;
  assign new_new_n983__ = ~G37 & G4089;
  assign new_new_n984__ = G4090 & ~new_new_n982__;
  assign new_new_n985__ = ~new_new_n983__ & new_new_n984__;
  assign new_new_n986__ = ~new_new_n981__ & ~new_new_n985__;
  assign G787 = new_new_n980__ | ~new_new_n986__;
  assign new_new_n988__ = new_new_n771__ & ~G873;
  assign new_new_n989__ = ~G834 & new_new_n769__;
  assign new_new_n990__ = ~G76 & ~G4089;
  assign new_new_n991__ = ~G20 & G4089;
  assign new_new_n992__ = G4090 & ~new_new_n990__;
  assign new_new_n993__ = ~new_new_n991__ & new_new_n992__;
  assign new_new_n994__ = ~new_new_n989__ & ~new_new_n993__;
  assign G792 = new_new_n988__ | ~new_new_n994__;
  assign new_new_n996__ = ~G836 & new_new_n769__;
  assign new_new_n997__ = new_new_n771__ & ~G875;
  assign new_new_n998__ = ~G73 & ~G4089;
  assign new_new_n999__ = ~G17 & G4089;
  assign new_new_n1000__ = G4090 & ~new_new_n998__;
  assign new_new_n1001__ = ~new_new_n999__ & new_new_n1000__;
  assign new_new_n1002__ = ~new_new_n996__ & ~new_new_n1001__;
  assign G797 = new_new_n997__ | ~new_new_n1002__;
  assign new_new_n1004__ = ~G838 & new_new_n769__;
  assign new_new_n1005__ = new_new_n771__ & ~G877;
  assign new_new_n1006__ = ~G67 & ~G4089;
  assign new_new_n1007__ = ~G70 & G4089;
  assign new_new_n1008__ = G4090 & ~new_new_n1006__;
  assign new_new_n1009__ = ~new_new_n1007__ & new_new_n1008__;
  assign new_new_n1010__ = ~new_new_n1004__ & ~new_new_n1009__;
  assign G802 = new_new_n1005__ | ~new_new_n1010__;
  assign new_new_n1012__ = ~G871 & new_new_n928__;
  assign new_new_n1013__ = ~G832 & new_new_n926__;
  assign new_new_n1014__ = ~G200 & ~G1689;
  assign new_new_n1015__ = ~G170 & G1689;
  assign new_new_n1016__ = G1690 & ~new_new_n1014__;
  assign new_new_n1017__ = ~new_new_n1015__ & new_new_n1016__;
  assign new_new_n1018__ = ~new_new_n1013__ & ~new_new_n1017__;
  assign new_new_n1019__ = ~new_new_n1012__ & new_new_n1018__;
  assign G642 = G137 & ~new_new_n1019__;
  assign new_new_n1021__ = ~G838 & new_new_n926__;
  assign new_new_n1022__ = ~G877 & new_new_n928__;
  assign new_new_n1023__ = ~G188 & ~G1689;
  assign new_new_n1024__ = ~G158 & G1689;
  assign new_new_n1025__ = G1690 & ~new_new_n1023__;
  assign new_new_n1026__ = ~new_new_n1024__ & new_new_n1025__;
  assign new_new_n1027__ = ~new_new_n1021__ & ~new_new_n1026__;
  assign new_new_n1028__ = ~new_new_n1022__ & new_new_n1027__;
  assign G664 = G137 & ~new_new_n1028__;
  assign new_new_n1030__ = ~G836 & new_new_n926__;
  assign new_new_n1031__ = ~G875 & new_new_n928__;
  assign new_new_n1032__ = ~G155 & ~G1689;
  assign new_new_n1033__ = ~G152 & G1689;
  assign new_new_n1034__ = G1690 & ~new_new_n1032__;
  assign new_new_n1035__ = ~new_new_n1033__ & new_new_n1034__;
  assign new_new_n1036__ = ~new_new_n1030__ & ~new_new_n1035__;
  assign new_new_n1037__ = ~new_new_n1031__ & new_new_n1036__;
  assign G667 = G137 & ~new_new_n1037__;
  assign new_new_n1039__ = ~G873 & new_new_n928__;
  assign new_new_n1040__ = ~G834 & new_new_n926__;
  assign new_new_n1041__ = ~G149 & ~G1689;
  assign new_new_n1042__ = ~G146 & G1689;
  assign new_new_n1043__ = G1690 & ~new_new_n1041__;
  assign new_new_n1044__ = ~new_new_n1042__ & new_new_n1043__;
  assign new_new_n1045__ = ~new_new_n1040__ & ~new_new_n1044__;
  assign new_new_n1046__ = ~new_new_n1039__ & new_new_n1045__;
  assign G670 = G137 & ~new_new_n1046__;
  assign new_new_n1048__ = ~G871 & new_new_n939__;
  assign new_new_n1049__ = ~G832 & new_new_n937__;
  assign new_new_n1050__ = ~G200 & ~G1691;
  assign new_new_n1051__ = ~G170 & G1691;
  assign new_new_n1052__ = G1694 & ~new_new_n1050__;
  assign new_new_n1053__ = ~new_new_n1051__ & new_new_n1052__;
  assign new_new_n1054__ = ~new_new_n1049__ & ~new_new_n1053__;
  assign new_new_n1055__ = ~new_new_n1048__ & new_new_n1054__;
  assign G676 = G137 & ~new_new_n1055__;
  assign new_new_n1057__ = ~G838 & new_new_n937__;
  assign new_new_n1058__ = ~G877 & new_new_n939__;
  assign new_new_n1059__ = ~G188 & ~G1691;
  assign new_new_n1060__ = ~G158 & G1691;
  assign new_new_n1061__ = G1694 & ~new_new_n1059__;
  assign new_new_n1062__ = ~new_new_n1060__ & new_new_n1061__;
  assign new_new_n1063__ = ~new_new_n1057__ & ~new_new_n1062__;
  assign new_new_n1064__ = ~new_new_n1058__ & new_new_n1063__;
  assign G696 = G137 & ~new_new_n1064__;
  assign new_new_n1066__ = ~G836 & new_new_n937__;
  assign new_new_n1067__ = ~G875 & new_new_n939__;
  assign new_new_n1068__ = ~G155 & ~G1691;
  assign new_new_n1069__ = ~G152 & G1691;
  assign new_new_n1070__ = G1694 & ~new_new_n1068__;
  assign new_new_n1071__ = ~new_new_n1069__ & new_new_n1070__;
  assign new_new_n1072__ = ~new_new_n1066__ & ~new_new_n1071__;
  assign new_new_n1073__ = ~new_new_n1067__ & new_new_n1072__;
  assign G699 = G137 & ~new_new_n1073__;
  assign new_new_n1075__ = ~G873 & new_new_n939__;
  assign new_new_n1076__ = ~G834 & new_new_n937__;
  assign new_new_n1077__ = ~G149 & ~G1691;
  assign new_new_n1078__ = ~G146 & G1691;
  assign new_new_n1079__ = G1694 & ~new_new_n1077__;
  assign new_new_n1080__ = ~new_new_n1078__ & new_new_n1079__;
  assign new_new_n1081__ = ~new_new_n1076__ & ~new_new_n1080__;
  assign new_new_n1082__ = ~new_new_n1075__ & new_new_n1081__;
  assign G702 = G137 & ~new_new_n1082__;
  assign new_new_n1084__ = G135 & G4115;
  assign new_new_n1085__ = G3717 & ~G623;
  assign new_new_n1086__ = ~G132 & ~new_new_n561__;
  assign new_new_n1087__ = G132 & new_new_n561__;
  assign new_new_n1088__ = ~new_new_n1086__ & ~new_new_n1087__;
  assign new_new_n1089__ = ~G3717 & ~new_new_n1088__;
  assign new_new_n1090__ = G3724 & ~new_new_n1089__;
  assign new_new_n1091__ = ~new_new_n1085__ & new_new_n1090__;
  assign new_new_n1092__ = ~G3717 & new_new_n353__;
  assign new_new_n1093__ = G123 & G3717;
  assign new_new_n1094__ = ~G3724 & ~new_new_n1093__;
  assign new_new_n1095__ = ~new_new_n1092__ & new_new_n1094__;
  assign new_new_n1096__ = ~new_new_n1084__ & ~new_new_n1095__;
  assign G818 = ~new_new_n1091__ & new_new_n1096__;
  assign new_new_n1098__ = ~G132 & ~new_new_n915__;
  assign new_new_n1099__ = G132 & new_new_n915__;
  assign G813 = new_new_n1098__ | new_new_n1099__;
  assign new_new_n1101__ = new_new_n353__ & new_new_n690__;
  assign new_new_n1102__ = G123 & new_new_n697__;
  assign new_new_n1103__ = new_new_n695__ & ~G623;
  assign new_new_n1104__ = ~new_new_n1101__ & ~new_new_n1102__;
  assign G824 = ~new_new_n1103__ & new_new_n1104__;
  assign new_new_n1106__ = ~new_new_n350__ & new_new_n690__;
  assign new_new_n1107__ = new_new_n695__ & ~new_new_n917__;
  assign new_new_n1108__ = G121 & new_new_n697__;
  assign new_new_n1109__ = ~new_new_n1106__ & ~new_new_n1108__;
  assign G826 = ~new_new_n1107__ & new_new_n1109__;
  assign new_new_n1111__ = ~new_new_n395__ & new_new_n690__;
  assign new_new_n1112__ = new_new_n695__ & ~new_new_n914__;
  assign new_new_n1113__ = G116 & new_new_n697__;
  assign new_new_n1114__ = ~new_new_n1111__ & ~new_new_n1113__;
  assign G828 = ~new_new_n1112__ & new_new_n1114__;
  assign new_new_n1116__ = ~new_new_n386__ & new_new_n690__;
  assign new_new_n1117__ = new_new_n695__ & new_new_n909__;
  assign new_new_n1118__ = G112 & new_new_n697__;
  assign new_new_n1119__ = ~new_new_n1116__ & ~new_new_n1118__;
  assign G830 = ~new_new_n1117__ & new_new_n1119__;
  assign new_new_n1121__ = G245 & G559;
  assign new_new_n1122__ = G601 & new_new_n1121__;
  assign new_new_n1123__ = ~G847 & new_new_n1122__;
  assign new_new_n1124__ = ~G1002 & new_new_n1123__;
  assign new_new_n1125__ = ~G1004 & new_new_n1124__;
  assign new_new_n1126__ = ~G1000 & new_new_n1125__;
  assign G854 = ~G998 & new_new_n1126__;
  assign new_new_n1128__ = ~new_new_n431__ & new_new_n690__;
  assign new_new_n1129__ = new_new_n695__ & new_new_n888__;
  assign new_new_n1130__ = G115 & new_new_n697__;
  assign new_new_n1131__ = ~new_new_n1128__ & ~new_new_n1130__;
  assign G863 = ~new_new_n1129__ & new_new_n1131__;
  assign new_new_n1133__ = new_new_n469__ & new_new_n690__;
  assign new_new_n1134__ = new_new_n695__ & ~new_new_n898__;
  assign new_new_n1135__ = G114 & new_new_n697__;
  assign new_new_n1136__ = ~new_new_n1133__ & ~new_new_n1135__;
  assign G865 = ~new_new_n1134__ & new_new_n1136__;
  assign new_new_n1138__ = new_new_n488__ & new_new_n690__;
  assign new_new_n1139__ = new_new_n695__ & ~new_new_n883__;
  assign new_new_n1140__ = G53 & new_new_n697__;
  assign new_new_n1141__ = ~new_new_n1138__ & ~new_new_n1140__;
  assign G867 = ~new_new_n1139__ & new_new_n1141__;
  assign new_new_n1143__ = new_new_n441__ & new_new_n690__;
  assign new_new_n1144__ = new_new_n695__ & new_new_n891__;
  assign new_new_n1145__ = G113 & new_new_n697__;
  assign new_new_n1146__ = ~new_new_n1143__ & ~new_new_n1145__;
  assign G869 = ~new_new_n1144__ & new_new_n1146__;
  assign new_new_n1148__ = new_new_n771__ & ~G863;
  assign new_new_n1149__ = new_new_n769__ & ~G824;
  assign new_new_n1150__ = ~G109 & ~G4089;
  assign new_new_n1151__ = ~G106 & G4089;
  assign new_new_n1152__ = G4090 & ~new_new_n1150__;
  assign new_new_n1153__ = ~new_new_n1151__ & new_new_n1152__;
  assign new_new_n1154__ = ~new_new_n1149__ & ~new_new_n1153__;
  assign G712 = new_new_n1148__ | ~new_new_n1154__;
  assign new_new_n1156__ = new_new_n728__ & ~G863;
  assign new_new_n1157__ = new_new_n726__ & ~G824;
  assign new_new_n1158__ = ~G109 & ~G4088;
  assign new_new_n1159__ = ~G106 & G4088;
  assign new_new_n1160__ = G4087 & ~new_new_n1158__;
  assign new_new_n1161__ = ~new_new_n1159__ & new_new_n1160__;
  assign new_new_n1162__ = ~new_new_n1157__ & ~new_new_n1161__;
  assign G727 = new_new_n1156__ | ~new_new_n1162__;
  assign new_new_n1164__ = new_new_n728__ & ~G865;
  assign new_new_n1165__ = new_new_n726__ & ~G826;
  assign new_new_n1166__ = ~G46 & ~G4088;
  assign new_new_n1167__ = ~G49 & G4088;
  assign new_new_n1168__ = G4087 & ~new_new_n1166__;
  assign new_new_n1169__ = ~new_new_n1167__ & new_new_n1168__;
  assign new_new_n1170__ = ~new_new_n1165__ & ~new_new_n1169__;
  assign G732 = new_new_n1164__ | ~new_new_n1170__;
  assign new_new_n1172__ = new_new_n728__ & ~G867;
  assign new_new_n1173__ = new_new_n726__ & ~G828;
  assign new_new_n1174__ = ~G100 & ~G4088;
  assign new_new_n1175__ = ~G103 & G4088;
  assign new_new_n1176__ = G4087 & ~new_new_n1174__;
  assign new_new_n1177__ = ~new_new_n1175__ & new_new_n1176__;
  assign new_new_n1178__ = ~new_new_n1173__ & ~new_new_n1177__;
  assign G737 = new_new_n1172__ | ~new_new_n1178__;
  assign new_new_n1180__ = new_new_n728__ & ~G869;
  assign new_new_n1181__ = new_new_n726__ & ~G830;
  assign new_new_n1182__ = ~G91 & ~G4088;
  assign new_new_n1183__ = ~G40 & G4088;
  assign new_new_n1184__ = G4087 & ~new_new_n1182__;
  assign new_new_n1185__ = ~new_new_n1183__ & new_new_n1184__;
  assign new_new_n1186__ = ~new_new_n1181__ & ~new_new_n1185__;
  assign G742 = new_new_n1180__ | ~new_new_n1186__;
  assign new_new_n1188__ = new_new_n771__ & ~G865;
  assign new_new_n1189__ = new_new_n769__ & ~G826;
  assign new_new_n1190__ = ~G46 & ~G4089;
  assign new_new_n1191__ = ~G49 & G4089;
  assign new_new_n1192__ = G4090 & ~new_new_n1190__;
  assign new_new_n1193__ = ~new_new_n1191__ & new_new_n1192__;
  assign new_new_n1194__ = ~new_new_n1189__ & ~new_new_n1193__;
  assign G772 = new_new_n1188__ | ~new_new_n1194__;
  assign new_new_n1196__ = new_new_n771__ & ~G867;
  assign new_new_n1197__ = new_new_n769__ & ~G828;
  assign new_new_n1198__ = ~G100 & ~G4089;
  assign new_new_n1199__ = ~G103 & G4089;
  assign new_new_n1200__ = G4090 & ~new_new_n1198__;
  assign new_new_n1201__ = ~new_new_n1199__ & new_new_n1200__;
  assign new_new_n1202__ = ~new_new_n1197__ & ~new_new_n1201__;
  assign G777 = new_new_n1196__ | ~new_new_n1202__;
  assign new_new_n1204__ = new_new_n771__ & ~G869;
  assign new_new_n1205__ = new_new_n769__ & ~G830;
  assign new_new_n1206__ = ~G91 & ~G4089;
  assign new_new_n1207__ = ~G40 & G4089;
  assign new_new_n1208__ = G4090 & ~new_new_n1206__;
  assign new_new_n1209__ = ~new_new_n1207__ & new_new_n1208__;
  assign new_new_n1210__ = ~new_new_n1205__ & ~new_new_n1209__;
  assign G782 = new_new_n1204__ | ~new_new_n1210__;
  assign new_new_n1212__ = new_new_n928__ & ~G869;
  assign new_new_n1213__ = new_new_n926__ & ~G830;
  assign new_new_n1214__ = ~G203 & ~G1689;
  assign new_new_n1215__ = ~G173 & G1689;
  assign new_new_n1216__ = G1690 & ~new_new_n1214__;
  assign new_new_n1217__ = ~new_new_n1215__ & new_new_n1216__;
  assign new_new_n1218__ = ~new_new_n1213__ & ~new_new_n1217__;
  assign new_new_n1219__ = ~new_new_n1212__ & new_new_n1218__;
  assign G645 = G137 & ~new_new_n1219__;
  assign new_new_n1221__ = new_new_n928__ & ~G867;
  assign new_new_n1222__ = new_new_n926__ & ~G828;
  assign new_new_n1223__ = ~G197 & ~G1689;
  assign new_new_n1224__ = ~G167 & G1689;
  assign new_new_n1225__ = G1690 & ~new_new_n1223__;
  assign new_new_n1226__ = ~new_new_n1224__ & new_new_n1225__;
  assign new_new_n1227__ = ~new_new_n1222__ & ~new_new_n1226__;
  assign new_new_n1228__ = ~new_new_n1221__ & new_new_n1227__;
  assign G648 = G137 & ~new_new_n1228__;
  assign new_new_n1230__ = new_new_n928__ & ~G865;
  assign new_new_n1231__ = new_new_n926__ & ~G826;
  assign new_new_n1232__ = ~G194 & ~G1689;
  assign new_new_n1233__ = ~G164 & G1689;
  assign new_new_n1234__ = G1690 & ~new_new_n1232__;
  assign new_new_n1235__ = ~new_new_n1233__ & new_new_n1234__;
  assign new_new_n1236__ = ~new_new_n1231__ & ~new_new_n1235__;
  assign new_new_n1237__ = ~new_new_n1230__ & new_new_n1236__;
  assign G651 = G137 & ~new_new_n1237__;
  assign new_new_n1239__ = new_new_n928__ & ~G863;
  assign new_new_n1240__ = new_new_n926__ & ~G824;
  assign new_new_n1241__ = ~G191 & ~G1689;
  assign new_new_n1242__ = ~G161 & G1689;
  assign new_new_n1243__ = G1690 & ~new_new_n1241__;
  assign new_new_n1244__ = ~new_new_n1242__ & new_new_n1243__;
  assign new_new_n1245__ = ~new_new_n1240__ & ~new_new_n1244__;
  assign new_new_n1246__ = ~new_new_n1239__ & new_new_n1245__;
  assign G654 = G137 & ~new_new_n1246__;
  assign new_new_n1248__ = new_new_n939__ & ~G869;
  assign new_new_n1249__ = new_new_n937__ & ~G830;
  assign new_new_n1250__ = ~G203 & ~G1691;
  assign new_new_n1251__ = ~G173 & G1691;
  assign new_new_n1252__ = G1694 & ~new_new_n1250__;
  assign new_new_n1253__ = ~new_new_n1251__ & new_new_n1252__;
  assign new_new_n1254__ = ~new_new_n1249__ & ~new_new_n1253__;
  assign new_new_n1255__ = ~new_new_n1248__ & new_new_n1254__;
  assign G679 = G137 & ~new_new_n1255__;
  assign new_new_n1257__ = new_new_n939__ & ~G867;
  assign new_new_n1258__ = new_new_n937__ & ~G828;
  assign new_new_n1259__ = ~G197 & ~G1691;
  assign new_new_n1260__ = ~G167 & G1691;
  assign new_new_n1261__ = G1694 & ~new_new_n1259__;
  assign new_new_n1262__ = ~new_new_n1260__ & new_new_n1261__;
  assign new_new_n1263__ = ~new_new_n1258__ & ~new_new_n1262__;
  assign new_new_n1264__ = ~new_new_n1257__ & new_new_n1263__;
  assign G682 = G137 & ~new_new_n1264__;
  assign new_new_n1266__ = new_new_n939__ & ~G865;
  assign new_new_n1267__ = new_new_n937__ & ~G826;
  assign new_new_n1268__ = ~G194 & ~G1691;
  assign new_new_n1269__ = ~G164 & G1691;
  assign new_new_n1270__ = G1694 & ~new_new_n1268__;
  assign new_new_n1271__ = ~new_new_n1269__ & new_new_n1270__;
  assign new_new_n1272__ = ~new_new_n1267__ & ~new_new_n1271__;
  assign new_new_n1273__ = ~new_new_n1266__ & new_new_n1272__;
  assign G685 = G137 & ~new_new_n1273__;
  assign new_new_n1275__ = new_new_n939__ & ~G863;
  assign new_new_n1276__ = new_new_n937__ & ~G824;
  assign new_new_n1277__ = ~G191 & ~G1691;
  assign new_new_n1278__ = ~G161 & G1691;
  assign new_new_n1279__ = G1694 & ~new_new_n1277__;
  assign new_new_n1280__ = ~new_new_n1278__ & new_new_n1279__;
  assign new_new_n1281__ = ~new_new_n1276__ & ~new_new_n1280__;
  assign new_new_n1282__ = ~new_new_n1275__ & new_new_n1281__;
  assign G688 = G137 & ~new_new_n1282__;
  assign new_new_n1284__ = ~G120 & ~G4091;
  assign new_new_n1285__ = ~new_new_n350__ & new_new_n353__;
  assign new_new_n1286__ = ~new_new_n397__ & ~new_new_n1285__;
  assign new_new_n1287__ = G251 & ~G351;
  assign new_new_n1288__ = G248 & G351;
  assign new_new_n1289__ = G534 & ~new_new_n1287__;
  assign new_new_n1290__ = ~new_new_n1288__ & new_new_n1289__;
  assign new_new_n1291__ = ~G254 & ~G351;
  assign new_new_n1292__ = ~G242 & G351;
  assign new_new_n1293__ = ~G534 & ~new_new_n1291__;
  assign new_new_n1294__ = ~new_new_n1292__ & new_new_n1293__;
  assign new_new_n1295__ = ~new_new_n1290__ & ~new_new_n1294__;
  assign new_new_n1296__ = G251 & ~G341;
  assign new_new_n1297__ = G248 & G341;
  assign new_new_n1298__ = G523 & ~new_new_n1296__;
  assign new_new_n1299__ = ~new_new_n1297__ & new_new_n1298__;
  assign new_new_n1300__ = ~G254 & ~G341;
  assign new_new_n1301__ = ~G242 & G341;
  assign new_new_n1302__ = ~G523 & ~new_new_n1300__;
  assign new_new_n1303__ = ~new_new_n1301__ & new_new_n1302__;
  assign new_new_n1304__ = ~new_new_n1299__ & ~new_new_n1303__;
  assign new_new_n1305__ = ~new_new_n1295__ & new_new_n1304__;
  assign new_new_n1306__ = new_new_n1295__ & ~new_new_n1304__;
  assign new_new_n1307__ = ~new_new_n1305__ & ~new_new_n1306__;
  assign new_new_n1308__ = ~G248 & G514;
  assign new_new_n1309__ = G242 & ~G514;
  assign new_new_n1310__ = ~new_new_n1308__ & ~new_new_n1309__;
  assign new_new_n1311__ = new_new_n1307__ & ~new_new_n1310__;
  assign new_new_n1312__ = ~new_new_n1307__ & new_new_n1310__;
  assign new_new_n1313__ = ~new_new_n1311__ & ~new_new_n1312__;
  assign new_new_n1314__ = ~new_new_n386__ & ~new_new_n395__;
  assign new_new_n1315__ = ~new_new_n396__ & ~new_new_n1314__;
  assign new_new_n1316__ = G251 & ~G324;
  assign new_new_n1317__ = G248 & G324;
  assign new_new_n1318__ = G503 & ~new_new_n1316__;
  assign new_new_n1319__ = ~new_new_n1317__ & new_new_n1318__;
  assign new_new_n1320__ = ~G254 & ~G324;
  assign new_new_n1321__ = ~G242 & G324;
  assign new_new_n1322__ = ~G503 & ~new_new_n1320__;
  assign new_new_n1323__ = ~new_new_n1321__ & new_new_n1322__;
  assign new_new_n1324__ = ~new_new_n1319__ & ~new_new_n1323__;
  assign new_new_n1325__ = ~new_new_n356__ & new_new_n1324__;
  assign new_new_n1326__ = new_new_n356__ & ~new_new_n1324__;
  assign new_new_n1327__ = ~new_new_n1325__ & ~new_new_n1326__;
  assign new_new_n1328__ = new_new_n1315__ & ~new_new_n1327__;
  assign new_new_n1329__ = ~new_new_n1315__ & new_new_n1327__;
  assign new_new_n1330__ = ~new_new_n1328__ & ~new_new_n1329__;
  assign new_new_n1331__ = ~new_new_n1313__ & new_new_n1330__;
  assign new_new_n1332__ = new_new_n1313__ & ~new_new_n1330__;
  assign new_new_n1333__ = ~new_new_n1331__ & ~new_new_n1332__;
  assign new_new_n1334__ = new_new_n1286__ & new_new_n1333__;
  assign new_new_n1335__ = ~new_new_n1286__ & ~new_new_n1333__;
  assign new_new_n1336__ = ~G4091 & ~new_new_n1334__;
  assign new_new_n1337__ = ~new_new_n1335__ & new_new_n1336__;
  assign new_new_n1338__ = ~G4092 & ~new_new_n1337__;
  assign new_new_n1339__ = ~new_new_n1284__ & ~new_new_n1338__;
  assign new_new_n1340__ = G4092 & ~new_new_n1339__;
  assign new_new_n1341__ = G2174 & new_new_n607__;
  assign new_new_n1342__ = new_new_n684__ & ~new_new_n1341__;
  assign new_new_n1343__ = new_new_n564__ & new_new_n570__;
  assign new_new_n1344__ = new_new_n564__ & new_new_n686__;
  assign new_new_n1345__ = new_new_n571__ & ~new_new_n1344__;
  assign new_new_n1346__ = ~new_new_n1343__ & ~new_new_n1345__;
  assign new_new_n1347__ = ~new_new_n575__ & ~new_new_n1346__;
  assign new_new_n1348__ = new_new_n575__ & new_new_n1346__;
  assign new_new_n1349__ = ~new_new_n578__ & ~new_new_n1347__;
  assign new_new_n1350__ = ~new_new_n1348__ & new_new_n1349__;
  assign new_new_n1351__ = ~new_new_n1342__ & ~new_new_n1350__;
  assign new_new_n1352__ = new_new_n576__ & ~new_new_n1346__;
  assign new_new_n1353__ = ~new_new_n576__ & new_new_n1346__;
  assign new_new_n1354__ = ~new_new_n1352__ & ~new_new_n1353__;
  assign new_new_n1355__ = new_new_n1342__ & new_new_n1354__;
  assign new_new_n1356__ = ~new_new_n1351__ & ~new_new_n1355__;
  assign new_new_n1357__ = ~new_new_n598__ & ~new_new_n604__;
  assign new_new_n1358__ = ~new_new_n605__ & ~new_new_n1357__;
  assign new_new_n1359__ = new_new_n584__ & ~new_new_n750__;
  assign new_new_n1360__ = ~new_new_n584__ & new_new_n750__;
  assign new_new_n1361__ = ~new_new_n1359__ & ~new_new_n1360__;
  assign new_new_n1362__ = ~new_new_n588__ & new_new_n593__;
  assign new_new_n1363__ = new_new_n588__ & ~new_new_n593__;
  assign new_new_n1364__ = ~new_new_n1362__ & ~new_new_n1363__;
  assign new_new_n1365__ = new_new_n737__ & ~new_new_n1364__;
  assign new_new_n1366__ = ~new_new_n737__ & new_new_n1364__;
  assign new_new_n1367__ = ~new_new_n1365__ & ~new_new_n1366__;
  assign new_new_n1368__ = new_new_n1361__ & ~new_new_n1367__;
  assign new_new_n1369__ = ~new_new_n1361__ & new_new_n1367__;
  assign new_new_n1370__ = G2174 & ~new_new_n1368__;
  assign new_new_n1371__ = ~new_new_n1369__ & new_new_n1370__;
  assign new_new_n1372__ = ~new_new_n584__ & new_new_n682__;
  assign new_new_n1373__ = ~new_new_n683__ & ~new_new_n1372__;
  assign new_new_n1374__ = ~new_new_n589__ & ~new_new_n1362__;
  assign new_new_n1375__ = new_new_n680__ & ~new_new_n1374__;
  assign new_new_n1376__ = ~new_new_n680__ & new_new_n1374__;
  assign new_new_n1377__ = ~new_new_n1375__ & ~new_new_n1376__;
  assign new_new_n1378__ = new_new_n1373__ & new_new_n1377__;
  assign new_new_n1379__ = ~new_new_n1373__ & ~new_new_n1377__;
  assign new_new_n1380__ = ~G2174 & ~new_new_n1378__;
  assign new_new_n1381__ = ~new_new_n1379__ & new_new_n1380__;
  assign new_new_n1382__ = ~new_new_n1371__ & ~new_new_n1381__;
  assign new_new_n1383__ = new_new_n723__ & ~new_new_n1382__;
  assign new_new_n1384__ = ~new_new_n723__ & new_new_n1382__;
  assign new_new_n1385__ = ~new_new_n1383__ & ~new_new_n1384__;
  assign new_new_n1386__ = ~new_new_n1358__ & new_new_n1385__;
  assign new_new_n1387__ = new_new_n1358__ & ~new_new_n1385__;
  assign new_new_n1388__ = ~new_new_n1386__ & ~new_new_n1387__;
  assign new_new_n1389__ = new_new_n1356__ & new_new_n1388__;
  assign new_new_n1390__ = ~new_new_n1356__ & ~new_new_n1388__;
  assign new_new_n1391__ = G4091 & ~new_new_n1389__;
  assign new_new_n1392__ = ~new_new_n1390__ & new_new_n1391__;
  assign new_new_n1393__ = new_new_n1338__ & ~new_new_n1392__;
  assign G843 = ~new_new_n1340__ & ~new_new_n1393__;
  assign new_new_n1395__ = ~G118 & ~G4091;
  assign new_new_n1396__ = G251 & ~G257;
  assign new_new_n1397__ = G248 & G257;
  assign new_new_n1398__ = G389 & ~new_new_n1396__;
  assign new_new_n1399__ = ~new_new_n1397__ & new_new_n1398__;
  assign new_new_n1400__ = ~G254 & ~G257;
  assign new_new_n1401__ = ~G242 & G257;
  assign new_new_n1402__ = ~G389 & ~new_new_n1400__;
  assign new_new_n1403__ = ~new_new_n1401__ & new_new_n1402__;
  assign new_new_n1404__ = ~new_new_n1399__ & ~new_new_n1403__;
  assign new_new_n1405__ = G251 & ~G281;
  assign new_new_n1406__ = G248 & G281;
  assign new_new_n1407__ = G374 & ~new_new_n1405__;
  assign new_new_n1408__ = ~new_new_n1406__ & new_new_n1407__;
  assign new_new_n1409__ = ~G254 & ~G281;
  assign new_new_n1410__ = ~G242 & G281;
  assign new_new_n1411__ = ~G374 & ~new_new_n1409__;
  assign new_new_n1412__ = ~new_new_n1410__ & new_new_n1411__;
  assign new_new_n1413__ = ~new_new_n1408__ & ~new_new_n1412__;
  assign new_new_n1414__ = ~new_new_n1404__ & new_new_n1413__;
  assign new_new_n1415__ = new_new_n1404__ & ~new_new_n1413__;
  assign new_new_n1416__ = ~new_new_n1414__ & ~new_new_n1415__;
  assign new_new_n1417__ = G248 & new_new_n432__;
  assign new_new_n1418__ = G251 & new_new_n434__;
  assign new_new_n1419__ = ~G226 & G254;
  assign new_new_n1420__ = G226 & G242;
  assign new_new_n1421__ = ~G422 & ~new_new_n1419__;
  assign new_new_n1422__ = ~new_new_n1420__ & new_new_n1421__;
  assign new_new_n1423__ = ~new_new_n1417__ & ~new_new_n1418__;
  assign new_new_n1424__ = ~new_new_n1422__ & new_new_n1423__;
  assign new_new_n1425__ = new_new_n431__ & ~new_new_n1424__;
  assign new_new_n1426__ = ~new_new_n431__ & new_new_n1424__;
  assign new_new_n1427__ = ~new_new_n1425__ & ~new_new_n1426__;
  assign new_new_n1428__ = new_new_n1416__ & ~new_new_n1427__;
  assign new_new_n1429__ = ~new_new_n1416__ & new_new_n1427__;
  assign new_new_n1430__ = ~new_new_n1428__ & ~new_new_n1429__;
  assign new_new_n1431__ = G251 & ~G273;
  assign new_new_n1432__ = G248 & G273;
  assign new_new_n1433__ = G411 & ~new_new_n1431__;
  assign new_new_n1434__ = ~new_new_n1432__ & new_new_n1433__;
  assign new_new_n1435__ = ~G254 & ~G273;
  assign new_new_n1436__ = ~G242 & G273;
  assign new_new_n1437__ = ~G411 & ~new_new_n1435__;
  assign new_new_n1438__ = ~new_new_n1436__ & new_new_n1437__;
  assign new_new_n1439__ = ~new_new_n1434__ & ~new_new_n1438__;
  assign new_new_n1440__ = G251 & ~G265;
  assign new_new_n1441__ = G248 & G265;
  assign new_new_n1442__ = G400 & ~new_new_n1440__;
  assign new_new_n1443__ = ~new_new_n1441__ & new_new_n1442__;
  assign new_new_n1444__ = ~G254 & ~G265;
  assign new_new_n1445__ = ~G242 & G265;
  assign new_new_n1446__ = ~G400 & ~new_new_n1444__;
  assign new_new_n1447__ = ~new_new_n1445__ & new_new_n1446__;
  assign new_new_n1448__ = ~new_new_n1443__ & ~new_new_n1447__;
  assign new_new_n1449__ = ~new_new_n1439__ & new_new_n1448__;
  assign new_new_n1450__ = new_new_n1439__ & ~new_new_n1448__;
  assign new_new_n1451__ = ~new_new_n1449__ & ~new_new_n1450__;
  assign new_new_n1452__ = G248 & new_new_n413__;
  assign new_new_n1453__ = G251 & new_new_n415__;
  assign new_new_n1454__ = ~G234 & G254;
  assign new_new_n1455__ = G234 & G242;
  assign new_new_n1456__ = ~G435 & ~new_new_n1454__;
  assign new_new_n1457__ = ~new_new_n1455__ & new_new_n1456__;
  assign new_new_n1458__ = ~new_new_n1452__ & ~new_new_n1453__;
  assign new_new_n1459__ = ~new_new_n1457__ & new_new_n1458__;
  assign new_new_n1460__ = new_new_n1451__ & new_new_n1459__;
  assign new_new_n1461__ = ~new_new_n1451__ & ~new_new_n1459__;
  assign new_new_n1462__ = ~new_new_n1460__ & ~new_new_n1461__;
  assign new_new_n1463__ = G248 & new_new_n460__;
  assign new_new_n1464__ = G251 & new_new_n462__;
  assign new_new_n1465__ = ~G210 & G254;
  assign new_new_n1466__ = G210 & G242;
  assign new_new_n1467__ = ~G457 & ~new_new_n1465__;
  assign new_new_n1468__ = ~new_new_n1466__ & new_new_n1467__;
  assign new_new_n1469__ = ~new_new_n1463__ & ~new_new_n1464__;
  assign new_new_n1470__ = ~new_new_n1468__ & new_new_n1469__;
  assign new_new_n1471__ = G248 & new_new_n479__;
  assign new_new_n1472__ = G251 & new_new_n481__;
  assign new_new_n1473__ = ~G218 & G254;
  assign new_new_n1474__ = G218 & G242;
  assign new_new_n1475__ = ~G468 & ~new_new_n1473__;
  assign new_new_n1476__ = ~new_new_n1474__ & new_new_n1475__;
  assign new_new_n1477__ = ~new_new_n1471__ & ~new_new_n1472__;
  assign new_new_n1478__ = ~new_new_n1476__ & new_new_n1477__;
  assign new_new_n1479__ = new_new_n1470__ & ~new_new_n1478__;
  assign new_new_n1480__ = ~new_new_n1470__ & new_new_n1478__;
  assign new_new_n1481__ = ~new_new_n1479__ & ~new_new_n1480__;
  assign new_new_n1482__ = new_new_n1462__ & ~new_new_n1481__;
  assign new_new_n1483__ = ~new_new_n1462__ & new_new_n1481__;
  assign new_new_n1484__ = ~new_new_n1482__ & ~new_new_n1483__;
  assign new_new_n1485__ = new_new_n1430__ & ~new_new_n1484__;
  assign new_new_n1486__ = ~new_new_n1430__ & new_new_n1484__;
  assign new_new_n1487__ = ~G4091 & ~new_new_n1485__;
  assign new_new_n1488__ = ~new_new_n1486__ & new_new_n1487__;
  assign new_new_n1489__ = ~G4092 & ~new_new_n1488__;
  assign new_new_n1490__ = ~new_new_n1395__ & ~new_new_n1489__;
  assign new_new_n1491__ = G4092 & ~new_new_n1490__;
  assign new_new_n1492__ = ~new_new_n548__ & ~new_new_n554__;
  assign new_new_n1493__ = ~new_new_n555__ & ~new_new_n1492__;
  assign new_new_n1494__ = new_new_n514__ & ~new_new_n1493__;
  assign new_new_n1495__ = ~new_new_n514__ & new_new_n1493__;
  assign new_new_n1496__ = ~new_new_n1494__ & ~new_new_n1495__;
  assign new_new_n1497__ = G1497 & new_new_n557__;
  assign new_new_n1498__ = ~new_new_n673__ & ~new_new_n1497__;
  assign new_new_n1499__ = ~new_new_n513__ & ~new_new_n662__;
  assign new_new_n1500__ = ~new_new_n663__ & ~new_new_n1499__;
  assign new_new_n1501__ = new_new_n522__ & ~new_new_n1500__;
  assign new_new_n1502__ = ~new_new_n522__ & new_new_n1500__;
  assign new_new_n1503__ = ~new_new_n1501__ & ~new_new_n1502__;
  assign new_new_n1504__ = new_new_n501__ & ~new_new_n508__;
  assign new_new_n1505__ = ~new_new_n893__ & ~new_new_n1504__;
  assign new_new_n1506__ = new_new_n1503__ & new_new_n1505__;
  assign new_new_n1507__ = ~new_new_n1503__ & ~new_new_n1505__;
  assign new_new_n1508__ = ~new_new_n1506__ & ~new_new_n1507__;
  assign new_new_n1509__ = new_new_n1498__ & new_new_n1508__;
  assign new_new_n1510__ = ~new_new_n500__ & ~new_new_n508__;
  assign new_new_n1511__ = ~new_new_n661__ & ~new_new_n1510__;
  assign new_new_n1512__ = ~new_new_n513__ & ~new_new_n894__;
  assign new_new_n1513__ = ~new_new_n664__ & new_new_n894__;
  assign new_new_n1514__ = ~new_new_n1512__ & ~new_new_n1513__;
  assign new_new_n1515__ = ~new_new_n522__ & ~new_new_n1514__;
  assign new_new_n1516__ = new_new_n522__ & new_new_n1514__;
  assign new_new_n1517__ = ~new_new_n1515__ & ~new_new_n1516__;
  assign new_new_n1518__ = new_new_n1511__ & new_new_n1517__;
  assign new_new_n1519__ = ~new_new_n1511__ & ~new_new_n1517__;
  assign new_new_n1520__ = ~new_new_n1498__ & ~new_new_n1518__;
  assign new_new_n1521__ = ~new_new_n1519__ & new_new_n1520__;
  assign new_new_n1522__ = ~new_new_n1509__ & ~new_new_n1521__;
  assign new_new_n1523__ = ~new_new_n539__ & ~new_new_n666__;
  assign new_new_n1524__ = ~new_new_n542__ & new_new_n1523__;
  assign new_new_n1525__ = new_new_n529__ & ~new_new_n1524__;
  assign new_new_n1526__ = ~new_new_n529__ & new_new_n1524__;
  assign new_new_n1527__ = ~new_new_n1525__ & ~new_new_n1526__;
  assign new_new_n1528__ = ~new_new_n666__ & ~new_new_n813__;
  assign new_new_n1529__ = ~new_new_n546__ & new_new_n781__;
  assign new_new_n1530__ = ~new_new_n556__ & ~new_new_n671__;
  assign new_new_n1531__ = ~new_new_n781__ & ~new_new_n1530__;
  assign new_new_n1532__ = ~new_new_n1529__ & ~new_new_n1531__;
  assign new_new_n1533__ = new_new_n1528__ & ~new_new_n1532__;
  assign new_new_n1534__ = ~new_new_n1528__ & new_new_n1532__;
  assign new_new_n1535__ = ~new_new_n1533__ & ~new_new_n1534__;
  assign new_new_n1536__ = new_new_n1527__ & ~new_new_n1535__;
  assign new_new_n1537__ = ~new_new_n1527__ & new_new_n1535__;
  assign new_new_n1538__ = ~new_new_n1536__ & ~new_new_n1537__;
  assign new_new_n1539__ = G1497 & ~new_new_n1538__;
  assign new_new_n1540__ = new_new_n541__ & ~new_new_n671__;
  assign new_new_n1541__ = ~new_new_n541__ & new_new_n671__;
  assign new_new_n1542__ = ~new_new_n1540__ & ~new_new_n1541__;
  assign new_new_n1543__ = new_new_n533__ & ~new_new_n669__;
  assign new_new_n1544__ = ~new_new_n533__ & ~new_new_n553__;
  assign new_new_n1545__ = ~new_new_n667__ & new_new_n1544__;
  assign new_new_n1546__ = new_new_n535__ & ~new_new_n1545__;
  assign new_new_n1547__ = ~new_new_n535__ & new_new_n1545__;
  assign new_new_n1548__ = ~new_new_n1546__ & ~new_new_n1547__;
  assign new_new_n1549__ = ~new_new_n1543__ & new_new_n1548__;
  assign new_new_n1550__ = new_new_n529__ & ~new_new_n1523__;
  assign new_new_n1551__ = ~new_new_n529__ & new_new_n1523__;
  assign new_new_n1552__ = ~new_new_n1550__ & ~new_new_n1551__;
  assign new_new_n1553__ = ~new_new_n1549__ & new_new_n1552__;
  assign new_new_n1554__ = new_new_n1549__ & ~new_new_n1552__;
  assign new_new_n1555__ = ~new_new_n1553__ & ~new_new_n1554__;
  assign new_new_n1556__ = new_new_n1542__ & new_new_n1555__;
  assign new_new_n1557__ = ~new_new_n1542__ & ~new_new_n1555__;
  assign new_new_n1558__ = ~new_new_n1556__ & ~new_new_n1557__;
  assign new_new_n1559__ = ~G1497 & ~new_new_n1558__;
  assign new_new_n1560__ = ~new_new_n1539__ & ~new_new_n1559__;
  assign new_new_n1561__ = new_new_n1522__ & ~new_new_n1560__;
  assign new_new_n1562__ = ~new_new_n1522__ & new_new_n1560__;
  assign new_new_n1563__ = ~new_new_n1561__ & ~new_new_n1562__;
  assign new_new_n1564__ = new_new_n1496__ & ~new_new_n1563__;
  assign new_new_n1565__ = ~new_new_n1496__ & new_new_n1563__;
  assign new_new_n1566__ = G4091 & ~new_new_n1564__;
  assign new_new_n1567__ = ~new_new_n1565__ & new_new_n1566__;
  assign new_new_n1568__ = new_new_n1489__ & ~new_new_n1567__;
  assign G882 = ~new_new_n1491__ & ~new_new_n1568__;
  assign new_new_n1570__ = G94 & G4092;
  assign new_new_n1571__ = ~new_new_n1393__ & ~new_new_n1570__;
  assign new_new_n1572__ = new_new_n726__ & ~new_new_n1571__;
  assign new_new_n1573__ = G97 & G4092;
  assign new_new_n1574__ = ~new_new_n1568__ & ~new_new_n1573__;
  assign new_new_n1575__ = new_new_n728__ & ~new_new_n1574__;
  assign new_new_n1576__ = ~G14 & ~G4088;
  assign new_new_n1577__ = ~G64 & G4088;
  assign new_new_n1578__ = G4087 & ~new_new_n1576__;
  assign new_new_n1579__ = ~new_new_n1577__ & new_new_n1578__;
  assign new_new_n1580__ = ~new_new_n1572__ & ~new_new_n1579__;
  assign G767 = new_new_n1575__ | ~new_new_n1580__;
  assign new_new_n1582__ = new_new_n769__ & ~new_new_n1571__;
  assign new_new_n1583__ = new_new_n771__ & ~new_new_n1574__;
  assign new_new_n1584__ = ~G14 & ~G4089;
  assign new_new_n1585__ = ~G64 & G4089;
  assign new_new_n1586__ = G4090 & ~new_new_n1584__;
  assign new_new_n1587__ = ~new_new_n1585__ & new_new_n1586__;
  assign new_new_n1588__ = ~new_new_n1582__ & ~new_new_n1587__;
  assign G807 = new_new_n1583__ | ~new_new_n1588__;
  assign new_new_n1590__ = new_new_n926__ & ~new_new_n1571__;
  assign new_new_n1591__ = new_new_n928__ & ~new_new_n1574__;
  assign new_new_n1592__ = ~G176 & ~G1689;
  assign new_new_n1593__ = ~G179 & G1689;
  assign new_new_n1594__ = G1690 & ~new_new_n1592__;
  assign new_new_n1595__ = ~new_new_n1593__ & new_new_n1594__;
  assign new_new_n1596__ = ~new_new_n1590__ & ~new_new_n1595__;
  assign new_new_n1597__ = ~new_new_n1591__ & new_new_n1596__;
  assign G658 = ~G137 | new_new_n1597__;
  assign new_new_n1599__ = new_new_n937__ & ~new_new_n1571__;
  assign new_new_n1600__ = new_new_n939__ & ~new_new_n1574__;
  assign new_new_n1601__ = ~G176 & ~G1691;
  assign new_new_n1602__ = ~G179 & G1691;
  assign new_new_n1603__ = G1694 & ~new_new_n1601__;
  assign new_new_n1604__ = ~new_new_n1602__ & new_new_n1603__;
  assign new_new_n1605__ = ~new_new_n1599__ & ~new_new_n1604__;
  assign new_new_n1606__ = ~new_new_n1600__ & new_new_n1605__;
  assign G690 = ~G137 | new_new_n1606__;
  assign G594 = ~G545;
  assign G599 = ~G348;
  assign G600 = ~G366;
  assign G602 = ~G549;
  assign G611 = ~G338;
  assign G612 = ~G358;
  assign G848 = ~G245;
  assign G849 = ~G552;
  assign G850 = ~G562;
  assign G851 = ~G559;
  assign G593 = ~G299;
  // assign G144 = G141;
  // assign G298 = G293;
  // assign G973 = G3173;
  // assign G603 = G594;
  // assign G604 = G594;
  // assign G926 = G137;
  // assign G923 = G141;
  // assign G921 = G1;
  // assign G892 = G549;
  // assign G887 = G299;
  // assign G606 = G602;
  // assign G993 = G1;
  // assign G978 = G1;
  // assign G949 = G1;
  // assign G939 = G1;
  // assign G889 = G299;
  // assign G717 = G704;
  // assign G626 = G615;
  // assign G632 = G588;
  // assign G621 = G591;
  // assign G629 = G618;
endmodule


