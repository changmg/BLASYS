// Benchmark "ex" written by ABC on Fri Jul  1 14:06:52 2022

module ex ( 
    a, b, c, d, e, f, g, h, i, j, k, l,
    F  );
  input  a, b, c, d, e, f, g, h, i, j, k, l;
  output F;
  assign F = g & c;
endmodule


