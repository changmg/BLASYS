module mult16_19(pi0 , pi1 , pi2 , pi3 , pi4 , po0 , po1 , po2 );
  input pi0 , pi1 , pi2 , pi3 , pi4 ;
  output po0 , po1 , po2 ;
  wire new_n6, new_n7, new_n8, new_n9, new_n10, new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22;
  assign new_n6 = ~pi0 & pi1 ;
  assign new_n7 = pi0 & ~pi1 ;
  assign new_n8 = ~new_n6 & ~new_n7 ;
  assign new_n9 = ~pi2 & pi3 ;
  assign new_n10 = pi2 & ~pi3 ;
  assign new_n11 = ~new_n9 & ~new_n10 ;
  assign new_n12 = new_n8 & new_n11 ;
  assign new_n13 = ~new_n8 & ~new_n11 ;
  assign new_n14 = ~new_n12 & ~new_n13 ;
  assign new_n15 = ~new_n9 & ~new_n12 ;
  assign new_n16 = pi4 & ~new_n15 ;
  assign new_n17 = ~pi4 & new_n15 ;
  assign new_n18 = ~new_n16 & ~new_n17 ;
  assign new_n19 = new_n6 & new_n18 ;
  assign new_n20 = ~new_n6 & ~new_n18 ;
  assign new_n21 = ~new_n19 & ~new_n20 ;
  assign new_n22 = ~new_n16 & ~new_n19 ;
  assign po0 = new_n14 ;
  assign po1 = new_n21 ;
  assign po2 = new_n22 ;
endmodule
