// Benchmark "c1355" written by ABC on Thu Jul 14 21:13:49 2022

module c1355 ( 
    G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat,
    G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat,
    G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat,
    G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat,
    G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat,
    G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat,
    G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat,
    G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat,
    G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat,
    G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_new_n74__, new_new_n75__, new_new_n76__, new_new_n77__,
    new_new_n78__, new_new_n79__, new_new_n80__, new_new_n81__,
    new_new_n82__, new_new_n83__, new_new_n84__, new_new_n85__,
    new_new_n86__, new_new_n87__, new_new_n88__, new_new_n89__,
    new_new_n90__, new_new_n91__, new_new_n92__, new_new_n93__,
    new_new_n94__, new_new_n95__, new_new_n96__, new_new_n97__,
    new_new_n98__, new_new_n99__, new_new_n100__, new_new_n101__,
    new_new_n102__, new_new_n103__, new_new_n104__, new_new_n105__,
    new_new_n106__, new_new_n107__, new_new_n108__, new_new_n109__,
    new_new_n110__, new_new_n111__, new_new_n112__, new_new_n113__,
    new_new_n114__, new_new_n115__, new_new_n116__, new_new_n117__,
    new_new_n118__, new_new_n119__, new_new_n120__, new_new_n121__,
    new_new_n122__, new_new_n123__, new_new_n124__, new_new_n125__,
    new_new_n126__, new_new_n127__, new_new_n128__, new_new_n129__,
    new_new_n130__, new_new_n131__, new_new_n132__, new_new_n133__,
    new_new_n134__, new_new_n135__, new_new_n136__, new_new_n137__,
    new_new_n138__, new_new_n139__, new_new_n140__, new_new_n141__,
    new_new_n142__, new_new_n143__, new_new_n144__, new_new_n145__,
    new_new_n146__, new_new_n147__, new_new_n148__, new_new_n149__,
    new_new_n150__, new_new_n151__, new_new_n152__, new_new_n153__,
    new_new_n154__, new_new_n155__, new_new_n156__, new_new_n157__,
    new_new_n158__, new_new_n159__, new_new_n160__, new_new_n161__,
    new_new_n162__, new_new_n163__, new_new_n164__, new_new_n165__,
    new_new_n166__, new_new_n167__, new_new_n168__, new_new_n169__,
    new_new_n170__, new_new_n171__, new_new_n172__, new_new_n173__,
    new_new_n174__, new_new_n175__, new_new_n176__, new_new_n177__,
    new_new_n178__, new_new_n179__, new_new_n180__, new_new_n181__,
    new_new_n182__, new_new_n183__, new_new_n184__, new_new_n185__,
    new_new_n186__, new_new_n187__, new_new_n188__, new_new_n189__,
    new_new_n190__, new_new_n191__, new_new_n192__, new_new_n193__,
    new_new_n194__, new_new_n195__, new_new_n196__, new_new_n197__,
    new_new_n198__, new_new_n199__, new_new_n200__, new_new_n201__,
    new_new_n202__, new_new_n203__, new_new_n204__, new_new_n205__,
    new_new_n206__, new_new_n207__, new_new_n208__, new_new_n209__,
    new_new_n210__, new_new_n211__, new_new_n212__, new_new_n213__,
    new_new_n214__, new_new_n215__, new_new_n216__, new_new_n217__,
    new_new_n218__, new_new_n219__, new_new_n220__, new_new_n221__,
    new_new_n222__, new_new_n223__, new_new_n224__, new_new_n225__,
    new_new_n226__, new_new_n227__, new_new_n228__, new_new_n229__,
    new_new_n230__, new_new_n231__, new_new_n232__, new_new_n233__,
    new_new_n234__, new_new_n235__, new_new_n236__, new_new_n237__,
    new_new_n238__, new_new_n239__, new_new_n240__, new_new_n241__,
    new_new_n242__, new_new_n243__, new_new_n244__, new_new_n245__,
    new_new_n246__, new_new_n247__, new_new_n248__, new_new_n249__,
    new_new_n250__, new_new_n251__, new_new_n252__, new_new_n253__,
    new_new_n254__, new_new_n255__, new_new_n256__, new_new_n257__,
    new_new_n258__, new_new_n259__, new_new_n260__, new_new_n261__,
    new_new_n262__, new_new_n263__, new_new_n264__, new_new_n265__,
    new_new_n266__, new_new_n267__, new_new_n268__, new_new_n269__,
    new_new_n270__, new_new_n271__, new_new_n272__, new_new_n273__,
    new_new_n274__, new_new_n275__, new_new_n276__, new_new_n277__,
    new_new_n278__, new_new_n279__, new_new_n280__, new_new_n281__,
    new_new_n282__, new_new_n283__, new_new_n284__, new_new_n285__,
    new_new_n286__, new_new_n287__, new_new_n288__, new_new_n289__,
    new_new_n290__, new_new_n291__, new_new_n292__, new_new_n293__,
    new_new_n294__, new_new_n295__, new_new_n296__, new_new_n297__,
    new_new_n298__, new_new_n299__, new_new_n300__, new_new_n301__,
    new_new_n302__, new_new_n303__, new_new_n304__, new_new_n305__,
    new_new_n306__, new_new_n307__, new_new_n308__, new_new_n309__,
    new_new_n310__, new_new_n311__, new_new_n312__, new_new_n313__,
    new_new_n314__, new_new_n315__, new_new_n317__, new_new_n318__,
    new_new_n319__, new_new_n321__, new_new_n322__, new_new_n323__,
    new_new_n325__, new_new_n326__, new_new_n327__, new_new_n329__,
    new_new_n330__, new_new_n331__, new_new_n332__, new_new_n333__,
    new_new_n334__, new_new_n336__, new_new_n337__, new_new_n338__,
    new_new_n340__, new_new_n341__, new_new_n342__, new_new_n344__,
    new_new_n345__, new_new_n346__, new_new_n348__, new_new_n349__,
    new_new_n350__, new_new_n351__, new_new_n352__, new_new_n353__,
    new_new_n355__, new_new_n356__, new_new_n357__, new_new_n359__,
    new_new_n360__, new_new_n361__, new_new_n363__, new_new_n364__,
    new_new_n365__, new_new_n367__, new_new_n368__, new_new_n369__,
    new_new_n370__, new_new_n371__, new_new_n373__, new_new_n374__,
    new_new_n375__, new_new_n377__, new_new_n378__, new_new_n379__,
    new_new_n381__, new_new_n382__, new_new_n383__, new_new_n385__,
    new_new_n386__, new_new_n387__, new_new_n388__, new_new_n389__,
    new_new_n390__, new_new_n391__, new_new_n392__, new_new_n393__,
    new_new_n394__, new_new_n395__, new_new_n396__, new_new_n398__,
    new_new_n399__, new_new_n400__, new_new_n402__, new_new_n403__,
    new_new_n404__, new_new_n406__, new_new_n407__, new_new_n408__,
    new_new_n410__, new_new_n411__, new_new_n412__, new_new_n413__,
    new_new_n414__, new_new_n416__, new_new_n417__, new_new_n418__,
    new_new_n420__, new_new_n421__, new_new_n422__, new_new_n424__,
    new_new_n425__, new_new_n426__, new_new_n428__, new_new_n429__,
    new_new_n430__, new_new_n431__, new_new_n432__, new_new_n434__,
    new_new_n435__, new_new_n436__, new_new_n438__, new_new_n439__,
    new_new_n440__, new_new_n442__, new_new_n443__, new_new_n444__,
    new_new_n446__, new_new_n447__, new_new_n448__, new_new_n449__,
    new_new_n450__, new_new_n452__, new_new_n453__, new_new_n454__,
    new_new_n456__, new_new_n457__, new_new_n458__, new_new_n460__,
    new_new_n461__, new_new_n462__;
  assign new_new_n74__ = G225gat & G233gat;
  assign new_new_n75__ = ~G127gat & ~G134gat;
  assign new_new_n76__ = G127gat & G134gat;
  assign new_new_n77__ = ~new_new_n75__ & ~new_new_n76__;
  assign new_new_n78__ = G113gat & ~G120gat;
  assign new_new_n79__ = ~G113gat & G120gat;
  assign new_new_n80__ = ~new_new_n78__ & ~new_new_n79__;
  assign new_new_n81__ = new_new_n77__ & new_new_n80__;
  assign new_new_n82__ = ~new_new_n77__ & ~new_new_n80__;
  assign new_new_n83__ = ~new_new_n81__ & ~new_new_n82__;
  assign new_new_n84__ = new_new_n74__ & new_new_n83__;
  assign new_new_n85__ = ~new_new_n74__ & ~new_new_n83__;
  assign new_new_n86__ = ~new_new_n84__ & ~new_new_n85__;
  assign new_new_n87__ = ~G57gat & ~G85gat;
  assign new_new_n88__ = G57gat & G85gat;
  assign new_new_n89__ = ~new_new_n87__ & ~new_new_n88__;
  assign new_new_n90__ = G1gat & ~G29gat;
  assign new_new_n91__ = ~G1gat & G29gat;
  assign new_new_n92__ = ~new_new_n90__ & ~new_new_n91__;
  assign new_new_n93__ = new_new_n89__ & new_new_n92__;
  assign new_new_n94__ = ~new_new_n89__ & ~new_new_n92__;
  assign new_new_n95__ = ~new_new_n93__ & ~new_new_n94__;
  assign new_new_n96__ = ~G155gat & ~G162gat;
  assign new_new_n97__ = G155gat & G162gat;
  assign new_new_n98__ = ~new_new_n96__ & ~new_new_n97__;
  assign new_new_n99__ = G141gat & ~G148gat;
  assign new_new_n100__ = ~G141gat & G148gat;
  assign new_new_n101__ = ~new_new_n99__ & ~new_new_n100__;
  assign new_new_n102__ = new_new_n98__ & new_new_n101__;
  assign new_new_n103__ = ~new_new_n98__ & ~new_new_n101__;
  assign new_new_n104__ = ~new_new_n102__ & ~new_new_n103__;
  assign new_new_n105__ = new_new_n95__ & ~new_new_n104__;
  assign new_new_n106__ = ~new_new_n95__ & new_new_n104__;
  assign new_new_n107__ = ~new_new_n105__ & ~new_new_n106__;
  assign new_new_n108__ = new_new_n86__ & new_new_n107__;
  assign new_new_n109__ = ~new_new_n86__ & ~new_new_n107__;
  assign new_new_n110__ = ~new_new_n108__ & ~new_new_n109__;
  assign new_new_n111__ = G229gat & G233gat;
  assign new_new_n112__ = ~G43gat & ~G50gat;
  assign new_new_n113__ = G43gat & G50gat;
  assign new_new_n114__ = ~new_new_n112__ & ~new_new_n113__;
  assign new_new_n115__ = G29gat & ~G36gat;
  assign new_new_n116__ = ~G29gat & G36gat;
  assign new_new_n117__ = ~new_new_n115__ & ~new_new_n116__;
  assign new_new_n118__ = new_new_n114__ & new_new_n117__;
  assign new_new_n119__ = ~new_new_n114__ & ~new_new_n117__;
  assign new_new_n120__ = ~new_new_n118__ & ~new_new_n119__;
  assign new_new_n121__ = new_new_n111__ & new_new_n120__;
  assign new_new_n122__ = ~new_new_n111__ & ~new_new_n120__;
  assign new_new_n123__ = ~new_new_n121__ & ~new_new_n122__;
  assign new_new_n124__ = ~G15gat & ~G22gat;
  assign new_new_n125__ = G15gat & G22gat;
  assign new_new_n126__ = ~new_new_n124__ & ~new_new_n125__;
  assign new_new_n127__ = G1gat & ~G8gat;
  assign new_new_n128__ = ~G1gat & G8gat;
  assign new_new_n129__ = ~new_new_n127__ & ~new_new_n128__;
  assign new_new_n130__ = new_new_n126__ & new_new_n129__;
  assign new_new_n131__ = ~new_new_n126__ & ~new_new_n129__;
  assign new_new_n132__ = ~new_new_n130__ & ~new_new_n131__;
  assign new_new_n133__ = ~G169gat & ~G197gat;
  assign new_new_n134__ = G169gat & G197gat;
  assign new_new_n135__ = ~new_new_n133__ & ~new_new_n134__;
  assign new_new_n136__ = G113gat & ~G141gat;
  assign new_new_n137__ = ~G113gat & G141gat;
  assign new_new_n138__ = ~new_new_n136__ & ~new_new_n137__;
  assign new_new_n139__ = new_new_n135__ & ~new_new_n138__;
  assign new_new_n140__ = ~new_new_n135__ & new_new_n138__;
  assign new_new_n141__ = ~new_new_n139__ & ~new_new_n140__;
  assign new_new_n142__ = new_new_n132__ & ~new_new_n141__;
  assign new_new_n143__ = ~new_new_n132__ & new_new_n141__;
  assign new_new_n144__ = ~new_new_n142__ & ~new_new_n143__;
  assign new_new_n145__ = new_new_n123__ & new_new_n144__;
  assign new_new_n146__ = ~new_new_n123__ & ~new_new_n144__;
  assign new_new_n147__ = ~new_new_n145__ & ~new_new_n146__;
  assign new_new_n148__ = G230gat & G233gat;
  assign new_new_n149__ = ~G99gat & ~G106gat;
  assign new_new_n150__ = G99gat & G106gat;
  assign new_new_n151__ = ~new_new_n149__ & ~new_new_n150__;
  assign new_new_n152__ = G85gat & ~G92gat;
  assign new_new_n153__ = ~G85gat & G92gat;
  assign new_new_n154__ = ~new_new_n152__ & ~new_new_n153__;
  assign new_new_n155__ = new_new_n151__ & new_new_n154__;
  assign new_new_n156__ = ~new_new_n151__ & ~new_new_n154__;
  assign new_new_n157__ = ~new_new_n155__ & ~new_new_n156__;
  assign new_new_n158__ = new_new_n148__ & new_new_n157__;
  assign new_new_n159__ = ~new_new_n148__ & ~new_new_n157__;
  assign new_new_n160__ = ~new_new_n158__ & ~new_new_n159__;
  assign new_new_n161__ = ~G71gat & ~G78gat;
  assign new_new_n162__ = G71gat & G78gat;
  assign new_new_n163__ = ~new_new_n161__ & ~new_new_n162__;
  assign new_new_n164__ = G57gat & ~G64gat;
  assign new_new_n165__ = ~G57gat & G64gat;
  assign new_new_n166__ = ~new_new_n164__ & ~new_new_n165__;
  assign new_new_n167__ = new_new_n163__ & new_new_n166__;
  assign new_new_n168__ = ~new_new_n163__ & ~new_new_n166__;
  assign new_new_n169__ = ~new_new_n167__ & ~new_new_n168__;
  assign new_new_n170__ = ~G176gat & ~G204gat;
  assign new_new_n171__ = G176gat & G204gat;
  assign new_new_n172__ = ~new_new_n170__ & ~new_new_n171__;
  assign new_new_n173__ = G120gat & ~G148gat;
  assign new_new_n174__ = ~G120gat & G148gat;
  assign new_new_n175__ = ~new_new_n173__ & ~new_new_n174__;
  assign new_new_n176__ = new_new_n172__ & ~new_new_n175__;
  assign new_new_n177__ = ~new_new_n172__ & new_new_n175__;
  assign new_new_n178__ = ~new_new_n176__ & ~new_new_n177__;
  assign new_new_n179__ = new_new_n169__ & ~new_new_n178__;
  assign new_new_n180__ = ~new_new_n169__ & new_new_n178__;
  assign new_new_n181__ = ~new_new_n179__ & ~new_new_n180__;
  assign new_new_n182__ = new_new_n160__ & new_new_n181__;
  assign new_new_n183__ = ~new_new_n160__ & ~new_new_n181__;
  assign new_new_n184__ = ~new_new_n182__ & ~new_new_n183__;
  assign new_new_n185__ = ~new_new_n147__ & new_new_n184__;
  assign new_new_n186__ = G232gat & G233gat;
  assign new_new_n187__ = new_new_n120__ & new_new_n186__;
  assign new_new_n188__ = ~new_new_n120__ & ~new_new_n186__;
  assign new_new_n189__ = ~new_new_n187__ & ~new_new_n188__;
  assign new_new_n190__ = ~G190gat & ~G218gat;
  assign new_new_n191__ = G190gat & G218gat;
  assign new_new_n192__ = ~new_new_n190__ & ~new_new_n191__;
  assign new_new_n193__ = G134gat & ~G162gat;
  assign new_new_n194__ = ~G134gat & G162gat;
  assign new_new_n195__ = ~new_new_n193__ & ~new_new_n194__;
  assign new_new_n196__ = new_new_n192__ & ~new_new_n195__;
  assign new_new_n197__ = ~new_new_n192__ & new_new_n195__;
  assign new_new_n198__ = ~new_new_n196__ & ~new_new_n197__;
  assign new_new_n199__ = new_new_n157__ & ~new_new_n198__;
  assign new_new_n200__ = ~new_new_n157__ & new_new_n198__;
  assign new_new_n201__ = ~new_new_n199__ & ~new_new_n200__;
  assign new_new_n202__ = new_new_n189__ & new_new_n201__;
  assign new_new_n203__ = ~new_new_n189__ & ~new_new_n201__;
  assign new_new_n204__ = ~new_new_n202__ & ~new_new_n203__;
  assign new_new_n205__ = G231gat & G233gat;
  assign new_new_n206__ = new_new_n132__ & new_new_n205__;
  assign new_new_n207__ = ~new_new_n132__ & ~new_new_n205__;
  assign new_new_n208__ = ~new_new_n206__ & ~new_new_n207__;
  assign new_new_n209__ = ~G183gat & ~G211gat;
  assign new_new_n210__ = G183gat & G211gat;
  assign new_new_n211__ = ~new_new_n209__ & ~new_new_n210__;
  assign new_new_n212__ = G127gat & ~G155gat;
  assign new_new_n213__ = ~G127gat & G155gat;
  assign new_new_n214__ = ~new_new_n212__ & ~new_new_n213__;
  assign new_new_n215__ = new_new_n211__ & ~new_new_n214__;
  assign new_new_n216__ = ~new_new_n211__ & new_new_n214__;
  assign new_new_n217__ = ~new_new_n215__ & ~new_new_n216__;
  assign new_new_n218__ = new_new_n169__ & ~new_new_n217__;
  assign new_new_n219__ = ~new_new_n169__ & new_new_n217__;
  assign new_new_n220__ = ~new_new_n218__ & ~new_new_n219__;
  assign new_new_n221__ = new_new_n208__ & new_new_n220__;
  assign new_new_n222__ = ~new_new_n208__ & ~new_new_n220__;
  assign new_new_n223__ = ~new_new_n221__ & ~new_new_n222__;
  assign new_new_n224__ = new_new_n204__ & ~new_new_n223__;
  assign new_new_n225__ = G226gat & G233gat;
  assign new_new_n226__ = ~G211gat & ~G218gat;
  assign new_new_n227__ = G211gat & G218gat;
  assign new_new_n228__ = ~new_new_n226__ & ~new_new_n227__;
  assign new_new_n229__ = G197gat & ~G204gat;
  assign new_new_n230__ = ~G197gat & G204gat;
  assign new_new_n231__ = ~new_new_n229__ & ~new_new_n230__;
  assign new_new_n232__ = new_new_n228__ & new_new_n231__;
  assign new_new_n233__ = ~new_new_n228__ & ~new_new_n231__;
  assign new_new_n234__ = ~new_new_n232__ & ~new_new_n233__;
  assign new_new_n235__ = new_new_n225__ & new_new_n234__;
  assign new_new_n236__ = ~new_new_n225__ & ~new_new_n234__;
  assign new_new_n237__ = ~new_new_n235__ & ~new_new_n236__;
  assign new_new_n238__ = ~G183gat & ~G190gat;
  assign new_new_n239__ = G183gat & G190gat;
  assign new_new_n240__ = ~new_new_n238__ & ~new_new_n239__;
  assign new_new_n241__ = G169gat & ~G176gat;
  assign new_new_n242__ = ~G169gat & G176gat;
  assign new_new_n243__ = ~new_new_n241__ & ~new_new_n242__;
  assign new_new_n244__ = new_new_n240__ & new_new_n243__;
  assign new_new_n245__ = ~new_new_n240__ & ~new_new_n243__;
  assign new_new_n246__ = ~new_new_n244__ & ~new_new_n245__;
  assign new_new_n247__ = ~G64gat & ~G92gat;
  assign new_new_n248__ = G64gat & G92gat;
  assign new_new_n249__ = ~new_new_n247__ & ~new_new_n248__;
  assign new_new_n250__ = G8gat & ~G36gat;
  assign new_new_n251__ = ~G8gat & G36gat;
  assign new_new_n252__ = ~new_new_n250__ & ~new_new_n251__;
  assign new_new_n253__ = new_new_n249__ & ~new_new_n252__;
  assign new_new_n254__ = ~new_new_n249__ & new_new_n252__;
  assign new_new_n255__ = ~new_new_n253__ & ~new_new_n254__;
  assign new_new_n256__ = new_new_n246__ & ~new_new_n255__;
  assign new_new_n257__ = ~new_new_n246__ & new_new_n255__;
  assign new_new_n258__ = ~new_new_n256__ & ~new_new_n257__;
  assign new_new_n259__ = new_new_n237__ & new_new_n258__;
  assign new_new_n260__ = ~new_new_n237__ & ~new_new_n258__;
  assign new_new_n261__ = ~new_new_n259__ & ~new_new_n260__;
  assign new_new_n262__ = ~new_new_n110__ & ~new_new_n261__;
  assign new_new_n263__ = new_new_n110__ & new_new_n261__;
  assign new_new_n264__ = ~new_new_n262__ & ~new_new_n263__;
  assign new_new_n265__ = G227gat & G233gat;
  assign new_new_n266__ = new_new_n83__ & new_new_n265__;
  assign new_new_n267__ = ~new_new_n83__ & ~new_new_n265__;
  assign new_new_n268__ = ~new_new_n266__ & ~new_new_n267__;
  assign new_new_n269__ = ~G71gat & ~G99gat;
  assign new_new_n270__ = G71gat & G99gat;
  assign new_new_n271__ = ~new_new_n269__ & ~new_new_n270__;
  assign new_new_n272__ = G15gat & ~G43gat;
  assign new_new_n273__ = ~G15gat & G43gat;
  assign new_new_n274__ = ~new_new_n272__ & ~new_new_n273__;
  assign new_new_n275__ = new_new_n271__ & ~new_new_n274__;
  assign new_new_n276__ = ~new_new_n271__ & new_new_n274__;
  assign new_new_n277__ = ~new_new_n275__ & ~new_new_n276__;
  assign new_new_n278__ = new_new_n246__ & ~new_new_n277__;
  assign new_new_n279__ = ~new_new_n246__ & new_new_n277__;
  assign new_new_n280__ = ~new_new_n278__ & ~new_new_n279__;
  assign new_new_n281__ = new_new_n268__ & new_new_n280__;
  assign new_new_n282__ = ~new_new_n268__ & ~new_new_n280__;
  assign new_new_n283__ = ~new_new_n281__ & ~new_new_n282__;
  assign new_new_n284__ = G228gat & G233gat;
  assign new_new_n285__ = new_new_n104__ & new_new_n284__;
  assign new_new_n286__ = ~new_new_n104__ & ~new_new_n284__;
  assign new_new_n287__ = ~new_new_n285__ & ~new_new_n286__;
  assign new_new_n288__ = ~G78gat & ~G106gat;
  assign new_new_n289__ = G78gat & G106gat;
  assign new_new_n290__ = ~new_new_n288__ & ~new_new_n289__;
  assign new_new_n291__ = G22gat & ~G50gat;
  assign new_new_n292__ = ~G22gat & G50gat;
  assign new_new_n293__ = ~new_new_n291__ & ~new_new_n292__;
  assign new_new_n294__ = new_new_n290__ & ~new_new_n293__;
  assign new_new_n295__ = ~new_new_n290__ & new_new_n293__;
  assign new_new_n296__ = ~new_new_n294__ & ~new_new_n295__;
  assign new_new_n297__ = new_new_n234__ & ~new_new_n296__;
  assign new_new_n298__ = ~new_new_n234__ & new_new_n296__;
  assign new_new_n299__ = ~new_new_n297__ & ~new_new_n298__;
  assign new_new_n300__ = new_new_n287__ & new_new_n299__;
  assign new_new_n301__ = ~new_new_n287__ & ~new_new_n299__;
  assign new_new_n302__ = ~new_new_n300__ & ~new_new_n301__;
  assign new_new_n303__ = new_new_n283__ & new_new_n302__;
  assign new_new_n304__ = ~new_new_n264__ & new_new_n303__;
  assign new_new_n305__ = new_new_n283__ & ~new_new_n302__;
  assign new_new_n306__ = ~new_new_n283__ & new_new_n302__;
  assign new_new_n307__ = ~new_new_n305__ & ~new_new_n306__;
  assign new_new_n308__ = ~new_new_n110__ & new_new_n261__;
  assign new_new_n309__ = ~new_new_n307__ & new_new_n308__;
  assign new_new_n310__ = ~new_new_n304__ & ~new_new_n309__;
  assign new_new_n311__ = new_new_n185__ & new_new_n224__;
  assign new_new_n312__ = ~new_new_n310__ & new_new_n311__;
  assign new_new_n313__ = new_new_n110__ & new_new_n312__;
  assign new_new_n314__ = G1gat & ~new_new_n313__;
  assign new_new_n315__ = ~G1gat & new_new_n313__;
  assign G1324gat = new_new_n314__ | new_new_n315__;
  assign new_new_n317__ = ~new_new_n261__ & new_new_n312__;
  assign new_new_n318__ = G8gat & ~new_new_n317__;
  assign new_new_n319__ = ~G8gat & new_new_n317__;
  assign G1325gat = new_new_n318__ | new_new_n319__;
  assign new_new_n321__ = ~new_new_n283__ & new_new_n312__;
  assign new_new_n322__ = G15gat & ~new_new_n321__;
  assign new_new_n323__ = ~G15gat & new_new_n321__;
  assign G1326gat = new_new_n322__ | new_new_n323__;
  assign new_new_n325__ = ~new_new_n302__ & new_new_n312__;
  assign new_new_n326__ = G22gat & ~new_new_n325__;
  assign new_new_n327__ = ~G22gat & new_new_n325__;
  assign G1327gat = new_new_n326__ | new_new_n327__;
  assign new_new_n329__ = ~new_new_n204__ & new_new_n223__;
  assign new_new_n330__ = new_new_n185__ & new_new_n329__;
  assign new_new_n331__ = ~new_new_n310__ & new_new_n330__;
  assign new_new_n332__ = new_new_n110__ & new_new_n331__;
  assign new_new_n333__ = G29gat & ~new_new_n332__;
  assign new_new_n334__ = ~G29gat & new_new_n332__;
  assign G1328gat = new_new_n333__ | new_new_n334__;
  assign new_new_n336__ = ~new_new_n261__ & new_new_n331__;
  assign new_new_n337__ = G36gat & ~new_new_n336__;
  assign new_new_n338__ = ~G36gat & new_new_n336__;
  assign G1329gat = new_new_n337__ | new_new_n338__;
  assign new_new_n340__ = ~new_new_n283__ & new_new_n331__;
  assign new_new_n341__ = G43gat & ~new_new_n340__;
  assign new_new_n342__ = ~G43gat & new_new_n340__;
  assign G1330gat = new_new_n341__ | new_new_n342__;
  assign new_new_n344__ = ~new_new_n302__ & new_new_n331__;
  assign new_new_n345__ = G50gat & ~new_new_n344__;
  assign new_new_n346__ = ~G50gat & new_new_n344__;
  assign G1331gat = new_new_n345__ | new_new_n346__;
  assign new_new_n348__ = new_new_n147__ & ~new_new_n184__;
  assign new_new_n349__ = new_new_n224__ & new_new_n348__;
  assign new_new_n350__ = ~new_new_n310__ & new_new_n349__;
  assign new_new_n351__ = new_new_n110__ & new_new_n350__;
  assign new_new_n352__ = G57gat & ~new_new_n351__;
  assign new_new_n353__ = ~G57gat & new_new_n351__;
  assign G1332gat = new_new_n352__ | new_new_n353__;
  assign new_new_n355__ = ~new_new_n261__ & new_new_n350__;
  assign new_new_n356__ = G64gat & ~new_new_n355__;
  assign new_new_n357__ = ~G64gat & new_new_n355__;
  assign G1333gat = new_new_n356__ | new_new_n357__;
  assign new_new_n359__ = ~new_new_n283__ & new_new_n350__;
  assign new_new_n360__ = G71gat & ~new_new_n359__;
  assign new_new_n361__ = ~G71gat & new_new_n359__;
  assign G1334gat = new_new_n360__ | new_new_n361__;
  assign new_new_n363__ = ~new_new_n302__ & new_new_n350__;
  assign new_new_n364__ = G78gat & ~new_new_n363__;
  assign new_new_n365__ = ~G78gat & new_new_n363__;
  assign G1335gat = new_new_n364__ | new_new_n365__;
  assign new_new_n367__ = new_new_n329__ & new_new_n348__;
  assign new_new_n368__ = ~new_new_n310__ & new_new_n367__;
  assign new_new_n369__ = new_new_n110__ & new_new_n368__;
  assign new_new_n370__ = G85gat & ~new_new_n369__;
  assign new_new_n371__ = ~G85gat & new_new_n369__;
  assign G1336gat = new_new_n370__ | new_new_n371__;
  assign new_new_n373__ = ~new_new_n261__ & new_new_n368__;
  assign new_new_n374__ = G92gat & ~new_new_n373__;
  assign new_new_n375__ = ~G92gat & new_new_n373__;
  assign G1337gat = new_new_n374__ | new_new_n375__;
  assign new_new_n377__ = ~new_new_n283__ & new_new_n368__;
  assign new_new_n378__ = G99gat & ~new_new_n377__;
  assign new_new_n379__ = ~G99gat & new_new_n377__;
  assign G1338gat = new_new_n378__ | new_new_n379__;
  assign new_new_n381__ = ~new_new_n302__ & new_new_n368__;
  assign new_new_n382__ = G106gat & ~new_new_n381__;
  assign new_new_n383__ = ~G106gat & new_new_n381__;
  assign G1339gat = new_new_n382__ | new_new_n383__;
  assign new_new_n385__ = ~new_new_n185__ & ~new_new_n348__;
  assign new_new_n386__ = new_new_n204__ & new_new_n223__;
  assign new_new_n387__ = ~new_new_n385__ & new_new_n386__;
  assign new_new_n388__ = ~new_new_n224__ & ~new_new_n329__;
  assign new_new_n389__ = new_new_n147__ & new_new_n184__;
  assign new_new_n390__ = ~new_new_n388__ & new_new_n389__;
  assign new_new_n391__ = ~new_new_n387__ & ~new_new_n390__;
  assign new_new_n392__ = new_new_n263__ & new_new_n306__;
  assign new_new_n393__ = ~new_new_n391__ & new_new_n392__;
  assign new_new_n394__ = ~new_new_n147__ & new_new_n393__;
  assign new_new_n395__ = G113gat & ~new_new_n394__;
  assign new_new_n396__ = ~G113gat & new_new_n394__;
  assign G1340gat = new_new_n395__ | new_new_n396__;
  assign new_new_n398__ = ~new_new_n184__ & new_new_n393__;
  assign new_new_n399__ = G120gat & ~new_new_n398__;
  assign new_new_n400__ = ~G120gat & new_new_n398__;
  assign G1341gat = new_new_n399__ | new_new_n400__;
  assign new_new_n402__ = ~new_new_n223__ & new_new_n393__;
  assign new_new_n403__ = G127gat & ~new_new_n402__;
  assign new_new_n404__ = ~G127gat & new_new_n402__;
  assign G1342gat = new_new_n403__ | new_new_n404__;
  assign new_new_n406__ = ~new_new_n204__ & new_new_n393__;
  assign new_new_n407__ = G134gat & ~new_new_n406__;
  assign new_new_n408__ = ~G134gat & new_new_n406__;
  assign G1343gat = new_new_n407__ | new_new_n408__;
  assign new_new_n410__ = new_new_n263__ & new_new_n305__;
  assign new_new_n411__ = ~new_new_n391__ & new_new_n410__;
  assign new_new_n412__ = ~new_new_n147__ & new_new_n411__;
  assign new_new_n413__ = G141gat & ~new_new_n412__;
  assign new_new_n414__ = ~G141gat & new_new_n412__;
  assign G1344gat = new_new_n413__ | new_new_n414__;
  assign new_new_n416__ = ~new_new_n184__ & new_new_n411__;
  assign new_new_n417__ = G148gat & ~new_new_n416__;
  assign new_new_n418__ = ~G148gat & new_new_n416__;
  assign G1345gat = new_new_n417__ | new_new_n418__;
  assign new_new_n420__ = ~new_new_n223__ & new_new_n411__;
  assign new_new_n421__ = G155gat & ~new_new_n420__;
  assign new_new_n422__ = ~G155gat & new_new_n420__;
  assign G1346gat = new_new_n421__ | new_new_n422__;
  assign new_new_n424__ = ~new_new_n204__ & new_new_n411__;
  assign new_new_n425__ = G162gat & ~new_new_n424__;
  assign new_new_n426__ = ~G162gat & new_new_n424__;
  assign G1347gat = new_new_n425__ | new_new_n426__;
  assign new_new_n428__ = new_new_n262__ & new_new_n306__;
  assign new_new_n429__ = ~new_new_n391__ & new_new_n428__;
  assign new_new_n430__ = ~new_new_n147__ & new_new_n429__;
  assign new_new_n431__ = G169gat & ~new_new_n430__;
  assign new_new_n432__ = ~G169gat & new_new_n430__;
  assign G1348gat = new_new_n431__ | new_new_n432__;
  assign new_new_n434__ = ~new_new_n184__ & new_new_n429__;
  assign new_new_n435__ = G176gat & ~new_new_n434__;
  assign new_new_n436__ = ~G176gat & new_new_n434__;
  assign G1349gat = new_new_n435__ | new_new_n436__;
  assign new_new_n438__ = ~new_new_n223__ & new_new_n429__;
  assign new_new_n439__ = G183gat & ~new_new_n438__;
  assign new_new_n440__ = ~G183gat & new_new_n438__;
  assign G1350gat = new_new_n439__ | new_new_n440__;
  assign new_new_n442__ = ~new_new_n204__ & new_new_n429__;
  assign new_new_n443__ = G190gat & ~new_new_n442__;
  assign new_new_n444__ = ~G190gat & new_new_n442__;
  assign G1351gat = new_new_n443__ | new_new_n444__;
  assign new_new_n446__ = new_new_n262__ & new_new_n305__;
  assign new_new_n447__ = ~new_new_n391__ & new_new_n446__;
  assign new_new_n448__ = ~new_new_n147__ & new_new_n447__;
  assign new_new_n449__ = G197gat & ~new_new_n448__;
  assign new_new_n450__ = ~G197gat & new_new_n448__;
  assign G1352gat = new_new_n449__ | new_new_n450__;
  assign new_new_n452__ = ~new_new_n184__ & new_new_n447__;
  assign new_new_n453__ = G204gat & ~new_new_n452__;
  assign new_new_n454__ = ~G204gat & new_new_n452__;
  assign G1353gat = new_new_n453__ | new_new_n454__;
  assign new_new_n456__ = ~new_new_n223__ & new_new_n447__;
  assign new_new_n457__ = G211gat & ~new_new_n456__;
  assign new_new_n458__ = ~G211gat & new_new_n456__;
  assign G1354gat = new_new_n457__ | new_new_n458__;
  assign new_new_n460__ = ~new_new_n204__ & new_new_n447__;
  assign new_new_n461__ = G218gat & ~new_new_n460__;
  assign new_new_n462__ = ~G218gat & new_new_n460__;
  assign G1355gat = new_new_n461__ | new_new_n462__;
endmodule


