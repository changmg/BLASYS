// Benchmark "ex" written by ABC on Thu Jul 14 00:21:06 2022

module ex ( 
    a, b, c, d, e, f,
    F  );
  input  a, b, c, d, e, f;
  output F;
  assign F = f;
endmodule


