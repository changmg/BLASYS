// Benchmark "c6288" written by ABC on Thu Jul 14 21:14:36 2022

module c6288 ( 
    G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat,
    G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat,
    G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat,
    G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat,
    G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat  );
  input  G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat,
    G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat,
    G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat,
    G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat;
  output G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat;
  wire new_new_n66__, new_new_n67__, new_new_n68__, new_new_n69__,
    new_new_n70__, new_new_n72__, new_new_n73__, new_new_n74__,
    new_new_n75__, new_new_n76__, new_new_n77__, new_new_n78__,
    new_new_n79__, new_new_n80__, new_new_n81__, new_new_n82__,
    new_new_n84__, new_new_n85__, new_new_n86__, new_new_n87__,
    new_new_n88__, new_new_n89__, new_new_n90__, new_new_n91__,
    new_new_n92__, new_new_n93__, new_new_n94__, new_new_n95__,
    new_new_n96__, new_new_n97__, new_new_n98__, new_new_n99__,
    new_new_n100__, new_new_n101__, new_new_n102__, new_new_n104__,
    new_new_n105__, new_new_n106__, new_new_n107__, new_new_n108__,
    new_new_n109__, new_new_n110__, new_new_n111__, new_new_n112__,
    new_new_n113__, new_new_n114__, new_new_n115__, new_new_n116__,
    new_new_n117__, new_new_n118__, new_new_n119__, new_new_n120__,
    new_new_n121__, new_new_n122__, new_new_n123__, new_new_n124__,
    new_new_n125__, new_new_n126__, new_new_n127__, new_new_n128__,
    new_new_n129__, new_new_n130__, new_new_n132__, new_new_n133__,
    new_new_n134__, new_new_n135__, new_new_n136__, new_new_n137__,
    new_new_n138__, new_new_n139__, new_new_n140__, new_new_n141__,
    new_new_n142__, new_new_n143__, new_new_n144__, new_new_n145__,
    new_new_n146__, new_new_n147__, new_new_n148__, new_new_n149__,
    new_new_n150__, new_new_n151__, new_new_n152__, new_new_n153__,
    new_new_n154__, new_new_n155__, new_new_n156__, new_new_n157__,
    new_new_n158__, new_new_n159__, new_new_n160__, new_new_n161__,
    new_new_n162__, new_new_n163__, new_new_n164__, new_new_n165__,
    new_new_n166__, new_new_n168__, new_new_n169__, new_new_n170__,
    new_new_n171__, new_new_n172__, new_new_n173__, new_new_n174__,
    new_new_n175__, new_new_n176__, new_new_n177__, new_new_n178__,
    new_new_n179__, new_new_n180__, new_new_n181__, new_new_n182__,
    new_new_n183__, new_new_n184__, new_new_n185__, new_new_n186__,
    new_new_n187__, new_new_n188__, new_new_n189__, new_new_n190__,
    new_new_n191__, new_new_n192__, new_new_n193__, new_new_n194__,
    new_new_n195__, new_new_n196__, new_new_n197__, new_new_n198__,
    new_new_n199__, new_new_n200__, new_new_n201__, new_new_n202__,
    new_new_n203__, new_new_n204__, new_new_n205__, new_new_n206__,
    new_new_n207__, new_new_n208__, new_new_n209__, new_new_n210__,
    new_new_n212__, new_new_n213__, new_new_n214__, new_new_n215__,
    new_new_n216__, new_new_n217__, new_new_n218__, new_new_n219__,
    new_new_n220__, new_new_n221__, new_new_n222__, new_new_n223__,
    new_new_n224__, new_new_n225__, new_new_n226__, new_new_n227__,
    new_new_n228__, new_new_n229__, new_new_n230__, new_new_n231__,
    new_new_n232__, new_new_n233__, new_new_n234__, new_new_n235__,
    new_new_n236__, new_new_n237__, new_new_n238__, new_new_n239__,
    new_new_n240__, new_new_n241__, new_new_n242__, new_new_n243__,
    new_new_n244__, new_new_n245__, new_new_n246__, new_new_n247__,
    new_new_n248__, new_new_n249__, new_new_n250__, new_new_n251__,
    new_new_n252__, new_new_n253__, new_new_n254__, new_new_n255__,
    new_new_n256__, new_new_n257__, new_new_n258__, new_new_n259__,
    new_new_n260__, new_new_n261__, new_new_n262__, new_new_n264__,
    new_new_n265__, new_new_n266__, new_new_n267__, new_new_n268__,
    new_new_n269__, new_new_n270__, new_new_n271__, new_new_n272__,
    new_new_n273__, new_new_n274__, new_new_n275__, new_new_n276__,
    new_new_n277__, new_new_n278__, new_new_n279__, new_new_n280__,
    new_new_n281__, new_new_n282__, new_new_n283__, new_new_n284__,
    new_new_n285__, new_new_n286__, new_new_n287__, new_new_n288__,
    new_new_n289__, new_new_n290__, new_new_n291__, new_new_n292__,
    new_new_n293__, new_new_n294__, new_new_n295__, new_new_n296__,
    new_new_n297__, new_new_n298__, new_new_n299__, new_new_n300__,
    new_new_n301__, new_new_n302__, new_new_n303__, new_new_n304__,
    new_new_n305__, new_new_n306__, new_new_n307__, new_new_n308__,
    new_new_n309__, new_new_n310__, new_new_n311__, new_new_n312__,
    new_new_n313__, new_new_n314__, new_new_n315__, new_new_n316__,
    new_new_n317__, new_new_n318__, new_new_n319__, new_new_n320__,
    new_new_n321__, new_new_n322__, new_new_n324__, new_new_n325__,
    new_new_n326__, new_new_n327__, new_new_n328__, new_new_n329__,
    new_new_n330__, new_new_n331__, new_new_n332__, new_new_n333__,
    new_new_n334__, new_new_n335__, new_new_n336__, new_new_n337__,
    new_new_n338__, new_new_n339__, new_new_n340__, new_new_n341__,
    new_new_n342__, new_new_n343__, new_new_n344__, new_new_n345__,
    new_new_n346__, new_new_n347__, new_new_n348__, new_new_n349__,
    new_new_n350__, new_new_n351__, new_new_n352__, new_new_n353__,
    new_new_n354__, new_new_n355__, new_new_n356__, new_new_n357__,
    new_new_n358__, new_new_n359__, new_new_n360__, new_new_n361__,
    new_new_n362__, new_new_n363__, new_new_n364__, new_new_n365__,
    new_new_n366__, new_new_n367__, new_new_n368__, new_new_n369__,
    new_new_n370__, new_new_n371__, new_new_n372__, new_new_n373__,
    new_new_n374__, new_new_n375__, new_new_n376__, new_new_n377__,
    new_new_n378__, new_new_n379__, new_new_n380__, new_new_n381__,
    new_new_n382__, new_new_n383__, new_new_n384__, new_new_n385__,
    new_new_n386__, new_new_n387__, new_new_n388__, new_new_n389__,
    new_new_n390__, new_new_n392__, new_new_n393__, new_new_n394__,
    new_new_n395__, new_new_n396__, new_new_n397__, new_new_n398__,
    new_new_n399__, new_new_n400__, new_new_n401__, new_new_n402__,
    new_new_n403__, new_new_n404__, new_new_n405__, new_new_n406__,
    new_new_n407__, new_new_n408__, new_new_n409__, new_new_n410__,
    new_new_n411__, new_new_n412__, new_new_n413__, new_new_n414__,
    new_new_n415__, new_new_n416__, new_new_n417__, new_new_n418__,
    new_new_n419__, new_new_n420__, new_new_n421__, new_new_n422__,
    new_new_n423__, new_new_n424__, new_new_n425__, new_new_n426__,
    new_new_n427__, new_new_n428__, new_new_n429__, new_new_n430__,
    new_new_n431__, new_new_n432__, new_new_n433__, new_new_n434__,
    new_new_n435__, new_new_n436__, new_new_n437__, new_new_n438__,
    new_new_n439__, new_new_n440__, new_new_n441__, new_new_n442__,
    new_new_n443__, new_new_n444__, new_new_n445__, new_new_n446__,
    new_new_n447__, new_new_n448__, new_new_n449__, new_new_n450__,
    new_new_n451__, new_new_n452__, new_new_n453__, new_new_n454__,
    new_new_n455__, new_new_n456__, new_new_n457__, new_new_n458__,
    new_new_n459__, new_new_n460__, new_new_n461__, new_new_n462__,
    new_new_n463__, new_new_n464__, new_new_n465__, new_new_n466__,
    new_new_n468__, new_new_n469__, new_new_n470__, new_new_n471__,
    new_new_n472__, new_new_n473__, new_new_n474__, new_new_n475__,
    new_new_n476__, new_new_n477__, new_new_n478__, new_new_n479__,
    new_new_n480__, new_new_n481__, new_new_n482__, new_new_n483__,
    new_new_n484__, new_new_n485__, new_new_n486__, new_new_n487__,
    new_new_n488__, new_new_n489__, new_new_n490__, new_new_n491__,
    new_new_n492__, new_new_n493__, new_new_n494__, new_new_n495__,
    new_new_n496__, new_new_n497__, new_new_n498__, new_new_n499__,
    new_new_n500__, new_new_n501__, new_new_n502__, new_new_n503__,
    new_new_n504__, new_new_n505__, new_new_n506__, new_new_n507__,
    new_new_n508__, new_new_n509__, new_new_n510__, new_new_n511__,
    new_new_n512__, new_new_n513__, new_new_n514__, new_new_n515__,
    new_new_n516__, new_new_n517__, new_new_n518__, new_new_n519__,
    new_new_n520__, new_new_n521__, new_new_n522__, new_new_n523__,
    new_new_n524__, new_new_n525__, new_new_n526__, new_new_n527__,
    new_new_n528__, new_new_n529__, new_new_n530__, new_new_n531__,
    new_new_n532__, new_new_n533__, new_new_n534__, new_new_n535__,
    new_new_n536__, new_new_n537__, new_new_n538__, new_new_n539__,
    new_new_n540__, new_new_n541__, new_new_n542__, new_new_n543__,
    new_new_n544__, new_new_n545__, new_new_n546__, new_new_n547__,
    new_new_n548__, new_new_n549__, new_new_n550__, new_new_n552__,
    new_new_n553__, new_new_n554__, new_new_n555__, new_new_n556__,
    new_new_n557__, new_new_n558__, new_new_n559__, new_new_n560__,
    new_new_n561__, new_new_n562__, new_new_n563__, new_new_n564__,
    new_new_n565__, new_new_n566__, new_new_n567__, new_new_n568__,
    new_new_n569__, new_new_n570__, new_new_n571__, new_new_n572__,
    new_new_n573__, new_new_n574__, new_new_n575__, new_new_n576__,
    new_new_n577__, new_new_n578__, new_new_n579__, new_new_n580__,
    new_new_n581__, new_new_n582__, new_new_n583__, new_new_n584__,
    new_new_n585__, new_new_n586__, new_new_n587__, new_new_n588__,
    new_new_n589__, new_new_n590__, new_new_n591__, new_new_n592__,
    new_new_n593__, new_new_n594__, new_new_n595__, new_new_n596__,
    new_new_n597__, new_new_n598__, new_new_n599__, new_new_n600__,
    new_new_n601__, new_new_n602__, new_new_n603__, new_new_n604__,
    new_new_n605__, new_new_n606__, new_new_n607__, new_new_n608__,
    new_new_n609__, new_new_n610__, new_new_n611__, new_new_n612__,
    new_new_n613__, new_new_n614__, new_new_n615__, new_new_n616__,
    new_new_n617__, new_new_n618__, new_new_n619__, new_new_n620__,
    new_new_n621__, new_new_n622__, new_new_n623__, new_new_n624__,
    new_new_n625__, new_new_n626__, new_new_n627__, new_new_n628__,
    new_new_n629__, new_new_n630__, new_new_n631__, new_new_n632__,
    new_new_n633__, new_new_n634__, new_new_n635__, new_new_n636__,
    new_new_n637__, new_new_n638__, new_new_n639__, new_new_n640__,
    new_new_n641__, new_new_n642__, new_new_n644__, new_new_n645__,
    new_new_n646__, new_new_n647__, new_new_n648__, new_new_n649__,
    new_new_n650__, new_new_n651__, new_new_n652__, new_new_n653__,
    new_new_n654__, new_new_n655__, new_new_n656__, new_new_n657__,
    new_new_n658__, new_new_n659__, new_new_n660__, new_new_n661__,
    new_new_n662__, new_new_n663__, new_new_n664__, new_new_n665__,
    new_new_n666__, new_new_n667__, new_new_n668__, new_new_n669__,
    new_new_n670__, new_new_n671__, new_new_n672__, new_new_n673__,
    new_new_n674__, new_new_n675__, new_new_n676__, new_new_n677__,
    new_new_n678__, new_new_n679__, new_new_n680__, new_new_n681__,
    new_new_n682__, new_new_n683__, new_new_n684__, new_new_n685__,
    new_new_n686__, new_new_n687__, new_new_n688__, new_new_n689__,
    new_new_n690__, new_new_n691__, new_new_n692__, new_new_n693__,
    new_new_n694__, new_new_n695__, new_new_n696__, new_new_n697__,
    new_new_n698__, new_new_n699__, new_new_n700__, new_new_n701__,
    new_new_n702__, new_new_n703__, new_new_n704__, new_new_n705__,
    new_new_n706__, new_new_n707__, new_new_n708__, new_new_n709__,
    new_new_n710__, new_new_n711__, new_new_n712__, new_new_n713__,
    new_new_n714__, new_new_n715__, new_new_n716__, new_new_n717__,
    new_new_n718__, new_new_n719__, new_new_n720__, new_new_n721__,
    new_new_n722__, new_new_n723__, new_new_n724__, new_new_n725__,
    new_new_n726__, new_new_n727__, new_new_n728__, new_new_n729__,
    new_new_n730__, new_new_n731__, new_new_n732__, new_new_n733__,
    new_new_n734__, new_new_n735__, new_new_n736__, new_new_n737__,
    new_new_n738__, new_new_n739__, new_new_n740__, new_new_n741__,
    new_new_n742__, new_new_n744__, new_new_n745__, new_new_n746__,
    new_new_n747__, new_new_n748__, new_new_n749__, new_new_n750__,
    new_new_n751__, new_new_n752__, new_new_n753__, new_new_n754__,
    new_new_n755__, new_new_n756__, new_new_n757__, new_new_n758__,
    new_new_n759__, new_new_n760__, new_new_n761__, new_new_n762__,
    new_new_n763__, new_new_n764__, new_new_n765__, new_new_n766__,
    new_new_n767__, new_new_n768__, new_new_n769__, new_new_n770__,
    new_new_n771__, new_new_n772__, new_new_n773__, new_new_n774__,
    new_new_n775__, new_new_n776__, new_new_n777__, new_new_n778__,
    new_new_n779__, new_new_n780__, new_new_n781__, new_new_n782__,
    new_new_n783__, new_new_n784__, new_new_n785__, new_new_n786__,
    new_new_n787__, new_new_n788__, new_new_n789__, new_new_n790__,
    new_new_n791__, new_new_n792__, new_new_n793__, new_new_n794__,
    new_new_n795__, new_new_n796__, new_new_n797__, new_new_n798__,
    new_new_n799__, new_new_n800__, new_new_n801__, new_new_n802__,
    new_new_n803__, new_new_n804__, new_new_n805__, new_new_n806__,
    new_new_n807__, new_new_n808__, new_new_n809__, new_new_n810__,
    new_new_n811__, new_new_n812__, new_new_n813__, new_new_n814__,
    new_new_n815__, new_new_n816__, new_new_n817__, new_new_n818__,
    new_new_n819__, new_new_n820__, new_new_n821__, new_new_n822__,
    new_new_n823__, new_new_n824__, new_new_n825__, new_new_n826__,
    new_new_n827__, new_new_n828__, new_new_n829__, new_new_n830__,
    new_new_n831__, new_new_n832__, new_new_n833__, new_new_n834__,
    new_new_n835__, new_new_n836__, new_new_n837__, new_new_n838__,
    new_new_n839__, new_new_n840__, new_new_n841__, new_new_n842__,
    new_new_n843__, new_new_n844__, new_new_n845__, new_new_n846__,
    new_new_n847__, new_new_n848__, new_new_n849__, new_new_n850__,
    new_new_n852__, new_new_n853__, new_new_n854__, new_new_n855__,
    new_new_n856__, new_new_n857__, new_new_n858__, new_new_n859__,
    new_new_n860__, new_new_n861__, new_new_n862__, new_new_n863__,
    new_new_n864__, new_new_n865__, new_new_n866__, new_new_n867__,
    new_new_n868__, new_new_n869__, new_new_n870__, new_new_n871__,
    new_new_n872__, new_new_n873__, new_new_n874__, new_new_n875__,
    new_new_n876__, new_new_n877__, new_new_n878__, new_new_n879__,
    new_new_n880__, new_new_n881__, new_new_n882__, new_new_n883__,
    new_new_n884__, new_new_n885__, new_new_n886__, new_new_n887__,
    new_new_n888__, new_new_n889__, new_new_n890__, new_new_n891__,
    new_new_n892__, new_new_n893__, new_new_n894__, new_new_n895__,
    new_new_n896__, new_new_n897__, new_new_n898__, new_new_n899__,
    new_new_n900__, new_new_n901__, new_new_n902__, new_new_n903__,
    new_new_n904__, new_new_n905__, new_new_n906__, new_new_n907__,
    new_new_n908__, new_new_n909__, new_new_n910__, new_new_n911__,
    new_new_n912__, new_new_n913__, new_new_n914__, new_new_n915__,
    new_new_n916__, new_new_n917__, new_new_n918__, new_new_n919__,
    new_new_n920__, new_new_n921__, new_new_n922__, new_new_n923__,
    new_new_n924__, new_new_n925__, new_new_n926__, new_new_n927__,
    new_new_n928__, new_new_n929__, new_new_n930__, new_new_n931__,
    new_new_n932__, new_new_n933__, new_new_n934__, new_new_n935__,
    new_new_n936__, new_new_n937__, new_new_n938__, new_new_n939__,
    new_new_n940__, new_new_n941__, new_new_n942__, new_new_n943__,
    new_new_n944__, new_new_n945__, new_new_n946__, new_new_n947__,
    new_new_n948__, new_new_n949__, new_new_n950__, new_new_n951__,
    new_new_n952__, new_new_n953__, new_new_n954__, new_new_n955__,
    new_new_n956__, new_new_n957__, new_new_n958__, new_new_n959__,
    new_new_n960__, new_new_n961__, new_new_n962__, new_new_n963__,
    new_new_n964__, new_new_n965__, new_new_n967__, new_new_n968__,
    new_new_n969__, new_new_n970__, new_new_n971__, new_new_n972__,
    new_new_n973__, new_new_n974__, new_new_n975__, new_new_n976__,
    new_new_n977__, new_new_n978__, new_new_n979__, new_new_n980__,
    new_new_n981__, new_new_n982__, new_new_n983__, new_new_n984__,
    new_new_n985__, new_new_n986__, new_new_n987__, new_new_n988__,
    new_new_n989__, new_new_n990__, new_new_n991__, new_new_n992__,
    new_new_n993__, new_new_n994__, new_new_n995__, new_new_n996__,
    new_new_n997__, new_new_n998__, new_new_n999__, new_new_n1000__,
    new_new_n1001__, new_new_n1002__, new_new_n1003__, new_new_n1004__,
    new_new_n1005__, new_new_n1006__, new_new_n1007__, new_new_n1008__,
    new_new_n1009__, new_new_n1010__, new_new_n1011__, new_new_n1012__,
    new_new_n1013__, new_new_n1014__, new_new_n1015__, new_new_n1016__,
    new_new_n1017__, new_new_n1018__, new_new_n1019__, new_new_n1020__,
    new_new_n1021__, new_new_n1022__, new_new_n1023__, new_new_n1024__,
    new_new_n1025__, new_new_n1026__, new_new_n1027__, new_new_n1028__,
    new_new_n1029__, new_new_n1030__, new_new_n1031__, new_new_n1032__,
    new_new_n1033__, new_new_n1034__, new_new_n1035__, new_new_n1036__,
    new_new_n1037__, new_new_n1038__, new_new_n1039__, new_new_n1040__,
    new_new_n1041__, new_new_n1042__, new_new_n1043__, new_new_n1044__,
    new_new_n1045__, new_new_n1046__, new_new_n1047__, new_new_n1048__,
    new_new_n1049__, new_new_n1050__, new_new_n1051__, new_new_n1052__,
    new_new_n1053__, new_new_n1054__, new_new_n1055__, new_new_n1056__,
    new_new_n1057__, new_new_n1058__, new_new_n1059__, new_new_n1060__,
    new_new_n1061__, new_new_n1062__, new_new_n1063__, new_new_n1064__,
    new_new_n1065__, new_new_n1066__, new_new_n1067__, new_new_n1068__,
    new_new_n1069__, new_new_n1070__, new_new_n1071__, new_new_n1072__,
    new_new_n1073__, new_new_n1074__, new_new_n1075__, new_new_n1076__,
    new_new_n1077__, new_new_n1078__, new_new_n1079__, new_new_n1081__,
    new_new_n1082__, new_new_n1083__, new_new_n1084__, new_new_n1085__,
    new_new_n1086__, new_new_n1087__, new_new_n1088__, new_new_n1089__,
    new_new_n1090__, new_new_n1091__, new_new_n1092__, new_new_n1093__,
    new_new_n1094__, new_new_n1095__, new_new_n1096__, new_new_n1097__,
    new_new_n1098__, new_new_n1099__, new_new_n1100__, new_new_n1101__,
    new_new_n1102__, new_new_n1103__, new_new_n1104__, new_new_n1105__,
    new_new_n1106__, new_new_n1107__, new_new_n1108__, new_new_n1109__,
    new_new_n1110__, new_new_n1111__, new_new_n1112__, new_new_n1113__,
    new_new_n1114__, new_new_n1115__, new_new_n1116__, new_new_n1117__,
    new_new_n1118__, new_new_n1119__, new_new_n1120__, new_new_n1121__,
    new_new_n1122__, new_new_n1123__, new_new_n1124__, new_new_n1125__,
    new_new_n1126__, new_new_n1127__, new_new_n1128__, new_new_n1129__,
    new_new_n1130__, new_new_n1131__, new_new_n1132__, new_new_n1133__,
    new_new_n1134__, new_new_n1135__, new_new_n1136__, new_new_n1137__,
    new_new_n1138__, new_new_n1139__, new_new_n1140__, new_new_n1141__,
    new_new_n1142__, new_new_n1143__, new_new_n1144__, new_new_n1145__,
    new_new_n1146__, new_new_n1147__, new_new_n1148__, new_new_n1149__,
    new_new_n1150__, new_new_n1151__, new_new_n1152__, new_new_n1153__,
    new_new_n1154__, new_new_n1155__, new_new_n1156__, new_new_n1157__,
    new_new_n1158__, new_new_n1159__, new_new_n1160__, new_new_n1161__,
    new_new_n1162__, new_new_n1163__, new_new_n1164__, new_new_n1165__,
    new_new_n1166__, new_new_n1167__, new_new_n1168__, new_new_n1169__,
    new_new_n1170__, new_new_n1171__, new_new_n1172__, new_new_n1173__,
    new_new_n1174__, new_new_n1175__, new_new_n1176__, new_new_n1177__,
    new_new_n1178__, new_new_n1179__, new_new_n1180__, new_new_n1181__,
    new_new_n1182__, new_new_n1183__, new_new_n1184__, new_new_n1185__,
    new_new_n1186__, new_new_n1187__, new_new_n1188__, new_new_n1189__,
    new_new_n1190__, new_new_n1191__, new_new_n1193__, new_new_n1194__,
    new_new_n1195__, new_new_n1196__, new_new_n1197__, new_new_n1198__,
    new_new_n1199__, new_new_n1200__, new_new_n1201__, new_new_n1202__,
    new_new_n1203__, new_new_n1204__, new_new_n1205__, new_new_n1206__,
    new_new_n1207__, new_new_n1208__, new_new_n1209__, new_new_n1210__,
    new_new_n1211__, new_new_n1212__, new_new_n1213__, new_new_n1214__,
    new_new_n1215__, new_new_n1216__, new_new_n1217__, new_new_n1218__,
    new_new_n1219__, new_new_n1220__, new_new_n1221__, new_new_n1222__,
    new_new_n1223__, new_new_n1224__, new_new_n1225__, new_new_n1226__,
    new_new_n1227__, new_new_n1228__, new_new_n1229__, new_new_n1230__,
    new_new_n1231__, new_new_n1232__, new_new_n1233__, new_new_n1234__,
    new_new_n1235__, new_new_n1236__, new_new_n1237__, new_new_n1238__,
    new_new_n1239__, new_new_n1240__, new_new_n1241__, new_new_n1242__,
    new_new_n1243__, new_new_n1244__, new_new_n1245__, new_new_n1246__,
    new_new_n1247__, new_new_n1248__, new_new_n1249__, new_new_n1250__,
    new_new_n1251__, new_new_n1252__, new_new_n1253__, new_new_n1254__,
    new_new_n1255__, new_new_n1256__, new_new_n1257__, new_new_n1258__,
    new_new_n1259__, new_new_n1260__, new_new_n1261__, new_new_n1262__,
    new_new_n1263__, new_new_n1264__, new_new_n1265__, new_new_n1266__,
    new_new_n1267__, new_new_n1268__, new_new_n1269__, new_new_n1270__,
    new_new_n1271__, new_new_n1272__, new_new_n1273__, new_new_n1274__,
    new_new_n1275__, new_new_n1276__, new_new_n1277__, new_new_n1278__,
    new_new_n1279__, new_new_n1280__, new_new_n1281__, new_new_n1282__,
    new_new_n1283__, new_new_n1284__, new_new_n1285__, new_new_n1286__,
    new_new_n1287__, new_new_n1288__, new_new_n1289__, new_new_n1290__,
    new_new_n1291__, new_new_n1292__, new_new_n1293__, new_new_n1294__,
    new_new_n1295__, new_new_n1296__, new_new_n1298__, new_new_n1299__,
    new_new_n1300__, new_new_n1301__, new_new_n1302__, new_new_n1303__,
    new_new_n1304__, new_new_n1305__, new_new_n1306__, new_new_n1307__,
    new_new_n1308__, new_new_n1309__, new_new_n1310__, new_new_n1311__,
    new_new_n1312__, new_new_n1313__, new_new_n1314__, new_new_n1315__,
    new_new_n1316__, new_new_n1317__, new_new_n1318__, new_new_n1319__,
    new_new_n1320__, new_new_n1321__, new_new_n1322__, new_new_n1323__,
    new_new_n1324__, new_new_n1325__, new_new_n1326__, new_new_n1327__,
    new_new_n1328__, new_new_n1329__, new_new_n1330__, new_new_n1331__,
    new_new_n1332__, new_new_n1333__, new_new_n1334__, new_new_n1335__,
    new_new_n1336__, new_new_n1337__, new_new_n1338__, new_new_n1339__,
    new_new_n1340__, new_new_n1341__, new_new_n1342__, new_new_n1343__,
    new_new_n1344__, new_new_n1345__, new_new_n1346__, new_new_n1347__,
    new_new_n1348__, new_new_n1349__, new_new_n1350__, new_new_n1351__,
    new_new_n1352__, new_new_n1353__, new_new_n1354__, new_new_n1355__,
    new_new_n1356__, new_new_n1357__, new_new_n1358__, new_new_n1359__,
    new_new_n1360__, new_new_n1361__, new_new_n1362__, new_new_n1363__,
    new_new_n1364__, new_new_n1365__, new_new_n1366__, new_new_n1367__,
    new_new_n1368__, new_new_n1369__, new_new_n1370__, new_new_n1371__,
    new_new_n1372__, new_new_n1373__, new_new_n1374__, new_new_n1375__,
    new_new_n1376__, new_new_n1377__, new_new_n1378__, new_new_n1379__,
    new_new_n1380__, new_new_n1381__, new_new_n1382__, new_new_n1383__,
    new_new_n1384__, new_new_n1385__, new_new_n1386__, new_new_n1387__,
    new_new_n1388__, new_new_n1389__, new_new_n1390__, new_new_n1391__,
    new_new_n1392__, new_new_n1393__, new_new_n1395__, new_new_n1396__,
    new_new_n1397__, new_new_n1398__, new_new_n1399__, new_new_n1400__,
    new_new_n1401__, new_new_n1402__, new_new_n1403__, new_new_n1404__,
    new_new_n1405__, new_new_n1406__, new_new_n1407__, new_new_n1408__,
    new_new_n1409__, new_new_n1410__, new_new_n1411__, new_new_n1412__,
    new_new_n1413__, new_new_n1414__, new_new_n1415__, new_new_n1416__,
    new_new_n1417__, new_new_n1418__, new_new_n1419__, new_new_n1420__,
    new_new_n1421__, new_new_n1422__, new_new_n1423__, new_new_n1424__,
    new_new_n1425__, new_new_n1426__, new_new_n1427__, new_new_n1428__,
    new_new_n1429__, new_new_n1430__, new_new_n1431__, new_new_n1432__,
    new_new_n1433__, new_new_n1434__, new_new_n1435__, new_new_n1436__,
    new_new_n1437__, new_new_n1438__, new_new_n1439__, new_new_n1440__,
    new_new_n1441__, new_new_n1442__, new_new_n1443__, new_new_n1444__,
    new_new_n1445__, new_new_n1446__, new_new_n1447__, new_new_n1448__,
    new_new_n1449__, new_new_n1450__, new_new_n1451__, new_new_n1452__,
    new_new_n1453__, new_new_n1454__, new_new_n1455__, new_new_n1456__,
    new_new_n1457__, new_new_n1458__, new_new_n1459__, new_new_n1460__,
    new_new_n1461__, new_new_n1462__, new_new_n1463__, new_new_n1464__,
    new_new_n1465__, new_new_n1466__, new_new_n1467__, new_new_n1468__,
    new_new_n1469__, new_new_n1470__, new_new_n1471__, new_new_n1472__,
    new_new_n1473__, new_new_n1474__, new_new_n1475__, new_new_n1476__,
    new_new_n1477__, new_new_n1478__, new_new_n1479__, new_new_n1480__,
    new_new_n1481__, new_new_n1482__, new_new_n1484__, new_new_n1485__,
    new_new_n1486__, new_new_n1487__, new_new_n1488__, new_new_n1489__,
    new_new_n1490__, new_new_n1491__, new_new_n1492__, new_new_n1493__,
    new_new_n1494__, new_new_n1495__, new_new_n1496__, new_new_n1497__,
    new_new_n1498__, new_new_n1499__, new_new_n1500__, new_new_n1501__,
    new_new_n1502__, new_new_n1503__, new_new_n1504__, new_new_n1505__,
    new_new_n1506__, new_new_n1507__, new_new_n1508__, new_new_n1509__,
    new_new_n1510__, new_new_n1511__, new_new_n1512__, new_new_n1513__,
    new_new_n1514__, new_new_n1515__, new_new_n1516__, new_new_n1517__,
    new_new_n1518__, new_new_n1519__, new_new_n1520__, new_new_n1521__,
    new_new_n1522__, new_new_n1523__, new_new_n1524__, new_new_n1525__,
    new_new_n1526__, new_new_n1527__, new_new_n1528__, new_new_n1529__,
    new_new_n1530__, new_new_n1531__, new_new_n1532__, new_new_n1533__,
    new_new_n1534__, new_new_n1535__, new_new_n1536__, new_new_n1537__,
    new_new_n1538__, new_new_n1539__, new_new_n1540__, new_new_n1541__,
    new_new_n1542__, new_new_n1543__, new_new_n1544__, new_new_n1545__,
    new_new_n1546__, new_new_n1547__, new_new_n1548__, new_new_n1549__,
    new_new_n1550__, new_new_n1551__, new_new_n1552__, new_new_n1553__,
    new_new_n1554__, new_new_n1555__, new_new_n1556__, new_new_n1557__,
    new_new_n1558__, new_new_n1559__, new_new_n1560__, new_new_n1561__,
    new_new_n1562__, new_new_n1563__, new_new_n1565__, new_new_n1566__,
    new_new_n1567__, new_new_n1568__, new_new_n1569__, new_new_n1570__,
    new_new_n1571__, new_new_n1572__, new_new_n1573__, new_new_n1574__,
    new_new_n1575__, new_new_n1576__, new_new_n1577__, new_new_n1578__,
    new_new_n1579__, new_new_n1580__, new_new_n1581__, new_new_n1582__,
    new_new_n1583__, new_new_n1584__, new_new_n1585__, new_new_n1586__,
    new_new_n1587__, new_new_n1588__, new_new_n1589__, new_new_n1590__,
    new_new_n1591__, new_new_n1592__, new_new_n1593__, new_new_n1594__,
    new_new_n1595__, new_new_n1596__, new_new_n1597__, new_new_n1598__,
    new_new_n1599__, new_new_n1600__, new_new_n1601__, new_new_n1602__,
    new_new_n1603__, new_new_n1604__, new_new_n1605__, new_new_n1606__,
    new_new_n1607__, new_new_n1608__, new_new_n1609__, new_new_n1610__,
    new_new_n1611__, new_new_n1612__, new_new_n1613__, new_new_n1614__,
    new_new_n1615__, new_new_n1616__, new_new_n1617__, new_new_n1618__,
    new_new_n1619__, new_new_n1620__, new_new_n1621__, new_new_n1622__,
    new_new_n1623__, new_new_n1624__, new_new_n1625__, new_new_n1626__,
    new_new_n1627__, new_new_n1628__, new_new_n1629__, new_new_n1630__,
    new_new_n1631__, new_new_n1632__, new_new_n1633__, new_new_n1634__,
    new_new_n1635__, new_new_n1636__, new_new_n1638__, new_new_n1639__,
    new_new_n1640__, new_new_n1641__, new_new_n1642__, new_new_n1643__,
    new_new_n1644__, new_new_n1645__, new_new_n1646__, new_new_n1647__,
    new_new_n1648__, new_new_n1649__, new_new_n1650__, new_new_n1651__,
    new_new_n1652__, new_new_n1653__, new_new_n1654__, new_new_n1655__,
    new_new_n1656__, new_new_n1657__, new_new_n1658__, new_new_n1659__,
    new_new_n1660__, new_new_n1661__, new_new_n1662__, new_new_n1663__,
    new_new_n1664__, new_new_n1665__, new_new_n1666__, new_new_n1667__,
    new_new_n1668__, new_new_n1669__, new_new_n1670__, new_new_n1671__,
    new_new_n1672__, new_new_n1673__, new_new_n1674__, new_new_n1675__,
    new_new_n1676__, new_new_n1677__, new_new_n1678__, new_new_n1679__,
    new_new_n1680__, new_new_n1681__, new_new_n1682__, new_new_n1683__,
    new_new_n1684__, new_new_n1685__, new_new_n1686__, new_new_n1687__,
    new_new_n1688__, new_new_n1689__, new_new_n1690__, new_new_n1691__,
    new_new_n1692__, new_new_n1693__, new_new_n1694__, new_new_n1695__,
    new_new_n1696__, new_new_n1697__, new_new_n1698__, new_new_n1699__,
    new_new_n1700__, new_new_n1701__, new_new_n1703__, new_new_n1704__,
    new_new_n1705__, new_new_n1706__, new_new_n1707__, new_new_n1708__,
    new_new_n1709__, new_new_n1710__, new_new_n1711__, new_new_n1712__,
    new_new_n1713__, new_new_n1714__, new_new_n1715__, new_new_n1716__,
    new_new_n1717__, new_new_n1718__, new_new_n1719__, new_new_n1720__,
    new_new_n1721__, new_new_n1722__, new_new_n1723__, new_new_n1724__,
    new_new_n1725__, new_new_n1726__, new_new_n1727__, new_new_n1728__,
    new_new_n1729__, new_new_n1730__, new_new_n1731__, new_new_n1732__,
    new_new_n1733__, new_new_n1734__, new_new_n1735__, new_new_n1736__,
    new_new_n1737__, new_new_n1738__, new_new_n1739__, new_new_n1740__,
    new_new_n1741__, new_new_n1742__, new_new_n1743__, new_new_n1744__,
    new_new_n1745__, new_new_n1746__, new_new_n1747__, new_new_n1748__,
    new_new_n1749__, new_new_n1750__, new_new_n1751__, new_new_n1752__,
    new_new_n1753__, new_new_n1754__, new_new_n1755__, new_new_n1756__,
    new_new_n1757__, new_new_n1758__, new_new_n1760__, new_new_n1761__,
    new_new_n1762__, new_new_n1763__, new_new_n1764__, new_new_n1765__,
    new_new_n1766__, new_new_n1767__, new_new_n1768__, new_new_n1769__,
    new_new_n1770__, new_new_n1771__, new_new_n1772__, new_new_n1773__,
    new_new_n1774__, new_new_n1775__, new_new_n1776__, new_new_n1777__,
    new_new_n1778__, new_new_n1779__, new_new_n1780__, new_new_n1781__,
    new_new_n1782__, new_new_n1783__, new_new_n1784__, new_new_n1785__,
    new_new_n1786__, new_new_n1787__, new_new_n1788__, new_new_n1789__,
    new_new_n1790__, new_new_n1791__, new_new_n1792__, new_new_n1793__,
    new_new_n1794__, new_new_n1795__, new_new_n1796__, new_new_n1797__,
    new_new_n1798__, new_new_n1799__, new_new_n1800__, new_new_n1801__,
    new_new_n1802__, new_new_n1803__, new_new_n1804__, new_new_n1805__,
    new_new_n1806__, new_new_n1807__, new_new_n1809__, new_new_n1810__,
    new_new_n1811__, new_new_n1812__, new_new_n1813__, new_new_n1814__,
    new_new_n1815__, new_new_n1816__, new_new_n1817__, new_new_n1818__,
    new_new_n1819__, new_new_n1820__, new_new_n1821__, new_new_n1822__,
    new_new_n1823__, new_new_n1824__, new_new_n1825__, new_new_n1826__,
    new_new_n1827__, new_new_n1828__, new_new_n1829__, new_new_n1830__,
    new_new_n1831__, new_new_n1832__, new_new_n1833__, new_new_n1834__,
    new_new_n1835__, new_new_n1836__, new_new_n1837__, new_new_n1838__,
    new_new_n1839__, new_new_n1840__, new_new_n1841__, new_new_n1842__,
    new_new_n1843__, new_new_n1844__, new_new_n1845__, new_new_n1846__,
    new_new_n1847__, new_new_n1848__, new_new_n1850__, new_new_n1851__,
    new_new_n1852__, new_new_n1853__, new_new_n1854__, new_new_n1855__,
    new_new_n1856__, new_new_n1857__, new_new_n1858__, new_new_n1859__,
    new_new_n1860__, new_new_n1861__, new_new_n1862__, new_new_n1863__,
    new_new_n1864__, new_new_n1865__, new_new_n1866__, new_new_n1867__,
    new_new_n1868__, new_new_n1869__, new_new_n1870__, new_new_n1871__,
    new_new_n1872__, new_new_n1873__, new_new_n1874__, new_new_n1875__,
    new_new_n1876__, new_new_n1877__, new_new_n1878__, new_new_n1879__,
    new_new_n1880__, new_new_n1881__, new_new_n1883__, new_new_n1884__,
    new_new_n1885__, new_new_n1886__, new_new_n1887__, new_new_n1888__,
    new_new_n1889__, new_new_n1890__, new_new_n1891__, new_new_n1892__,
    new_new_n1893__, new_new_n1894__, new_new_n1895__, new_new_n1896__,
    new_new_n1897__, new_new_n1898__, new_new_n1899__, new_new_n1900__,
    new_new_n1901__, new_new_n1902__, new_new_n1903__, new_new_n1904__,
    new_new_n1905__, new_new_n1906__, new_new_n1908__, new_new_n1909__,
    new_new_n1910__, new_new_n1911__, new_new_n1912__, new_new_n1913__,
    new_new_n1914__, new_new_n1915__, new_new_n1916__, new_new_n1917__,
    new_new_n1918__, new_new_n1919__, new_new_n1920__, new_new_n1921__,
    new_new_n1922__, new_new_n1923__, new_new_n1925__, new_new_n1926__,
    new_new_n1927__, new_new_n1928__, new_new_n1929__, new_new_n1930__,
    new_new_n1931__, new_new_n1933__;
  assign G545gat = G1gat & G273gat;
  assign new_new_n66__ = G18gat & G273gat;
  assign new_new_n67__ = G1gat & G290gat;
  assign new_new_n68__ = ~new_new_n66__ & ~new_new_n67__;
  assign new_new_n69__ = G18gat & G290gat;
  assign new_new_n70__ = G545gat & new_new_n69__;
  assign G1581gat = ~new_new_n68__ & ~new_new_n70__;
  assign new_new_n72__ = G1gat & G307gat;
  assign new_new_n73__ = G35gat & G273gat;
  assign new_new_n74__ = ~new_new_n69__ & ~new_new_n73__;
  assign new_new_n75__ = G35gat & G290gat;
  assign new_new_n76__ = new_new_n66__ & new_new_n75__;
  assign new_new_n77__ = ~new_new_n74__ & ~new_new_n76__;
  assign new_new_n78__ = ~new_new_n70__ & ~new_new_n77__;
  assign new_new_n79__ = new_new_n70__ & ~new_new_n76__;
  assign new_new_n80__ = ~new_new_n78__ & ~new_new_n79__;
  assign new_new_n81__ = ~new_new_n72__ & new_new_n80__;
  assign new_new_n82__ = new_new_n72__ & ~new_new_n80__;
  assign G1901gat = new_new_n81__ | new_new_n82__;
  assign new_new_n84__ = G1gat & G324gat;
  assign new_new_n85__ = ~new_new_n78__ & ~new_new_n81__;
  assign new_new_n86__ = G18gat & G307gat;
  assign new_new_n87__ = G52gat & G273gat;
  assign new_new_n88__ = ~new_new_n75__ & ~new_new_n87__;
  assign new_new_n89__ = G52gat & G290gat;
  assign new_new_n90__ = new_new_n73__ & new_new_n89__;
  assign new_new_n91__ = ~new_new_n88__ & ~new_new_n90__;
  assign new_new_n92__ = ~new_new_n76__ & ~new_new_n91__;
  assign new_new_n93__ = new_new_n76__ & ~new_new_n90__;
  assign new_new_n94__ = ~new_new_n92__ & ~new_new_n93__;
  assign new_new_n95__ = ~new_new_n86__ & new_new_n94__;
  assign new_new_n96__ = new_new_n86__ & ~new_new_n94__;
  assign new_new_n97__ = ~new_new_n95__ & ~new_new_n96__;
  assign new_new_n98__ = ~new_new_n85__ & new_new_n97__;
  assign new_new_n99__ = new_new_n85__ & ~new_new_n97__;
  assign new_new_n100__ = ~new_new_n98__ & ~new_new_n99__;
  assign new_new_n101__ = ~new_new_n84__ & new_new_n100__;
  assign new_new_n102__ = new_new_n84__ & ~new_new_n100__;
  assign G2223gat = new_new_n101__ | new_new_n102__;
  assign new_new_n104__ = G1gat & G341gat;
  assign new_new_n105__ = ~new_new_n98__ & ~new_new_n101__;
  assign new_new_n106__ = G18gat & G324gat;
  assign new_new_n107__ = ~new_new_n92__ & ~new_new_n95__;
  assign new_new_n108__ = G35gat & G307gat;
  assign new_new_n109__ = G69gat & G273gat;
  assign new_new_n110__ = ~new_new_n89__ & ~new_new_n109__;
  assign new_new_n111__ = G69gat & G290gat;
  assign new_new_n112__ = new_new_n87__ & new_new_n111__;
  assign new_new_n113__ = ~new_new_n110__ & ~new_new_n112__;
  assign new_new_n114__ = ~new_new_n90__ & ~new_new_n113__;
  assign new_new_n115__ = new_new_n90__ & ~new_new_n112__;
  assign new_new_n116__ = ~new_new_n114__ & ~new_new_n115__;
  assign new_new_n117__ = ~new_new_n108__ & new_new_n116__;
  assign new_new_n118__ = new_new_n108__ & ~new_new_n116__;
  assign new_new_n119__ = ~new_new_n117__ & ~new_new_n118__;
  assign new_new_n120__ = ~new_new_n107__ & new_new_n119__;
  assign new_new_n121__ = new_new_n107__ & ~new_new_n119__;
  assign new_new_n122__ = ~new_new_n120__ & ~new_new_n121__;
  assign new_new_n123__ = ~new_new_n106__ & new_new_n122__;
  assign new_new_n124__ = new_new_n106__ & ~new_new_n122__;
  assign new_new_n125__ = ~new_new_n123__ & ~new_new_n124__;
  assign new_new_n126__ = ~new_new_n105__ & new_new_n125__;
  assign new_new_n127__ = new_new_n105__ & ~new_new_n125__;
  assign new_new_n128__ = ~new_new_n126__ & ~new_new_n127__;
  assign new_new_n129__ = ~new_new_n104__ & new_new_n128__;
  assign new_new_n130__ = new_new_n104__ & ~new_new_n128__;
  assign G2548gat = new_new_n129__ | new_new_n130__;
  assign new_new_n132__ = G1gat & G358gat;
  assign new_new_n133__ = ~new_new_n126__ & ~new_new_n129__;
  assign new_new_n134__ = G18gat & G341gat;
  assign new_new_n135__ = ~new_new_n120__ & ~new_new_n123__;
  assign new_new_n136__ = G35gat & G324gat;
  assign new_new_n137__ = ~new_new_n114__ & ~new_new_n117__;
  assign new_new_n138__ = G52gat & G307gat;
  assign new_new_n139__ = G86gat & G273gat;
  assign new_new_n140__ = ~new_new_n111__ & ~new_new_n139__;
  assign new_new_n141__ = G86gat & G290gat;
  assign new_new_n142__ = new_new_n109__ & new_new_n141__;
  assign new_new_n143__ = ~new_new_n140__ & ~new_new_n142__;
  assign new_new_n144__ = ~new_new_n112__ & ~new_new_n143__;
  assign new_new_n145__ = new_new_n112__ & ~new_new_n142__;
  assign new_new_n146__ = ~new_new_n144__ & ~new_new_n145__;
  assign new_new_n147__ = ~new_new_n138__ & new_new_n146__;
  assign new_new_n148__ = new_new_n138__ & ~new_new_n146__;
  assign new_new_n149__ = ~new_new_n147__ & ~new_new_n148__;
  assign new_new_n150__ = ~new_new_n137__ & new_new_n149__;
  assign new_new_n151__ = new_new_n137__ & ~new_new_n149__;
  assign new_new_n152__ = ~new_new_n150__ & ~new_new_n151__;
  assign new_new_n153__ = ~new_new_n136__ & new_new_n152__;
  assign new_new_n154__ = new_new_n136__ & ~new_new_n152__;
  assign new_new_n155__ = ~new_new_n153__ & ~new_new_n154__;
  assign new_new_n156__ = ~new_new_n135__ & new_new_n155__;
  assign new_new_n157__ = new_new_n135__ & ~new_new_n155__;
  assign new_new_n158__ = ~new_new_n156__ & ~new_new_n157__;
  assign new_new_n159__ = ~new_new_n134__ & new_new_n158__;
  assign new_new_n160__ = new_new_n134__ & ~new_new_n158__;
  assign new_new_n161__ = ~new_new_n159__ & ~new_new_n160__;
  assign new_new_n162__ = ~new_new_n133__ & new_new_n161__;
  assign new_new_n163__ = new_new_n133__ & ~new_new_n161__;
  assign new_new_n164__ = ~new_new_n162__ & ~new_new_n163__;
  assign new_new_n165__ = ~new_new_n132__ & new_new_n164__;
  assign new_new_n166__ = new_new_n132__ & ~new_new_n164__;
  assign G2877gat = new_new_n165__ | new_new_n166__;
  assign new_new_n168__ = G1gat & G375gat;
  assign new_new_n169__ = ~new_new_n162__ & ~new_new_n165__;
  assign new_new_n170__ = G18gat & G358gat;
  assign new_new_n171__ = ~new_new_n156__ & ~new_new_n159__;
  assign new_new_n172__ = G35gat & G341gat;
  assign new_new_n173__ = ~new_new_n150__ & ~new_new_n153__;
  assign new_new_n174__ = G52gat & G324gat;
  assign new_new_n175__ = ~new_new_n144__ & ~new_new_n147__;
  assign new_new_n176__ = G69gat & G307gat;
  assign new_new_n177__ = G103gat & G273gat;
  assign new_new_n178__ = ~new_new_n141__ & ~new_new_n177__;
  assign new_new_n179__ = G103gat & G290gat;
  assign new_new_n180__ = new_new_n139__ & new_new_n179__;
  assign new_new_n181__ = ~new_new_n178__ & ~new_new_n180__;
  assign new_new_n182__ = ~new_new_n142__ & ~new_new_n181__;
  assign new_new_n183__ = new_new_n142__ & ~new_new_n180__;
  assign new_new_n184__ = ~new_new_n182__ & ~new_new_n183__;
  assign new_new_n185__ = ~new_new_n176__ & new_new_n184__;
  assign new_new_n186__ = new_new_n176__ & ~new_new_n184__;
  assign new_new_n187__ = ~new_new_n185__ & ~new_new_n186__;
  assign new_new_n188__ = ~new_new_n175__ & new_new_n187__;
  assign new_new_n189__ = new_new_n175__ & ~new_new_n187__;
  assign new_new_n190__ = ~new_new_n188__ & ~new_new_n189__;
  assign new_new_n191__ = ~new_new_n174__ & new_new_n190__;
  assign new_new_n192__ = new_new_n174__ & ~new_new_n190__;
  assign new_new_n193__ = ~new_new_n191__ & ~new_new_n192__;
  assign new_new_n194__ = ~new_new_n173__ & new_new_n193__;
  assign new_new_n195__ = new_new_n173__ & ~new_new_n193__;
  assign new_new_n196__ = ~new_new_n194__ & ~new_new_n195__;
  assign new_new_n197__ = ~new_new_n172__ & new_new_n196__;
  assign new_new_n198__ = new_new_n172__ & ~new_new_n196__;
  assign new_new_n199__ = ~new_new_n197__ & ~new_new_n198__;
  assign new_new_n200__ = ~new_new_n171__ & new_new_n199__;
  assign new_new_n201__ = new_new_n171__ & ~new_new_n199__;
  assign new_new_n202__ = ~new_new_n200__ & ~new_new_n201__;
  assign new_new_n203__ = ~new_new_n170__ & new_new_n202__;
  assign new_new_n204__ = new_new_n170__ & ~new_new_n202__;
  assign new_new_n205__ = ~new_new_n203__ & ~new_new_n204__;
  assign new_new_n206__ = ~new_new_n169__ & new_new_n205__;
  assign new_new_n207__ = new_new_n169__ & ~new_new_n205__;
  assign new_new_n208__ = ~new_new_n206__ & ~new_new_n207__;
  assign new_new_n209__ = ~new_new_n168__ & new_new_n208__;
  assign new_new_n210__ = new_new_n168__ & ~new_new_n208__;
  assign G3211gat = new_new_n209__ | new_new_n210__;
  assign new_new_n212__ = G1gat & G392gat;
  assign new_new_n213__ = ~new_new_n206__ & ~new_new_n209__;
  assign new_new_n214__ = G18gat & G375gat;
  assign new_new_n215__ = ~new_new_n200__ & ~new_new_n203__;
  assign new_new_n216__ = G35gat & G358gat;
  assign new_new_n217__ = ~new_new_n194__ & ~new_new_n197__;
  assign new_new_n218__ = G52gat & G341gat;
  assign new_new_n219__ = ~new_new_n188__ & ~new_new_n191__;
  assign new_new_n220__ = G69gat & G324gat;
  assign new_new_n221__ = ~new_new_n182__ & ~new_new_n185__;
  assign new_new_n222__ = G86gat & G307gat;
  assign new_new_n223__ = G120gat & G273gat;
  assign new_new_n224__ = ~new_new_n179__ & ~new_new_n223__;
  assign new_new_n225__ = G120gat & G290gat;
  assign new_new_n226__ = new_new_n177__ & new_new_n225__;
  assign new_new_n227__ = ~new_new_n224__ & ~new_new_n226__;
  assign new_new_n228__ = ~new_new_n180__ & ~new_new_n227__;
  assign new_new_n229__ = new_new_n180__ & ~new_new_n226__;
  assign new_new_n230__ = ~new_new_n228__ & ~new_new_n229__;
  assign new_new_n231__ = ~new_new_n222__ & new_new_n230__;
  assign new_new_n232__ = new_new_n222__ & ~new_new_n230__;
  assign new_new_n233__ = ~new_new_n231__ & ~new_new_n232__;
  assign new_new_n234__ = ~new_new_n221__ & new_new_n233__;
  assign new_new_n235__ = new_new_n221__ & ~new_new_n233__;
  assign new_new_n236__ = ~new_new_n234__ & ~new_new_n235__;
  assign new_new_n237__ = ~new_new_n220__ & new_new_n236__;
  assign new_new_n238__ = new_new_n220__ & ~new_new_n236__;
  assign new_new_n239__ = ~new_new_n237__ & ~new_new_n238__;
  assign new_new_n240__ = ~new_new_n219__ & new_new_n239__;
  assign new_new_n241__ = new_new_n219__ & ~new_new_n239__;
  assign new_new_n242__ = ~new_new_n240__ & ~new_new_n241__;
  assign new_new_n243__ = ~new_new_n218__ & new_new_n242__;
  assign new_new_n244__ = new_new_n218__ & ~new_new_n242__;
  assign new_new_n245__ = ~new_new_n243__ & ~new_new_n244__;
  assign new_new_n246__ = ~new_new_n217__ & new_new_n245__;
  assign new_new_n247__ = new_new_n217__ & ~new_new_n245__;
  assign new_new_n248__ = ~new_new_n246__ & ~new_new_n247__;
  assign new_new_n249__ = ~new_new_n216__ & new_new_n248__;
  assign new_new_n250__ = new_new_n216__ & ~new_new_n248__;
  assign new_new_n251__ = ~new_new_n249__ & ~new_new_n250__;
  assign new_new_n252__ = ~new_new_n215__ & new_new_n251__;
  assign new_new_n253__ = new_new_n215__ & ~new_new_n251__;
  assign new_new_n254__ = ~new_new_n252__ & ~new_new_n253__;
  assign new_new_n255__ = ~new_new_n214__ & new_new_n254__;
  assign new_new_n256__ = new_new_n214__ & ~new_new_n254__;
  assign new_new_n257__ = ~new_new_n255__ & ~new_new_n256__;
  assign new_new_n258__ = ~new_new_n213__ & new_new_n257__;
  assign new_new_n259__ = new_new_n213__ & ~new_new_n257__;
  assign new_new_n260__ = ~new_new_n258__ & ~new_new_n259__;
  assign new_new_n261__ = ~new_new_n212__ & new_new_n260__;
  assign new_new_n262__ = new_new_n212__ & ~new_new_n260__;
  assign G3552gat = new_new_n261__ | new_new_n262__;
  assign new_new_n264__ = G1gat & G409gat;
  assign new_new_n265__ = ~new_new_n258__ & ~new_new_n261__;
  assign new_new_n266__ = G18gat & G392gat;
  assign new_new_n267__ = ~new_new_n252__ & ~new_new_n255__;
  assign new_new_n268__ = G35gat & G375gat;
  assign new_new_n269__ = ~new_new_n246__ & ~new_new_n249__;
  assign new_new_n270__ = G52gat & G358gat;
  assign new_new_n271__ = ~new_new_n240__ & ~new_new_n243__;
  assign new_new_n272__ = G69gat & G341gat;
  assign new_new_n273__ = ~new_new_n234__ & ~new_new_n237__;
  assign new_new_n274__ = G86gat & G324gat;
  assign new_new_n275__ = ~new_new_n228__ & ~new_new_n231__;
  assign new_new_n276__ = G103gat & G307gat;
  assign new_new_n277__ = G137gat & G273gat;
  assign new_new_n278__ = ~new_new_n225__ & ~new_new_n277__;
  assign new_new_n279__ = G137gat & G290gat;
  assign new_new_n280__ = new_new_n223__ & new_new_n279__;
  assign new_new_n281__ = ~new_new_n278__ & ~new_new_n280__;
  assign new_new_n282__ = ~new_new_n226__ & ~new_new_n281__;
  assign new_new_n283__ = new_new_n226__ & ~new_new_n280__;
  assign new_new_n284__ = ~new_new_n282__ & ~new_new_n283__;
  assign new_new_n285__ = ~new_new_n276__ & new_new_n284__;
  assign new_new_n286__ = new_new_n276__ & ~new_new_n284__;
  assign new_new_n287__ = ~new_new_n285__ & ~new_new_n286__;
  assign new_new_n288__ = ~new_new_n275__ & new_new_n287__;
  assign new_new_n289__ = new_new_n275__ & ~new_new_n287__;
  assign new_new_n290__ = ~new_new_n288__ & ~new_new_n289__;
  assign new_new_n291__ = ~new_new_n274__ & new_new_n290__;
  assign new_new_n292__ = new_new_n274__ & ~new_new_n290__;
  assign new_new_n293__ = ~new_new_n291__ & ~new_new_n292__;
  assign new_new_n294__ = ~new_new_n273__ & new_new_n293__;
  assign new_new_n295__ = new_new_n273__ & ~new_new_n293__;
  assign new_new_n296__ = ~new_new_n294__ & ~new_new_n295__;
  assign new_new_n297__ = ~new_new_n272__ & new_new_n296__;
  assign new_new_n298__ = new_new_n272__ & ~new_new_n296__;
  assign new_new_n299__ = ~new_new_n297__ & ~new_new_n298__;
  assign new_new_n300__ = ~new_new_n271__ & new_new_n299__;
  assign new_new_n301__ = new_new_n271__ & ~new_new_n299__;
  assign new_new_n302__ = ~new_new_n300__ & ~new_new_n301__;
  assign new_new_n303__ = ~new_new_n270__ & new_new_n302__;
  assign new_new_n304__ = new_new_n270__ & ~new_new_n302__;
  assign new_new_n305__ = ~new_new_n303__ & ~new_new_n304__;
  assign new_new_n306__ = ~new_new_n269__ & new_new_n305__;
  assign new_new_n307__ = new_new_n269__ & ~new_new_n305__;
  assign new_new_n308__ = ~new_new_n306__ & ~new_new_n307__;
  assign new_new_n309__ = ~new_new_n268__ & new_new_n308__;
  assign new_new_n310__ = new_new_n268__ & ~new_new_n308__;
  assign new_new_n311__ = ~new_new_n309__ & ~new_new_n310__;
  assign new_new_n312__ = ~new_new_n267__ & new_new_n311__;
  assign new_new_n313__ = new_new_n267__ & ~new_new_n311__;
  assign new_new_n314__ = ~new_new_n312__ & ~new_new_n313__;
  assign new_new_n315__ = ~new_new_n266__ & new_new_n314__;
  assign new_new_n316__ = new_new_n266__ & ~new_new_n314__;
  assign new_new_n317__ = ~new_new_n315__ & ~new_new_n316__;
  assign new_new_n318__ = ~new_new_n265__ & new_new_n317__;
  assign new_new_n319__ = new_new_n265__ & ~new_new_n317__;
  assign new_new_n320__ = ~new_new_n318__ & ~new_new_n319__;
  assign new_new_n321__ = ~new_new_n264__ & new_new_n320__;
  assign new_new_n322__ = new_new_n264__ & ~new_new_n320__;
  assign G3895gat = new_new_n321__ | new_new_n322__;
  assign new_new_n324__ = G1gat & G426gat;
  assign new_new_n325__ = ~new_new_n318__ & ~new_new_n321__;
  assign new_new_n326__ = G18gat & G409gat;
  assign new_new_n327__ = ~new_new_n312__ & ~new_new_n315__;
  assign new_new_n328__ = G35gat & G392gat;
  assign new_new_n329__ = ~new_new_n306__ & ~new_new_n309__;
  assign new_new_n330__ = G52gat & G375gat;
  assign new_new_n331__ = ~new_new_n300__ & ~new_new_n303__;
  assign new_new_n332__ = G69gat & G358gat;
  assign new_new_n333__ = ~new_new_n294__ & ~new_new_n297__;
  assign new_new_n334__ = G86gat & G341gat;
  assign new_new_n335__ = ~new_new_n288__ & ~new_new_n291__;
  assign new_new_n336__ = G103gat & G324gat;
  assign new_new_n337__ = ~new_new_n282__ & ~new_new_n285__;
  assign new_new_n338__ = G120gat & G307gat;
  assign new_new_n339__ = G154gat & G273gat;
  assign new_new_n340__ = ~new_new_n279__ & ~new_new_n339__;
  assign new_new_n341__ = G154gat & G290gat;
  assign new_new_n342__ = new_new_n277__ & new_new_n341__;
  assign new_new_n343__ = ~new_new_n340__ & ~new_new_n342__;
  assign new_new_n344__ = ~new_new_n280__ & ~new_new_n343__;
  assign new_new_n345__ = new_new_n280__ & ~new_new_n342__;
  assign new_new_n346__ = ~new_new_n344__ & ~new_new_n345__;
  assign new_new_n347__ = ~new_new_n338__ & new_new_n346__;
  assign new_new_n348__ = new_new_n338__ & ~new_new_n346__;
  assign new_new_n349__ = ~new_new_n347__ & ~new_new_n348__;
  assign new_new_n350__ = ~new_new_n337__ & new_new_n349__;
  assign new_new_n351__ = new_new_n337__ & ~new_new_n349__;
  assign new_new_n352__ = ~new_new_n350__ & ~new_new_n351__;
  assign new_new_n353__ = ~new_new_n336__ & new_new_n352__;
  assign new_new_n354__ = new_new_n336__ & ~new_new_n352__;
  assign new_new_n355__ = ~new_new_n353__ & ~new_new_n354__;
  assign new_new_n356__ = ~new_new_n335__ & new_new_n355__;
  assign new_new_n357__ = new_new_n335__ & ~new_new_n355__;
  assign new_new_n358__ = ~new_new_n356__ & ~new_new_n357__;
  assign new_new_n359__ = ~new_new_n334__ & new_new_n358__;
  assign new_new_n360__ = new_new_n334__ & ~new_new_n358__;
  assign new_new_n361__ = ~new_new_n359__ & ~new_new_n360__;
  assign new_new_n362__ = ~new_new_n333__ & new_new_n361__;
  assign new_new_n363__ = new_new_n333__ & ~new_new_n361__;
  assign new_new_n364__ = ~new_new_n362__ & ~new_new_n363__;
  assign new_new_n365__ = ~new_new_n332__ & new_new_n364__;
  assign new_new_n366__ = new_new_n332__ & ~new_new_n364__;
  assign new_new_n367__ = ~new_new_n365__ & ~new_new_n366__;
  assign new_new_n368__ = ~new_new_n331__ & new_new_n367__;
  assign new_new_n369__ = new_new_n331__ & ~new_new_n367__;
  assign new_new_n370__ = ~new_new_n368__ & ~new_new_n369__;
  assign new_new_n371__ = ~new_new_n330__ & new_new_n370__;
  assign new_new_n372__ = new_new_n330__ & ~new_new_n370__;
  assign new_new_n373__ = ~new_new_n371__ & ~new_new_n372__;
  assign new_new_n374__ = ~new_new_n329__ & new_new_n373__;
  assign new_new_n375__ = new_new_n329__ & ~new_new_n373__;
  assign new_new_n376__ = ~new_new_n374__ & ~new_new_n375__;
  assign new_new_n377__ = ~new_new_n328__ & new_new_n376__;
  assign new_new_n378__ = new_new_n328__ & ~new_new_n376__;
  assign new_new_n379__ = ~new_new_n377__ & ~new_new_n378__;
  assign new_new_n380__ = ~new_new_n327__ & new_new_n379__;
  assign new_new_n381__ = new_new_n327__ & ~new_new_n379__;
  assign new_new_n382__ = ~new_new_n380__ & ~new_new_n381__;
  assign new_new_n383__ = ~new_new_n326__ & new_new_n382__;
  assign new_new_n384__ = new_new_n326__ & ~new_new_n382__;
  assign new_new_n385__ = ~new_new_n383__ & ~new_new_n384__;
  assign new_new_n386__ = ~new_new_n325__ & new_new_n385__;
  assign new_new_n387__ = new_new_n325__ & ~new_new_n385__;
  assign new_new_n388__ = ~new_new_n386__ & ~new_new_n387__;
  assign new_new_n389__ = ~new_new_n324__ & new_new_n388__;
  assign new_new_n390__ = new_new_n324__ & ~new_new_n388__;
  assign G4241gat = new_new_n389__ | new_new_n390__;
  assign new_new_n392__ = G1gat & G443gat;
  assign new_new_n393__ = ~new_new_n386__ & ~new_new_n389__;
  assign new_new_n394__ = G18gat & G426gat;
  assign new_new_n395__ = ~new_new_n380__ & ~new_new_n383__;
  assign new_new_n396__ = G35gat & G409gat;
  assign new_new_n397__ = ~new_new_n374__ & ~new_new_n377__;
  assign new_new_n398__ = G52gat & G392gat;
  assign new_new_n399__ = ~new_new_n368__ & ~new_new_n371__;
  assign new_new_n400__ = G69gat & G375gat;
  assign new_new_n401__ = ~new_new_n362__ & ~new_new_n365__;
  assign new_new_n402__ = G86gat & G358gat;
  assign new_new_n403__ = ~new_new_n356__ & ~new_new_n359__;
  assign new_new_n404__ = G103gat & G341gat;
  assign new_new_n405__ = ~new_new_n350__ & ~new_new_n353__;
  assign new_new_n406__ = G120gat & G324gat;
  assign new_new_n407__ = ~new_new_n344__ & ~new_new_n347__;
  assign new_new_n408__ = G137gat & G307gat;
  assign new_new_n409__ = G171gat & G273gat;
  assign new_new_n410__ = ~new_new_n341__ & ~new_new_n409__;
  assign new_new_n411__ = G171gat & G290gat;
  assign new_new_n412__ = new_new_n339__ & new_new_n411__;
  assign new_new_n413__ = ~new_new_n410__ & ~new_new_n412__;
  assign new_new_n414__ = ~new_new_n342__ & ~new_new_n413__;
  assign new_new_n415__ = new_new_n342__ & ~new_new_n412__;
  assign new_new_n416__ = ~new_new_n414__ & ~new_new_n415__;
  assign new_new_n417__ = ~new_new_n408__ & new_new_n416__;
  assign new_new_n418__ = new_new_n408__ & ~new_new_n416__;
  assign new_new_n419__ = ~new_new_n417__ & ~new_new_n418__;
  assign new_new_n420__ = ~new_new_n407__ & new_new_n419__;
  assign new_new_n421__ = new_new_n407__ & ~new_new_n419__;
  assign new_new_n422__ = ~new_new_n420__ & ~new_new_n421__;
  assign new_new_n423__ = ~new_new_n406__ & new_new_n422__;
  assign new_new_n424__ = new_new_n406__ & ~new_new_n422__;
  assign new_new_n425__ = ~new_new_n423__ & ~new_new_n424__;
  assign new_new_n426__ = ~new_new_n405__ & new_new_n425__;
  assign new_new_n427__ = new_new_n405__ & ~new_new_n425__;
  assign new_new_n428__ = ~new_new_n426__ & ~new_new_n427__;
  assign new_new_n429__ = ~new_new_n404__ & new_new_n428__;
  assign new_new_n430__ = new_new_n404__ & ~new_new_n428__;
  assign new_new_n431__ = ~new_new_n429__ & ~new_new_n430__;
  assign new_new_n432__ = ~new_new_n403__ & new_new_n431__;
  assign new_new_n433__ = new_new_n403__ & ~new_new_n431__;
  assign new_new_n434__ = ~new_new_n432__ & ~new_new_n433__;
  assign new_new_n435__ = ~new_new_n402__ & new_new_n434__;
  assign new_new_n436__ = new_new_n402__ & ~new_new_n434__;
  assign new_new_n437__ = ~new_new_n435__ & ~new_new_n436__;
  assign new_new_n438__ = ~new_new_n401__ & new_new_n437__;
  assign new_new_n439__ = new_new_n401__ & ~new_new_n437__;
  assign new_new_n440__ = ~new_new_n438__ & ~new_new_n439__;
  assign new_new_n441__ = ~new_new_n400__ & new_new_n440__;
  assign new_new_n442__ = new_new_n400__ & ~new_new_n440__;
  assign new_new_n443__ = ~new_new_n441__ & ~new_new_n442__;
  assign new_new_n444__ = ~new_new_n399__ & new_new_n443__;
  assign new_new_n445__ = new_new_n399__ & ~new_new_n443__;
  assign new_new_n446__ = ~new_new_n444__ & ~new_new_n445__;
  assign new_new_n447__ = ~new_new_n398__ & new_new_n446__;
  assign new_new_n448__ = new_new_n398__ & ~new_new_n446__;
  assign new_new_n449__ = ~new_new_n447__ & ~new_new_n448__;
  assign new_new_n450__ = ~new_new_n397__ & new_new_n449__;
  assign new_new_n451__ = new_new_n397__ & ~new_new_n449__;
  assign new_new_n452__ = ~new_new_n450__ & ~new_new_n451__;
  assign new_new_n453__ = ~new_new_n396__ & new_new_n452__;
  assign new_new_n454__ = new_new_n396__ & ~new_new_n452__;
  assign new_new_n455__ = ~new_new_n453__ & ~new_new_n454__;
  assign new_new_n456__ = ~new_new_n395__ & new_new_n455__;
  assign new_new_n457__ = new_new_n395__ & ~new_new_n455__;
  assign new_new_n458__ = ~new_new_n456__ & ~new_new_n457__;
  assign new_new_n459__ = ~new_new_n394__ & new_new_n458__;
  assign new_new_n460__ = new_new_n394__ & ~new_new_n458__;
  assign new_new_n461__ = ~new_new_n459__ & ~new_new_n460__;
  assign new_new_n462__ = ~new_new_n393__ & new_new_n461__;
  assign new_new_n463__ = new_new_n393__ & ~new_new_n461__;
  assign new_new_n464__ = ~new_new_n462__ & ~new_new_n463__;
  assign new_new_n465__ = ~new_new_n392__ & new_new_n464__;
  assign new_new_n466__ = new_new_n392__ & ~new_new_n464__;
  assign G4591gat = new_new_n465__ | new_new_n466__;
  assign new_new_n468__ = G1gat & G460gat;
  assign new_new_n469__ = ~new_new_n462__ & ~new_new_n465__;
  assign new_new_n470__ = G18gat & G443gat;
  assign new_new_n471__ = ~new_new_n456__ & ~new_new_n459__;
  assign new_new_n472__ = G35gat & G426gat;
  assign new_new_n473__ = ~new_new_n450__ & ~new_new_n453__;
  assign new_new_n474__ = G52gat & G409gat;
  assign new_new_n475__ = ~new_new_n444__ & ~new_new_n447__;
  assign new_new_n476__ = G69gat & G392gat;
  assign new_new_n477__ = ~new_new_n438__ & ~new_new_n441__;
  assign new_new_n478__ = G86gat & G375gat;
  assign new_new_n479__ = ~new_new_n432__ & ~new_new_n435__;
  assign new_new_n480__ = G103gat & G358gat;
  assign new_new_n481__ = ~new_new_n426__ & ~new_new_n429__;
  assign new_new_n482__ = G120gat & G341gat;
  assign new_new_n483__ = ~new_new_n420__ & ~new_new_n423__;
  assign new_new_n484__ = G137gat & G324gat;
  assign new_new_n485__ = ~new_new_n414__ & ~new_new_n417__;
  assign new_new_n486__ = G154gat & G307gat;
  assign new_new_n487__ = G188gat & G273gat;
  assign new_new_n488__ = ~new_new_n411__ & ~new_new_n487__;
  assign new_new_n489__ = G188gat & G290gat;
  assign new_new_n490__ = new_new_n409__ & new_new_n489__;
  assign new_new_n491__ = ~new_new_n488__ & ~new_new_n490__;
  assign new_new_n492__ = ~new_new_n412__ & ~new_new_n491__;
  assign new_new_n493__ = new_new_n412__ & ~new_new_n490__;
  assign new_new_n494__ = ~new_new_n492__ & ~new_new_n493__;
  assign new_new_n495__ = ~new_new_n486__ & new_new_n494__;
  assign new_new_n496__ = new_new_n486__ & ~new_new_n494__;
  assign new_new_n497__ = ~new_new_n495__ & ~new_new_n496__;
  assign new_new_n498__ = ~new_new_n485__ & new_new_n497__;
  assign new_new_n499__ = new_new_n485__ & ~new_new_n497__;
  assign new_new_n500__ = ~new_new_n498__ & ~new_new_n499__;
  assign new_new_n501__ = ~new_new_n484__ & new_new_n500__;
  assign new_new_n502__ = new_new_n484__ & ~new_new_n500__;
  assign new_new_n503__ = ~new_new_n501__ & ~new_new_n502__;
  assign new_new_n504__ = ~new_new_n483__ & new_new_n503__;
  assign new_new_n505__ = new_new_n483__ & ~new_new_n503__;
  assign new_new_n506__ = ~new_new_n504__ & ~new_new_n505__;
  assign new_new_n507__ = ~new_new_n482__ & new_new_n506__;
  assign new_new_n508__ = new_new_n482__ & ~new_new_n506__;
  assign new_new_n509__ = ~new_new_n507__ & ~new_new_n508__;
  assign new_new_n510__ = ~new_new_n481__ & new_new_n509__;
  assign new_new_n511__ = new_new_n481__ & ~new_new_n509__;
  assign new_new_n512__ = ~new_new_n510__ & ~new_new_n511__;
  assign new_new_n513__ = ~new_new_n480__ & new_new_n512__;
  assign new_new_n514__ = new_new_n480__ & ~new_new_n512__;
  assign new_new_n515__ = ~new_new_n513__ & ~new_new_n514__;
  assign new_new_n516__ = ~new_new_n479__ & new_new_n515__;
  assign new_new_n517__ = new_new_n479__ & ~new_new_n515__;
  assign new_new_n518__ = ~new_new_n516__ & ~new_new_n517__;
  assign new_new_n519__ = ~new_new_n478__ & new_new_n518__;
  assign new_new_n520__ = new_new_n478__ & ~new_new_n518__;
  assign new_new_n521__ = ~new_new_n519__ & ~new_new_n520__;
  assign new_new_n522__ = ~new_new_n477__ & new_new_n521__;
  assign new_new_n523__ = new_new_n477__ & ~new_new_n521__;
  assign new_new_n524__ = ~new_new_n522__ & ~new_new_n523__;
  assign new_new_n525__ = ~new_new_n476__ & new_new_n524__;
  assign new_new_n526__ = new_new_n476__ & ~new_new_n524__;
  assign new_new_n527__ = ~new_new_n525__ & ~new_new_n526__;
  assign new_new_n528__ = ~new_new_n475__ & new_new_n527__;
  assign new_new_n529__ = new_new_n475__ & ~new_new_n527__;
  assign new_new_n530__ = ~new_new_n528__ & ~new_new_n529__;
  assign new_new_n531__ = ~new_new_n474__ & new_new_n530__;
  assign new_new_n532__ = new_new_n474__ & ~new_new_n530__;
  assign new_new_n533__ = ~new_new_n531__ & ~new_new_n532__;
  assign new_new_n534__ = ~new_new_n473__ & new_new_n533__;
  assign new_new_n535__ = new_new_n473__ & ~new_new_n533__;
  assign new_new_n536__ = ~new_new_n534__ & ~new_new_n535__;
  assign new_new_n537__ = ~new_new_n472__ & new_new_n536__;
  assign new_new_n538__ = new_new_n472__ & ~new_new_n536__;
  assign new_new_n539__ = ~new_new_n537__ & ~new_new_n538__;
  assign new_new_n540__ = ~new_new_n471__ & new_new_n539__;
  assign new_new_n541__ = new_new_n471__ & ~new_new_n539__;
  assign new_new_n542__ = ~new_new_n540__ & ~new_new_n541__;
  assign new_new_n543__ = ~new_new_n470__ & new_new_n542__;
  assign new_new_n544__ = new_new_n470__ & ~new_new_n542__;
  assign new_new_n545__ = ~new_new_n543__ & ~new_new_n544__;
  assign new_new_n546__ = ~new_new_n469__ & new_new_n545__;
  assign new_new_n547__ = new_new_n469__ & ~new_new_n545__;
  assign new_new_n548__ = ~new_new_n546__ & ~new_new_n547__;
  assign new_new_n549__ = ~new_new_n468__ & new_new_n548__;
  assign new_new_n550__ = new_new_n468__ & ~new_new_n548__;
  assign G4946gat = new_new_n549__ | new_new_n550__;
  assign new_new_n552__ = G1gat & G477gat;
  assign new_new_n553__ = ~new_new_n546__ & ~new_new_n549__;
  assign new_new_n554__ = G18gat & G460gat;
  assign new_new_n555__ = ~new_new_n540__ & ~new_new_n543__;
  assign new_new_n556__ = G35gat & G443gat;
  assign new_new_n557__ = ~new_new_n534__ & ~new_new_n537__;
  assign new_new_n558__ = G52gat & G426gat;
  assign new_new_n559__ = ~new_new_n528__ & ~new_new_n531__;
  assign new_new_n560__ = G69gat & G409gat;
  assign new_new_n561__ = ~new_new_n522__ & ~new_new_n525__;
  assign new_new_n562__ = G86gat & G392gat;
  assign new_new_n563__ = ~new_new_n516__ & ~new_new_n519__;
  assign new_new_n564__ = G103gat & G375gat;
  assign new_new_n565__ = ~new_new_n510__ & ~new_new_n513__;
  assign new_new_n566__ = G120gat & G358gat;
  assign new_new_n567__ = ~new_new_n504__ & ~new_new_n507__;
  assign new_new_n568__ = G137gat & G341gat;
  assign new_new_n569__ = ~new_new_n498__ & ~new_new_n501__;
  assign new_new_n570__ = G154gat & G324gat;
  assign new_new_n571__ = ~new_new_n492__ & ~new_new_n495__;
  assign new_new_n572__ = G171gat & G307gat;
  assign new_new_n573__ = G205gat & G273gat;
  assign new_new_n574__ = ~new_new_n489__ & ~new_new_n573__;
  assign new_new_n575__ = G205gat & G290gat;
  assign new_new_n576__ = new_new_n487__ & new_new_n575__;
  assign new_new_n577__ = ~new_new_n574__ & ~new_new_n576__;
  assign new_new_n578__ = ~new_new_n490__ & ~new_new_n577__;
  assign new_new_n579__ = new_new_n490__ & ~new_new_n576__;
  assign new_new_n580__ = ~new_new_n578__ & ~new_new_n579__;
  assign new_new_n581__ = ~new_new_n572__ & new_new_n580__;
  assign new_new_n582__ = new_new_n572__ & ~new_new_n580__;
  assign new_new_n583__ = ~new_new_n581__ & ~new_new_n582__;
  assign new_new_n584__ = ~new_new_n571__ & new_new_n583__;
  assign new_new_n585__ = new_new_n571__ & ~new_new_n583__;
  assign new_new_n586__ = ~new_new_n584__ & ~new_new_n585__;
  assign new_new_n587__ = ~new_new_n570__ & new_new_n586__;
  assign new_new_n588__ = new_new_n570__ & ~new_new_n586__;
  assign new_new_n589__ = ~new_new_n587__ & ~new_new_n588__;
  assign new_new_n590__ = ~new_new_n569__ & new_new_n589__;
  assign new_new_n591__ = new_new_n569__ & ~new_new_n589__;
  assign new_new_n592__ = ~new_new_n590__ & ~new_new_n591__;
  assign new_new_n593__ = ~new_new_n568__ & new_new_n592__;
  assign new_new_n594__ = new_new_n568__ & ~new_new_n592__;
  assign new_new_n595__ = ~new_new_n593__ & ~new_new_n594__;
  assign new_new_n596__ = ~new_new_n567__ & new_new_n595__;
  assign new_new_n597__ = new_new_n567__ & ~new_new_n595__;
  assign new_new_n598__ = ~new_new_n596__ & ~new_new_n597__;
  assign new_new_n599__ = ~new_new_n566__ & new_new_n598__;
  assign new_new_n600__ = new_new_n566__ & ~new_new_n598__;
  assign new_new_n601__ = ~new_new_n599__ & ~new_new_n600__;
  assign new_new_n602__ = ~new_new_n565__ & new_new_n601__;
  assign new_new_n603__ = new_new_n565__ & ~new_new_n601__;
  assign new_new_n604__ = ~new_new_n602__ & ~new_new_n603__;
  assign new_new_n605__ = ~new_new_n564__ & new_new_n604__;
  assign new_new_n606__ = new_new_n564__ & ~new_new_n604__;
  assign new_new_n607__ = ~new_new_n605__ & ~new_new_n606__;
  assign new_new_n608__ = ~new_new_n563__ & new_new_n607__;
  assign new_new_n609__ = new_new_n563__ & ~new_new_n607__;
  assign new_new_n610__ = ~new_new_n608__ & ~new_new_n609__;
  assign new_new_n611__ = ~new_new_n562__ & new_new_n610__;
  assign new_new_n612__ = new_new_n562__ & ~new_new_n610__;
  assign new_new_n613__ = ~new_new_n611__ & ~new_new_n612__;
  assign new_new_n614__ = ~new_new_n561__ & new_new_n613__;
  assign new_new_n615__ = new_new_n561__ & ~new_new_n613__;
  assign new_new_n616__ = ~new_new_n614__ & ~new_new_n615__;
  assign new_new_n617__ = ~new_new_n560__ & new_new_n616__;
  assign new_new_n618__ = new_new_n560__ & ~new_new_n616__;
  assign new_new_n619__ = ~new_new_n617__ & ~new_new_n618__;
  assign new_new_n620__ = ~new_new_n559__ & new_new_n619__;
  assign new_new_n621__ = new_new_n559__ & ~new_new_n619__;
  assign new_new_n622__ = ~new_new_n620__ & ~new_new_n621__;
  assign new_new_n623__ = ~new_new_n558__ & new_new_n622__;
  assign new_new_n624__ = new_new_n558__ & ~new_new_n622__;
  assign new_new_n625__ = ~new_new_n623__ & ~new_new_n624__;
  assign new_new_n626__ = ~new_new_n557__ & new_new_n625__;
  assign new_new_n627__ = new_new_n557__ & ~new_new_n625__;
  assign new_new_n628__ = ~new_new_n626__ & ~new_new_n627__;
  assign new_new_n629__ = ~new_new_n556__ & new_new_n628__;
  assign new_new_n630__ = new_new_n556__ & ~new_new_n628__;
  assign new_new_n631__ = ~new_new_n629__ & ~new_new_n630__;
  assign new_new_n632__ = ~new_new_n555__ & new_new_n631__;
  assign new_new_n633__ = new_new_n555__ & ~new_new_n631__;
  assign new_new_n634__ = ~new_new_n632__ & ~new_new_n633__;
  assign new_new_n635__ = ~new_new_n554__ & new_new_n634__;
  assign new_new_n636__ = new_new_n554__ & ~new_new_n634__;
  assign new_new_n637__ = ~new_new_n635__ & ~new_new_n636__;
  assign new_new_n638__ = ~new_new_n553__ & new_new_n637__;
  assign new_new_n639__ = new_new_n553__ & ~new_new_n637__;
  assign new_new_n640__ = ~new_new_n638__ & ~new_new_n639__;
  assign new_new_n641__ = ~new_new_n552__ & new_new_n640__;
  assign new_new_n642__ = new_new_n552__ & ~new_new_n640__;
  assign G5308gat = new_new_n641__ | new_new_n642__;
  assign new_new_n644__ = G1gat & G494gat;
  assign new_new_n645__ = ~new_new_n638__ & ~new_new_n641__;
  assign new_new_n646__ = G18gat & G477gat;
  assign new_new_n647__ = ~new_new_n632__ & ~new_new_n635__;
  assign new_new_n648__ = G35gat & G460gat;
  assign new_new_n649__ = ~new_new_n626__ & ~new_new_n629__;
  assign new_new_n650__ = G52gat & G443gat;
  assign new_new_n651__ = ~new_new_n620__ & ~new_new_n623__;
  assign new_new_n652__ = G69gat & G426gat;
  assign new_new_n653__ = ~new_new_n614__ & ~new_new_n617__;
  assign new_new_n654__ = G86gat & G409gat;
  assign new_new_n655__ = ~new_new_n608__ & ~new_new_n611__;
  assign new_new_n656__ = G103gat & G392gat;
  assign new_new_n657__ = ~new_new_n602__ & ~new_new_n605__;
  assign new_new_n658__ = G120gat & G375gat;
  assign new_new_n659__ = ~new_new_n596__ & ~new_new_n599__;
  assign new_new_n660__ = G137gat & G358gat;
  assign new_new_n661__ = ~new_new_n590__ & ~new_new_n593__;
  assign new_new_n662__ = G154gat & G341gat;
  assign new_new_n663__ = ~new_new_n584__ & ~new_new_n587__;
  assign new_new_n664__ = G171gat & G324gat;
  assign new_new_n665__ = ~new_new_n578__ & ~new_new_n581__;
  assign new_new_n666__ = G188gat & G307gat;
  assign new_new_n667__ = G222gat & G273gat;
  assign new_new_n668__ = ~new_new_n575__ & ~new_new_n667__;
  assign new_new_n669__ = G222gat & G290gat;
  assign new_new_n670__ = new_new_n573__ & new_new_n669__;
  assign new_new_n671__ = ~new_new_n668__ & ~new_new_n670__;
  assign new_new_n672__ = ~new_new_n576__ & ~new_new_n671__;
  assign new_new_n673__ = new_new_n576__ & ~new_new_n670__;
  assign new_new_n674__ = ~new_new_n672__ & ~new_new_n673__;
  assign new_new_n675__ = ~new_new_n666__ & new_new_n674__;
  assign new_new_n676__ = new_new_n666__ & ~new_new_n674__;
  assign new_new_n677__ = ~new_new_n675__ & ~new_new_n676__;
  assign new_new_n678__ = ~new_new_n665__ & new_new_n677__;
  assign new_new_n679__ = new_new_n665__ & ~new_new_n677__;
  assign new_new_n680__ = ~new_new_n678__ & ~new_new_n679__;
  assign new_new_n681__ = ~new_new_n664__ & new_new_n680__;
  assign new_new_n682__ = new_new_n664__ & ~new_new_n680__;
  assign new_new_n683__ = ~new_new_n681__ & ~new_new_n682__;
  assign new_new_n684__ = ~new_new_n663__ & new_new_n683__;
  assign new_new_n685__ = new_new_n663__ & ~new_new_n683__;
  assign new_new_n686__ = ~new_new_n684__ & ~new_new_n685__;
  assign new_new_n687__ = ~new_new_n662__ & new_new_n686__;
  assign new_new_n688__ = new_new_n662__ & ~new_new_n686__;
  assign new_new_n689__ = ~new_new_n687__ & ~new_new_n688__;
  assign new_new_n690__ = ~new_new_n661__ & new_new_n689__;
  assign new_new_n691__ = new_new_n661__ & ~new_new_n689__;
  assign new_new_n692__ = ~new_new_n690__ & ~new_new_n691__;
  assign new_new_n693__ = ~new_new_n660__ & new_new_n692__;
  assign new_new_n694__ = new_new_n660__ & ~new_new_n692__;
  assign new_new_n695__ = ~new_new_n693__ & ~new_new_n694__;
  assign new_new_n696__ = ~new_new_n659__ & new_new_n695__;
  assign new_new_n697__ = new_new_n659__ & ~new_new_n695__;
  assign new_new_n698__ = ~new_new_n696__ & ~new_new_n697__;
  assign new_new_n699__ = ~new_new_n658__ & new_new_n698__;
  assign new_new_n700__ = new_new_n658__ & ~new_new_n698__;
  assign new_new_n701__ = ~new_new_n699__ & ~new_new_n700__;
  assign new_new_n702__ = ~new_new_n657__ & new_new_n701__;
  assign new_new_n703__ = new_new_n657__ & ~new_new_n701__;
  assign new_new_n704__ = ~new_new_n702__ & ~new_new_n703__;
  assign new_new_n705__ = ~new_new_n656__ & new_new_n704__;
  assign new_new_n706__ = new_new_n656__ & ~new_new_n704__;
  assign new_new_n707__ = ~new_new_n705__ & ~new_new_n706__;
  assign new_new_n708__ = ~new_new_n655__ & new_new_n707__;
  assign new_new_n709__ = new_new_n655__ & ~new_new_n707__;
  assign new_new_n710__ = ~new_new_n708__ & ~new_new_n709__;
  assign new_new_n711__ = ~new_new_n654__ & new_new_n710__;
  assign new_new_n712__ = new_new_n654__ & ~new_new_n710__;
  assign new_new_n713__ = ~new_new_n711__ & ~new_new_n712__;
  assign new_new_n714__ = ~new_new_n653__ & new_new_n713__;
  assign new_new_n715__ = new_new_n653__ & ~new_new_n713__;
  assign new_new_n716__ = ~new_new_n714__ & ~new_new_n715__;
  assign new_new_n717__ = ~new_new_n652__ & new_new_n716__;
  assign new_new_n718__ = new_new_n652__ & ~new_new_n716__;
  assign new_new_n719__ = ~new_new_n717__ & ~new_new_n718__;
  assign new_new_n720__ = ~new_new_n651__ & new_new_n719__;
  assign new_new_n721__ = new_new_n651__ & ~new_new_n719__;
  assign new_new_n722__ = ~new_new_n720__ & ~new_new_n721__;
  assign new_new_n723__ = ~new_new_n650__ & new_new_n722__;
  assign new_new_n724__ = new_new_n650__ & ~new_new_n722__;
  assign new_new_n725__ = ~new_new_n723__ & ~new_new_n724__;
  assign new_new_n726__ = ~new_new_n649__ & new_new_n725__;
  assign new_new_n727__ = new_new_n649__ & ~new_new_n725__;
  assign new_new_n728__ = ~new_new_n726__ & ~new_new_n727__;
  assign new_new_n729__ = ~new_new_n648__ & new_new_n728__;
  assign new_new_n730__ = new_new_n648__ & ~new_new_n728__;
  assign new_new_n731__ = ~new_new_n729__ & ~new_new_n730__;
  assign new_new_n732__ = ~new_new_n647__ & new_new_n731__;
  assign new_new_n733__ = new_new_n647__ & ~new_new_n731__;
  assign new_new_n734__ = ~new_new_n732__ & ~new_new_n733__;
  assign new_new_n735__ = ~new_new_n646__ & new_new_n734__;
  assign new_new_n736__ = new_new_n646__ & ~new_new_n734__;
  assign new_new_n737__ = ~new_new_n735__ & ~new_new_n736__;
  assign new_new_n738__ = ~new_new_n645__ & new_new_n737__;
  assign new_new_n739__ = new_new_n645__ & ~new_new_n737__;
  assign new_new_n740__ = ~new_new_n738__ & ~new_new_n739__;
  assign new_new_n741__ = ~new_new_n644__ & new_new_n740__;
  assign new_new_n742__ = new_new_n644__ & ~new_new_n740__;
  assign G5672gat = new_new_n741__ | new_new_n742__;
  assign new_new_n744__ = G1gat & G511gat;
  assign new_new_n745__ = ~new_new_n738__ & ~new_new_n741__;
  assign new_new_n746__ = G18gat & G494gat;
  assign new_new_n747__ = ~new_new_n732__ & ~new_new_n735__;
  assign new_new_n748__ = G35gat & G477gat;
  assign new_new_n749__ = ~new_new_n726__ & ~new_new_n729__;
  assign new_new_n750__ = G52gat & G460gat;
  assign new_new_n751__ = ~new_new_n720__ & ~new_new_n723__;
  assign new_new_n752__ = G69gat & G443gat;
  assign new_new_n753__ = ~new_new_n714__ & ~new_new_n717__;
  assign new_new_n754__ = G86gat & G426gat;
  assign new_new_n755__ = ~new_new_n708__ & ~new_new_n711__;
  assign new_new_n756__ = G103gat & G409gat;
  assign new_new_n757__ = ~new_new_n702__ & ~new_new_n705__;
  assign new_new_n758__ = G120gat & G392gat;
  assign new_new_n759__ = ~new_new_n696__ & ~new_new_n699__;
  assign new_new_n760__ = G137gat & G375gat;
  assign new_new_n761__ = ~new_new_n690__ & ~new_new_n693__;
  assign new_new_n762__ = G154gat & G358gat;
  assign new_new_n763__ = ~new_new_n684__ & ~new_new_n687__;
  assign new_new_n764__ = G171gat & G341gat;
  assign new_new_n765__ = ~new_new_n678__ & ~new_new_n681__;
  assign new_new_n766__ = G188gat & G324gat;
  assign new_new_n767__ = ~new_new_n672__ & ~new_new_n675__;
  assign new_new_n768__ = G205gat & G307gat;
  assign new_new_n769__ = G239gat & G273gat;
  assign new_new_n770__ = ~new_new_n669__ & ~new_new_n769__;
  assign new_new_n771__ = G239gat & G290gat;
  assign new_new_n772__ = new_new_n667__ & new_new_n771__;
  assign new_new_n773__ = ~new_new_n770__ & ~new_new_n772__;
  assign new_new_n774__ = ~new_new_n670__ & ~new_new_n773__;
  assign new_new_n775__ = new_new_n670__ & ~new_new_n772__;
  assign new_new_n776__ = ~new_new_n774__ & ~new_new_n775__;
  assign new_new_n777__ = ~new_new_n768__ & new_new_n776__;
  assign new_new_n778__ = new_new_n768__ & ~new_new_n776__;
  assign new_new_n779__ = ~new_new_n777__ & ~new_new_n778__;
  assign new_new_n780__ = ~new_new_n767__ & new_new_n779__;
  assign new_new_n781__ = new_new_n767__ & ~new_new_n779__;
  assign new_new_n782__ = ~new_new_n780__ & ~new_new_n781__;
  assign new_new_n783__ = ~new_new_n766__ & new_new_n782__;
  assign new_new_n784__ = new_new_n766__ & ~new_new_n782__;
  assign new_new_n785__ = ~new_new_n783__ & ~new_new_n784__;
  assign new_new_n786__ = ~new_new_n765__ & new_new_n785__;
  assign new_new_n787__ = new_new_n765__ & ~new_new_n785__;
  assign new_new_n788__ = ~new_new_n786__ & ~new_new_n787__;
  assign new_new_n789__ = ~new_new_n764__ & new_new_n788__;
  assign new_new_n790__ = new_new_n764__ & ~new_new_n788__;
  assign new_new_n791__ = ~new_new_n789__ & ~new_new_n790__;
  assign new_new_n792__ = ~new_new_n763__ & new_new_n791__;
  assign new_new_n793__ = new_new_n763__ & ~new_new_n791__;
  assign new_new_n794__ = ~new_new_n792__ & ~new_new_n793__;
  assign new_new_n795__ = ~new_new_n762__ & new_new_n794__;
  assign new_new_n796__ = new_new_n762__ & ~new_new_n794__;
  assign new_new_n797__ = ~new_new_n795__ & ~new_new_n796__;
  assign new_new_n798__ = ~new_new_n761__ & new_new_n797__;
  assign new_new_n799__ = new_new_n761__ & ~new_new_n797__;
  assign new_new_n800__ = ~new_new_n798__ & ~new_new_n799__;
  assign new_new_n801__ = ~new_new_n760__ & new_new_n800__;
  assign new_new_n802__ = new_new_n760__ & ~new_new_n800__;
  assign new_new_n803__ = ~new_new_n801__ & ~new_new_n802__;
  assign new_new_n804__ = ~new_new_n759__ & new_new_n803__;
  assign new_new_n805__ = new_new_n759__ & ~new_new_n803__;
  assign new_new_n806__ = ~new_new_n804__ & ~new_new_n805__;
  assign new_new_n807__ = ~new_new_n758__ & new_new_n806__;
  assign new_new_n808__ = new_new_n758__ & ~new_new_n806__;
  assign new_new_n809__ = ~new_new_n807__ & ~new_new_n808__;
  assign new_new_n810__ = ~new_new_n757__ & new_new_n809__;
  assign new_new_n811__ = new_new_n757__ & ~new_new_n809__;
  assign new_new_n812__ = ~new_new_n810__ & ~new_new_n811__;
  assign new_new_n813__ = ~new_new_n756__ & new_new_n812__;
  assign new_new_n814__ = new_new_n756__ & ~new_new_n812__;
  assign new_new_n815__ = ~new_new_n813__ & ~new_new_n814__;
  assign new_new_n816__ = ~new_new_n755__ & new_new_n815__;
  assign new_new_n817__ = new_new_n755__ & ~new_new_n815__;
  assign new_new_n818__ = ~new_new_n816__ & ~new_new_n817__;
  assign new_new_n819__ = ~new_new_n754__ & new_new_n818__;
  assign new_new_n820__ = new_new_n754__ & ~new_new_n818__;
  assign new_new_n821__ = ~new_new_n819__ & ~new_new_n820__;
  assign new_new_n822__ = ~new_new_n753__ & new_new_n821__;
  assign new_new_n823__ = new_new_n753__ & ~new_new_n821__;
  assign new_new_n824__ = ~new_new_n822__ & ~new_new_n823__;
  assign new_new_n825__ = ~new_new_n752__ & new_new_n824__;
  assign new_new_n826__ = new_new_n752__ & ~new_new_n824__;
  assign new_new_n827__ = ~new_new_n825__ & ~new_new_n826__;
  assign new_new_n828__ = ~new_new_n751__ & new_new_n827__;
  assign new_new_n829__ = new_new_n751__ & ~new_new_n827__;
  assign new_new_n830__ = ~new_new_n828__ & ~new_new_n829__;
  assign new_new_n831__ = ~new_new_n750__ & new_new_n830__;
  assign new_new_n832__ = new_new_n750__ & ~new_new_n830__;
  assign new_new_n833__ = ~new_new_n831__ & ~new_new_n832__;
  assign new_new_n834__ = ~new_new_n749__ & new_new_n833__;
  assign new_new_n835__ = new_new_n749__ & ~new_new_n833__;
  assign new_new_n836__ = ~new_new_n834__ & ~new_new_n835__;
  assign new_new_n837__ = ~new_new_n748__ & new_new_n836__;
  assign new_new_n838__ = new_new_n748__ & ~new_new_n836__;
  assign new_new_n839__ = ~new_new_n837__ & ~new_new_n838__;
  assign new_new_n840__ = ~new_new_n747__ & new_new_n839__;
  assign new_new_n841__ = new_new_n747__ & ~new_new_n839__;
  assign new_new_n842__ = ~new_new_n840__ & ~new_new_n841__;
  assign new_new_n843__ = ~new_new_n746__ & new_new_n842__;
  assign new_new_n844__ = new_new_n746__ & ~new_new_n842__;
  assign new_new_n845__ = ~new_new_n843__ & ~new_new_n844__;
  assign new_new_n846__ = ~new_new_n745__ & new_new_n845__;
  assign new_new_n847__ = new_new_n745__ & ~new_new_n845__;
  assign new_new_n848__ = ~new_new_n846__ & ~new_new_n847__;
  assign new_new_n849__ = ~new_new_n744__ & new_new_n848__;
  assign new_new_n850__ = new_new_n744__ & ~new_new_n848__;
  assign G5971gat = new_new_n849__ | new_new_n850__;
  assign new_new_n852__ = G1gat & G528gat;
  assign new_new_n853__ = ~new_new_n846__ & ~new_new_n849__;
  assign new_new_n854__ = G18gat & G511gat;
  assign new_new_n855__ = ~new_new_n840__ & ~new_new_n843__;
  assign new_new_n856__ = G35gat & G494gat;
  assign new_new_n857__ = ~new_new_n834__ & ~new_new_n837__;
  assign new_new_n858__ = G52gat & G477gat;
  assign new_new_n859__ = ~new_new_n828__ & ~new_new_n831__;
  assign new_new_n860__ = G69gat & G460gat;
  assign new_new_n861__ = ~new_new_n822__ & ~new_new_n825__;
  assign new_new_n862__ = G86gat & G443gat;
  assign new_new_n863__ = ~new_new_n816__ & ~new_new_n819__;
  assign new_new_n864__ = G103gat & G426gat;
  assign new_new_n865__ = ~new_new_n810__ & ~new_new_n813__;
  assign new_new_n866__ = G120gat & G409gat;
  assign new_new_n867__ = ~new_new_n804__ & ~new_new_n807__;
  assign new_new_n868__ = G137gat & G392gat;
  assign new_new_n869__ = ~new_new_n798__ & ~new_new_n801__;
  assign new_new_n870__ = G154gat & G375gat;
  assign new_new_n871__ = ~new_new_n792__ & ~new_new_n795__;
  assign new_new_n872__ = G171gat & G358gat;
  assign new_new_n873__ = ~new_new_n786__ & ~new_new_n789__;
  assign new_new_n874__ = G188gat & G341gat;
  assign new_new_n875__ = ~new_new_n780__ & ~new_new_n783__;
  assign new_new_n876__ = G205gat & G324gat;
  assign new_new_n877__ = ~new_new_n774__ & ~new_new_n777__;
  assign new_new_n878__ = G222gat & G307gat;
  assign new_new_n879__ = G256gat & G273gat;
  assign new_new_n880__ = ~new_new_n771__ & new_new_n879__;
  assign new_new_n881__ = new_new_n771__ & ~new_new_n879__;
  assign new_new_n882__ = ~new_new_n772__ & ~new_new_n880__;
  assign new_new_n883__ = ~new_new_n881__ & new_new_n882__;
  assign new_new_n884__ = new_new_n667__ & new_new_n881__;
  assign new_new_n885__ = ~new_new_n883__ & ~new_new_n884__;
  assign new_new_n886__ = ~new_new_n878__ & new_new_n885__;
  assign new_new_n887__ = new_new_n878__ & ~new_new_n885__;
  assign new_new_n888__ = ~new_new_n886__ & ~new_new_n887__;
  assign new_new_n889__ = ~new_new_n877__ & new_new_n888__;
  assign new_new_n890__ = new_new_n877__ & ~new_new_n888__;
  assign new_new_n891__ = ~new_new_n889__ & ~new_new_n890__;
  assign new_new_n892__ = ~new_new_n876__ & new_new_n891__;
  assign new_new_n893__ = new_new_n876__ & ~new_new_n891__;
  assign new_new_n894__ = ~new_new_n892__ & ~new_new_n893__;
  assign new_new_n895__ = ~new_new_n875__ & new_new_n894__;
  assign new_new_n896__ = new_new_n875__ & ~new_new_n894__;
  assign new_new_n897__ = ~new_new_n895__ & ~new_new_n896__;
  assign new_new_n898__ = ~new_new_n874__ & new_new_n897__;
  assign new_new_n899__ = new_new_n874__ & ~new_new_n897__;
  assign new_new_n900__ = ~new_new_n898__ & ~new_new_n899__;
  assign new_new_n901__ = ~new_new_n873__ & new_new_n900__;
  assign new_new_n902__ = new_new_n873__ & ~new_new_n900__;
  assign new_new_n903__ = ~new_new_n901__ & ~new_new_n902__;
  assign new_new_n904__ = ~new_new_n872__ & new_new_n903__;
  assign new_new_n905__ = new_new_n872__ & ~new_new_n903__;
  assign new_new_n906__ = ~new_new_n904__ & ~new_new_n905__;
  assign new_new_n907__ = ~new_new_n871__ & new_new_n906__;
  assign new_new_n908__ = new_new_n871__ & ~new_new_n906__;
  assign new_new_n909__ = ~new_new_n907__ & ~new_new_n908__;
  assign new_new_n910__ = ~new_new_n870__ & new_new_n909__;
  assign new_new_n911__ = new_new_n870__ & ~new_new_n909__;
  assign new_new_n912__ = ~new_new_n910__ & ~new_new_n911__;
  assign new_new_n913__ = ~new_new_n869__ & new_new_n912__;
  assign new_new_n914__ = new_new_n869__ & ~new_new_n912__;
  assign new_new_n915__ = ~new_new_n913__ & ~new_new_n914__;
  assign new_new_n916__ = ~new_new_n868__ & new_new_n915__;
  assign new_new_n917__ = new_new_n868__ & ~new_new_n915__;
  assign new_new_n918__ = ~new_new_n916__ & ~new_new_n917__;
  assign new_new_n919__ = ~new_new_n867__ & new_new_n918__;
  assign new_new_n920__ = new_new_n867__ & ~new_new_n918__;
  assign new_new_n921__ = ~new_new_n919__ & ~new_new_n920__;
  assign new_new_n922__ = ~new_new_n866__ & new_new_n921__;
  assign new_new_n923__ = new_new_n866__ & ~new_new_n921__;
  assign new_new_n924__ = ~new_new_n922__ & ~new_new_n923__;
  assign new_new_n925__ = ~new_new_n865__ & new_new_n924__;
  assign new_new_n926__ = new_new_n865__ & ~new_new_n924__;
  assign new_new_n927__ = ~new_new_n925__ & ~new_new_n926__;
  assign new_new_n928__ = ~new_new_n864__ & new_new_n927__;
  assign new_new_n929__ = new_new_n864__ & ~new_new_n927__;
  assign new_new_n930__ = ~new_new_n928__ & ~new_new_n929__;
  assign new_new_n931__ = ~new_new_n863__ & new_new_n930__;
  assign new_new_n932__ = new_new_n863__ & ~new_new_n930__;
  assign new_new_n933__ = ~new_new_n931__ & ~new_new_n932__;
  assign new_new_n934__ = ~new_new_n862__ & new_new_n933__;
  assign new_new_n935__ = new_new_n862__ & ~new_new_n933__;
  assign new_new_n936__ = ~new_new_n934__ & ~new_new_n935__;
  assign new_new_n937__ = ~new_new_n861__ & new_new_n936__;
  assign new_new_n938__ = new_new_n861__ & ~new_new_n936__;
  assign new_new_n939__ = ~new_new_n937__ & ~new_new_n938__;
  assign new_new_n940__ = ~new_new_n860__ & new_new_n939__;
  assign new_new_n941__ = new_new_n860__ & ~new_new_n939__;
  assign new_new_n942__ = ~new_new_n940__ & ~new_new_n941__;
  assign new_new_n943__ = ~new_new_n859__ & new_new_n942__;
  assign new_new_n944__ = new_new_n859__ & ~new_new_n942__;
  assign new_new_n945__ = ~new_new_n943__ & ~new_new_n944__;
  assign new_new_n946__ = ~new_new_n858__ & new_new_n945__;
  assign new_new_n947__ = new_new_n858__ & ~new_new_n945__;
  assign new_new_n948__ = ~new_new_n946__ & ~new_new_n947__;
  assign new_new_n949__ = ~new_new_n857__ & new_new_n948__;
  assign new_new_n950__ = new_new_n857__ & ~new_new_n948__;
  assign new_new_n951__ = ~new_new_n949__ & ~new_new_n950__;
  assign new_new_n952__ = ~new_new_n856__ & new_new_n951__;
  assign new_new_n953__ = new_new_n856__ & ~new_new_n951__;
  assign new_new_n954__ = ~new_new_n952__ & ~new_new_n953__;
  assign new_new_n955__ = ~new_new_n855__ & new_new_n954__;
  assign new_new_n956__ = new_new_n855__ & ~new_new_n954__;
  assign new_new_n957__ = ~new_new_n955__ & ~new_new_n956__;
  assign new_new_n958__ = ~new_new_n854__ & new_new_n957__;
  assign new_new_n959__ = new_new_n854__ & ~new_new_n957__;
  assign new_new_n960__ = ~new_new_n958__ & ~new_new_n959__;
  assign new_new_n961__ = ~new_new_n853__ & new_new_n960__;
  assign new_new_n962__ = new_new_n853__ & ~new_new_n960__;
  assign new_new_n963__ = ~new_new_n961__ & ~new_new_n962__;
  assign new_new_n964__ = ~new_new_n852__ & new_new_n963__;
  assign new_new_n965__ = new_new_n852__ & ~new_new_n963__;
  assign G6123gat = new_new_n964__ | new_new_n965__;
  assign new_new_n967__ = ~new_new_n961__ & ~new_new_n964__;
  assign new_new_n968__ = G18gat & G528gat;
  assign new_new_n969__ = ~new_new_n955__ & ~new_new_n958__;
  assign new_new_n970__ = G35gat & G511gat;
  assign new_new_n971__ = ~new_new_n949__ & ~new_new_n952__;
  assign new_new_n972__ = G52gat & G494gat;
  assign new_new_n973__ = ~new_new_n943__ & ~new_new_n946__;
  assign new_new_n974__ = G69gat & G477gat;
  assign new_new_n975__ = ~new_new_n937__ & ~new_new_n940__;
  assign new_new_n976__ = G86gat & G460gat;
  assign new_new_n977__ = ~new_new_n931__ & ~new_new_n934__;
  assign new_new_n978__ = G103gat & G443gat;
  assign new_new_n979__ = ~new_new_n925__ & ~new_new_n928__;
  assign new_new_n980__ = G120gat & G426gat;
  assign new_new_n981__ = ~new_new_n919__ & ~new_new_n922__;
  assign new_new_n982__ = G137gat & G409gat;
  assign new_new_n983__ = ~new_new_n913__ & ~new_new_n916__;
  assign new_new_n984__ = G154gat & G392gat;
  assign new_new_n985__ = ~new_new_n907__ & ~new_new_n910__;
  assign new_new_n986__ = G171gat & G375gat;
  assign new_new_n987__ = ~new_new_n901__ & ~new_new_n904__;
  assign new_new_n988__ = G188gat & G358gat;
  assign new_new_n989__ = ~new_new_n895__ & ~new_new_n898__;
  assign new_new_n990__ = G205gat & G341gat;
  assign new_new_n991__ = ~new_new_n889__ & ~new_new_n892__;
  assign new_new_n992__ = G222gat & G324gat;
  assign new_new_n993__ = ~new_new_n883__ & ~new_new_n886__;
  assign new_new_n994__ = G239gat & G307gat;
  assign new_new_n995__ = G256gat & G290gat;
  assign new_new_n996__ = ~new_new_n769__ & new_new_n995__;
  assign new_new_n997__ = ~new_new_n994__ & new_new_n996__;
  assign new_new_n998__ = new_new_n994__ & ~new_new_n996__;
  assign new_new_n999__ = ~new_new_n997__ & ~new_new_n998__;
  assign new_new_n1000__ = ~new_new_n993__ & new_new_n999__;
  assign new_new_n1001__ = new_new_n993__ & ~new_new_n999__;
  assign new_new_n1002__ = ~new_new_n1000__ & ~new_new_n1001__;
  assign new_new_n1003__ = ~new_new_n992__ & new_new_n1002__;
  assign new_new_n1004__ = new_new_n992__ & ~new_new_n1002__;
  assign new_new_n1005__ = ~new_new_n1003__ & ~new_new_n1004__;
  assign new_new_n1006__ = ~new_new_n991__ & new_new_n1005__;
  assign new_new_n1007__ = new_new_n991__ & ~new_new_n1005__;
  assign new_new_n1008__ = ~new_new_n1006__ & ~new_new_n1007__;
  assign new_new_n1009__ = ~new_new_n990__ & new_new_n1008__;
  assign new_new_n1010__ = new_new_n990__ & ~new_new_n1008__;
  assign new_new_n1011__ = ~new_new_n1009__ & ~new_new_n1010__;
  assign new_new_n1012__ = ~new_new_n989__ & new_new_n1011__;
  assign new_new_n1013__ = new_new_n989__ & ~new_new_n1011__;
  assign new_new_n1014__ = ~new_new_n1012__ & ~new_new_n1013__;
  assign new_new_n1015__ = ~new_new_n988__ & new_new_n1014__;
  assign new_new_n1016__ = new_new_n988__ & ~new_new_n1014__;
  assign new_new_n1017__ = ~new_new_n1015__ & ~new_new_n1016__;
  assign new_new_n1018__ = ~new_new_n987__ & new_new_n1017__;
  assign new_new_n1019__ = new_new_n987__ & ~new_new_n1017__;
  assign new_new_n1020__ = ~new_new_n1018__ & ~new_new_n1019__;
  assign new_new_n1021__ = ~new_new_n986__ & new_new_n1020__;
  assign new_new_n1022__ = new_new_n986__ & ~new_new_n1020__;
  assign new_new_n1023__ = ~new_new_n1021__ & ~new_new_n1022__;
  assign new_new_n1024__ = ~new_new_n985__ & new_new_n1023__;
  assign new_new_n1025__ = new_new_n985__ & ~new_new_n1023__;
  assign new_new_n1026__ = ~new_new_n1024__ & ~new_new_n1025__;
  assign new_new_n1027__ = ~new_new_n984__ & new_new_n1026__;
  assign new_new_n1028__ = new_new_n984__ & ~new_new_n1026__;
  assign new_new_n1029__ = ~new_new_n1027__ & ~new_new_n1028__;
  assign new_new_n1030__ = ~new_new_n983__ & new_new_n1029__;
  assign new_new_n1031__ = new_new_n983__ & ~new_new_n1029__;
  assign new_new_n1032__ = ~new_new_n1030__ & ~new_new_n1031__;
  assign new_new_n1033__ = ~new_new_n982__ & new_new_n1032__;
  assign new_new_n1034__ = new_new_n982__ & ~new_new_n1032__;
  assign new_new_n1035__ = ~new_new_n1033__ & ~new_new_n1034__;
  assign new_new_n1036__ = ~new_new_n981__ & new_new_n1035__;
  assign new_new_n1037__ = new_new_n981__ & ~new_new_n1035__;
  assign new_new_n1038__ = ~new_new_n1036__ & ~new_new_n1037__;
  assign new_new_n1039__ = ~new_new_n980__ & new_new_n1038__;
  assign new_new_n1040__ = new_new_n980__ & ~new_new_n1038__;
  assign new_new_n1041__ = ~new_new_n1039__ & ~new_new_n1040__;
  assign new_new_n1042__ = ~new_new_n979__ & new_new_n1041__;
  assign new_new_n1043__ = new_new_n979__ & ~new_new_n1041__;
  assign new_new_n1044__ = ~new_new_n1042__ & ~new_new_n1043__;
  assign new_new_n1045__ = ~new_new_n978__ & new_new_n1044__;
  assign new_new_n1046__ = new_new_n978__ & ~new_new_n1044__;
  assign new_new_n1047__ = ~new_new_n1045__ & ~new_new_n1046__;
  assign new_new_n1048__ = ~new_new_n977__ & new_new_n1047__;
  assign new_new_n1049__ = new_new_n977__ & ~new_new_n1047__;
  assign new_new_n1050__ = ~new_new_n1048__ & ~new_new_n1049__;
  assign new_new_n1051__ = ~new_new_n976__ & new_new_n1050__;
  assign new_new_n1052__ = new_new_n976__ & ~new_new_n1050__;
  assign new_new_n1053__ = ~new_new_n1051__ & ~new_new_n1052__;
  assign new_new_n1054__ = ~new_new_n975__ & new_new_n1053__;
  assign new_new_n1055__ = new_new_n975__ & ~new_new_n1053__;
  assign new_new_n1056__ = ~new_new_n1054__ & ~new_new_n1055__;
  assign new_new_n1057__ = ~new_new_n974__ & new_new_n1056__;
  assign new_new_n1058__ = new_new_n974__ & ~new_new_n1056__;
  assign new_new_n1059__ = ~new_new_n1057__ & ~new_new_n1058__;
  assign new_new_n1060__ = ~new_new_n973__ & new_new_n1059__;
  assign new_new_n1061__ = new_new_n973__ & ~new_new_n1059__;
  assign new_new_n1062__ = ~new_new_n1060__ & ~new_new_n1061__;
  assign new_new_n1063__ = ~new_new_n972__ & new_new_n1062__;
  assign new_new_n1064__ = new_new_n972__ & ~new_new_n1062__;
  assign new_new_n1065__ = ~new_new_n1063__ & ~new_new_n1064__;
  assign new_new_n1066__ = ~new_new_n971__ & new_new_n1065__;
  assign new_new_n1067__ = new_new_n971__ & ~new_new_n1065__;
  assign new_new_n1068__ = ~new_new_n1066__ & ~new_new_n1067__;
  assign new_new_n1069__ = ~new_new_n970__ & new_new_n1068__;
  assign new_new_n1070__ = new_new_n970__ & ~new_new_n1068__;
  assign new_new_n1071__ = ~new_new_n1069__ & ~new_new_n1070__;
  assign new_new_n1072__ = ~new_new_n969__ & new_new_n1071__;
  assign new_new_n1073__ = new_new_n969__ & ~new_new_n1071__;
  assign new_new_n1074__ = ~new_new_n1072__ & ~new_new_n1073__;
  assign new_new_n1075__ = ~new_new_n968__ & new_new_n1074__;
  assign new_new_n1076__ = new_new_n968__ & ~new_new_n1074__;
  assign new_new_n1077__ = ~new_new_n1075__ & ~new_new_n1076__;
  assign new_new_n1078__ = ~new_new_n967__ & new_new_n1077__;
  assign new_new_n1079__ = new_new_n967__ & ~new_new_n1077__;
  assign G6150gat = ~new_new_n1078__ & ~new_new_n1079__;
  assign new_new_n1081__ = ~new_new_n1072__ & ~new_new_n1075__;
  assign new_new_n1082__ = G35gat & G528gat;
  assign new_new_n1083__ = ~new_new_n1066__ & ~new_new_n1069__;
  assign new_new_n1084__ = G52gat & G511gat;
  assign new_new_n1085__ = ~new_new_n1060__ & ~new_new_n1063__;
  assign new_new_n1086__ = G69gat & G494gat;
  assign new_new_n1087__ = ~new_new_n1054__ & ~new_new_n1057__;
  assign new_new_n1088__ = G86gat & G477gat;
  assign new_new_n1089__ = ~new_new_n1048__ & ~new_new_n1051__;
  assign new_new_n1090__ = G103gat & G460gat;
  assign new_new_n1091__ = ~new_new_n1042__ & ~new_new_n1045__;
  assign new_new_n1092__ = G120gat & G443gat;
  assign new_new_n1093__ = ~new_new_n1036__ & ~new_new_n1039__;
  assign new_new_n1094__ = G137gat & G426gat;
  assign new_new_n1095__ = ~new_new_n1030__ & ~new_new_n1033__;
  assign new_new_n1096__ = G154gat & G409gat;
  assign new_new_n1097__ = ~new_new_n1024__ & ~new_new_n1027__;
  assign new_new_n1098__ = G171gat & G392gat;
  assign new_new_n1099__ = ~new_new_n1018__ & ~new_new_n1021__;
  assign new_new_n1100__ = G188gat & G375gat;
  assign new_new_n1101__ = ~new_new_n1012__ & ~new_new_n1015__;
  assign new_new_n1102__ = G205gat & G358gat;
  assign new_new_n1103__ = ~new_new_n1006__ & ~new_new_n1009__;
  assign new_new_n1104__ = G222gat & G341gat;
  assign new_new_n1105__ = ~new_new_n1000__ & ~new_new_n1003__;
  assign new_new_n1106__ = G239gat & G324gat;
  assign new_new_n1107__ = G256gat & G307gat;
  assign new_new_n1108__ = new_new_n995__ & ~new_new_n997__;
  assign new_new_n1109__ = ~new_new_n1107__ & ~new_new_n1108__;
  assign new_new_n1110__ = G307gat & new_new_n1108__;
  assign new_new_n1111__ = ~new_new_n1109__ & ~new_new_n1110__;
  assign new_new_n1112__ = ~new_new_n1106__ & new_new_n1111__;
  assign new_new_n1113__ = new_new_n1106__ & ~new_new_n1111__;
  assign new_new_n1114__ = ~new_new_n1112__ & ~new_new_n1113__;
  assign new_new_n1115__ = ~new_new_n1105__ & new_new_n1114__;
  assign new_new_n1116__ = new_new_n1105__ & ~new_new_n1114__;
  assign new_new_n1117__ = ~new_new_n1115__ & ~new_new_n1116__;
  assign new_new_n1118__ = ~new_new_n1104__ & new_new_n1117__;
  assign new_new_n1119__ = new_new_n1104__ & ~new_new_n1117__;
  assign new_new_n1120__ = ~new_new_n1118__ & ~new_new_n1119__;
  assign new_new_n1121__ = ~new_new_n1103__ & new_new_n1120__;
  assign new_new_n1122__ = new_new_n1103__ & ~new_new_n1120__;
  assign new_new_n1123__ = ~new_new_n1121__ & ~new_new_n1122__;
  assign new_new_n1124__ = ~new_new_n1102__ & new_new_n1123__;
  assign new_new_n1125__ = new_new_n1102__ & ~new_new_n1123__;
  assign new_new_n1126__ = ~new_new_n1124__ & ~new_new_n1125__;
  assign new_new_n1127__ = ~new_new_n1101__ & new_new_n1126__;
  assign new_new_n1128__ = new_new_n1101__ & ~new_new_n1126__;
  assign new_new_n1129__ = ~new_new_n1127__ & ~new_new_n1128__;
  assign new_new_n1130__ = ~new_new_n1100__ & new_new_n1129__;
  assign new_new_n1131__ = new_new_n1100__ & ~new_new_n1129__;
  assign new_new_n1132__ = ~new_new_n1130__ & ~new_new_n1131__;
  assign new_new_n1133__ = ~new_new_n1099__ & new_new_n1132__;
  assign new_new_n1134__ = new_new_n1099__ & ~new_new_n1132__;
  assign new_new_n1135__ = ~new_new_n1133__ & ~new_new_n1134__;
  assign new_new_n1136__ = ~new_new_n1098__ & new_new_n1135__;
  assign new_new_n1137__ = new_new_n1098__ & ~new_new_n1135__;
  assign new_new_n1138__ = ~new_new_n1136__ & ~new_new_n1137__;
  assign new_new_n1139__ = ~new_new_n1097__ & new_new_n1138__;
  assign new_new_n1140__ = new_new_n1097__ & ~new_new_n1138__;
  assign new_new_n1141__ = ~new_new_n1139__ & ~new_new_n1140__;
  assign new_new_n1142__ = ~new_new_n1096__ & new_new_n1141__;
  assign new_new_n1143__ = new_new_n1096__ & ~new_new_n1141__;
  assign new_new_n1144__ = ~new_new_n1142__ & ~new_new_n1143__;
  assign new_new_n1145__ = ~new_new_n1095__ & new_new_n1144__;
  assign new_new_n1146__ = new_new_n1095__ & ~new_new_n1144__;
  assign new_new_n1147__ = ~new_new_n1145__ & ~new_new_n1146__;
  assign new_new_n1148__ = ~new_new_n1094__ & new_new_n1147__;
  assign new_new_n1149__ = new_new_n1094__ & ~new_new_n1147__;
  assign new_new_n1150__ = ~new_new_n1148__ & ~new_new_n1149__;
  assign new_new_n1151__ = ~new_new_n1093__ & new_new_n1150__;
  assign new_new_n1152__ = new_new_n1093__ & ~new_new_n1150__;
  assign new_new_n1153__ = ~new_new_n1151__ & ~new_new_n1152__;
  assign new_new_n1154__ = ~new_new_n1092__ & new_new_n1153__;
  assign new_new_n1155__ = new_new_n1092__ & ~new_new_n1153__;
  assign new_new_n1156__ = ~new_new_n1154__ & ~new_new_n1155__;
  assign new_new_n1157__ = ~new_new_n1091__ & new_new_n1156__;
  assign new_new_n1158__ = new_new_n1091__ & ~new_new_n1156__;
  assign new_new_n1159__ = ~new_new_n1157__ & ~new_new_n1158__;
  assign new_new_n1160__ = ~new_new_n1090__ & new_new_n1159__;
  assign new_new_n1161__ = new_new_n1090__ & ~new_new_n1159__;
  assign new_new_n1162__ = ~new_new_n1160__ & ~new_new_n1161__;
  assign new_new_n1163__ = ~new_new_n1089__ & new_new_n1162__;
  assign new_new_n1164__ = new_new_n1089__ & ~new_new_n1162__;
  assign new_new_n1165__ = ~new_new_n1163__ & ~new_new_n1164__;
  assign new_new_n1166__ = ~new_new_n1088__ & new_new_n1165__;
  assign new_new_n1167__ = new_new_n1088__ & ~new_new_n1165__;
  assign new_new_n1168__ = ~new_new_n1166__ & ~new_new_n1167__;
  assign new_new_n1169__ = ~new_new_n1087__ & new_new_n1168__;
  assign new_new_n1170__ = new_new_n1087__ & ~new_new_n1168__;
  assign new_new_n1171__ = ~new_new_n1169__ & ~new_new_n1170__;
  assign new_new_n1172__ = ~new_new_n1086__ & new_new_n1171__;
  assign new_new_n1173__ = new_new_n1086__ & ~new_new_n1171__;
  assign new_new_n1174__ = ~new_new_n1172__ & ~new_new_n1173__;
  assign new_new_n1175__ = ~new_new_n1085__ & new_new_n1174__;
  assign new_new_n1176__ = new_new_n1085__ & ~new_new_n1174__;
  assign new_new_n1177__ = ~new_new_n1175__ & ~new_new_n1176__;
  assign new_new_n1178__ = ~new_new_n1084__ & new_new_n1177__;
  assign new_new_n1179__ = new_new_n1084__ & ~new_new_n1177__;
  assign new_new_n1180__ = ~new_new_n1178__ & ~new_new_n1179__;
  assign new_new_n1181__ = ~new_new_n1083__ & new_new_n1180__;
  assign new_new_n1182__ = new_new_n1083__ & ~new_new_n1180__;
  assign new_new_n1183__ = ~new_new_n1181__ & ~new_new_n1182__;
  assign new_new_n1184__ = ~new_new_n1082__ & new_new_n1183__;
  assign new_new_n1185__ = new_new_n1082__ & ~new_new_n1183__;
  assign new_new_n1186__ = ~new_new_n1184__ & ~new_new_n1185__;
  assign new_new_n1187__ = ~new_new_n1081__ & new_new_n1186__;
  assign new_new_n1188__ = new_new_n1081__ & ~new_new_n1186__;
  assign new_new_n1189__ = ~new_new_n1187__ & ~new_new_n1188__;
  assign new_new_n1190__ = ~new_new_n1079__ & new_new_n1189__;
  assign new_new_n1191__ = new_new_n1079__ & ~new_new_n1189__;
  assign G6160gat = new_new_n1190__ | new_new_n1191__;
  assign new_new_n1193__ = ~new_new_n1187__ & ~new_new_n1190__;
  assign new_new_n1194__ = ~new_new_n1181__ & ~new_new_n1184__;
  assign new_new_n1195__ = G52gat & G528gat;
  assign new_new_n1196__ = ~new_new_n1175__ & ~new_new_n1178__;
  assign new_new_n1197__ = G69gat & G511gat;
  assign new_new_n1198__ = ~new_new_n1169__ & ~new_new_n1172__;
  assign new_new_n1199__ = G86gat & G494gat;
  assign new_new_n1200__ = ~new_new_n1163__ & ~new_new_n1166__;
  assign new_new_n1201__ = G103gat & G477gat;
  assign new_new_n1202__ = ~new_new_n1157__ & ~new_new_n1160__;
  assign new_new_n1203__ = G120gat & G460gat;
  assign new_new_n1204__ = ~new_new_n1151__ & ~new_new_n1154__;
  assign new_new_n1205__ = G137gat & G443gat;
  assign new_new_n1206__ = ~new_new_n1145__ & ~new_new_n1148__;
  assign new_new_n1207__ = G154gat & G426gat;
  assign new_new_n1208__ = ~new_new_n1139__ & ~new_new_n1142__;
  assign new_new_n1209__ = G171gat & G409gat;
  assign new_new_n1210__ = ~new_new_n1133__ & ~new_new_n1136__;
  assign new_new_n1211__ = G188gat & G392gat;
  assign new_new_n1212__ = ~new_new_n1127__ & ~new_new_n1130__;
  assign new_new_n1213__ = G205gat & G375gat;
  assign new_new_n1214__ = ~new_new_n1121__ & ~new_new_n1124__;
  assign new_new_n1215__ = G222gat & G358gat;
  assign new_new_n1216__ = ~new_new_n1115__ & ~new_new_n1118__;
  assign new_new_n1217__ = G239gat & G341gat;
  assign new_new_n1218__ = G256gat & G324gat;
  assign new_new_n1219__ = ~new_new_n1109__ & ~new_new_n1112__;
  assign new_new_n1220__ = ~new_new_n1218__ & ~new_new_n1219__;
  assign new_new_n1221__ = new_new_n1218__ & new_new_n1219__;
  assign new_new_n1222__ = ~new_new_n1220__ & ~new_new_n1221__;
  assign new_new_n1223__ = ~new_new_n1217__ & new_new_n1222__;
  assign new_new_n1224__ = new_new_n1217__ & ~new_new_n1222__;
  assign new_new_n1225__ = ~new_new_n1223__ & ~new_new_n1224__;
  assign new_new_n1226__ = ~new_new_n1216__ & new_new_n1225__;
  assign new_new_n1227__ = new_new_n1216__ & ~new_new_n1225__;
  assign new_new_n1228__ = ~new_new_n1226__ & ~new_new_n1227__;
  assign new_new_n1229__ = ~new_new_n1215__ & new_new_n1228__;
  assign new_new_n1230__ = new_new_n1215__ & ~new_new_n1228__;
  assign new_new_n1231__ = ~new_new_n1229__ & ~new_new_n1230__;
  assign new_new_n1232__ = ~new_new_n1214__ & new_new_n1231__;
  assign new_new_n1233__ = new_new_n1214__ & ~new_new_n1231__;
  assign new_new_n1234__ = ~new_new_n1232__ & ~new_new_n1233__;
  assign new_new_n1235__ = ~new_new_n1213__ & new_new_n1234__;
  assign new_new_n1236__ = new_new_n1213__ & ~new_new_n1234__;
  assign new_new_n1237__ = ~new_new_n1235__ & ~new_new_n1236__;
  assign new_new_n1238__ = ~new_new_n1212__ & new_new_n1237__;
  assign new_new_n1239__ = new_new_n1212__ & ~new_new_n1237__;
  assign new_new_n1240__ = ~new_new_n1238__ & ~new_new_n1239__;
  assign new_new_n1241__ = ~new_new_n1211__ & new_new_n1240__;
  assign new_new_n1242__ = new_new_n1211__ & ~new_new_n1240__;
  assign new_new_n1243__ = ~new_new_n1241__ & ~new_new_n1242__;
  assign new_new_n1244__ = ~new_new_n1210__ & new_new_n1243__;
  assign new_new_n1245__ = new_new_n1210__ & ~new_new_n1243__;
  assign new_new_n1246__ = ~new_new_n1244__ & ~new_new_n1245__;
  assign new_new_n1247__ = ~new_new_n1209__ & new_new_n1246__;
  assign new_new_n1248__ = new_new_n1209__ & ~new_new_n1246__;
  assign new_new_n1249__ = ~new_new_n1247__ & ~new_new_n1248__;
  assign new_new_n1250__ = ~new_new_n1208__ & new_new_n1249__;
  assign new_new_n1251__ = new_new_n1208__ & ~new_new_n1249__;
  assign new_new_n1252__ = ~new_new_n1250__ & ~new_new_n1251__;
  assign new_new_n1253__ = ~new_new_n1207__ & new_new_n1252__;
  assign new_new_n1254__ = new_new_n1207__ & ~new_new_n1252__;
  assign new_new_n1255__ = ~new_new_n1253__ & ~new_new_n1254__;
  assign new_new_n1256__ = ~new_new_n1206__ & new_new_n1255__;
  assign new_new_n1257__ = new_new_n1206__ & ~new_new_n1255__;
  assign new_new_n1258__ = ~new_new_n1256__ & ~new_new_n1257__;
  assign new_new_n1259__ = ~new_new_n1205__ & new_new_n1258__;
  assign new_new_n1260__ = new_new_n1205__ & ~new_new_n1258__;
  assign new_new_n1261__ = ~new_new_n1259__ & ~new_new_n1260__;
  assign new_new_n1262__ = ~new_new_n1204__ & new_new_n1261__;
  assign new_new_n1263__ = new_new_n1204__ & ~new_new_n1261__;
  assign new_new_n1264__ = ~new_new_n1262__ & ~new_new_n1263__;
  assign new_new_n1265__ = ~new_new_n1203__ & new_new_n1264__;
  assign new_new_n1266__ = new_new_n1203__ & ~new_new_n1264__;
  assign new_new_n1267__ = ~new_new_n1265__ & ~new_new_n1266__;
  assign new_new_n1268__ = ~new_new_n1202__ & new_new_n1267__;
  assign new_new_n1269__ = new_new_n1202__ & ~new_new_n1267__;
  assign new_new_n1270__ = ~new_new_n1268__ & ~new_new_n1269__;
  assign new_new_n1271__ = ~new_new_n1201__ & new_new_n1270__;
  assign new_new_n1272__ = new_new_n1201__ & ~new_new_n1270__;
  assign new_new_n1273__ = ~new_new_n1271__ & ~new_new_n1272__;
  assign new_new_n1274__ = ~new_new_n1200__ & new_new_n1273__;
  assign new_new_n1275__ = new_new_n1200__ & ~new_new_n1273__;
  assign new_new_n1276__ = ~new_new_n1274__ & ~new_new_n1275__;
  assign new_new_n1277__ = ~new_new_n1199__ & new_new_n1276__;
  assign new_new_n1278__ = new_new_n1199__ & ~new_new_n1276__;
  assign new_new_n1279__ = ~new_new_n1277__ & ~new_new_n1278__;
  assign new_new_n1280__ = ~new_new_n1198__ & new_new_n1279__;
  assign new_new_n1281__ = new_new_n1198__ & ~new_new_n1279__;
  assign new_new_n1282__ = ~new_new_n1280__ & ~new_new_n1281__;
  assign new_new_n1283__ = ~new_new_n1197__ & new_new_n1282__;
  assign new_new_n1284__ = new_new_n1197__ & ~new_new_n1282__;
  assign new_new_n1285__ = ~new_new_n1283__ & ~new_new_n1284__;
  assign new_new_n1286__ = ~new_new_n1196__ & new_new_n1285__;
  assign new_new_n1287__ = new_new_n1196__ & ~new_new_n1285__;
  assign new_new_n1288__ = ~new_new_n1286__ & ~new_new_n1287__;
  assign new_new_n1289__ = ~new_new_n1195__ & new_new_n1288__;
  assign new_new_n1290__ = new_new_n1195__ & ~new_new_n1288__;
  assign new_new_n1291__ = ~new_new_n1289__ & ~new_new_n1290__;
  assign new_new_n1292__ = ~new_new_n1194__ & new_new_n1291__;
  assign new_new_n1293__ = new_new_n1194__ & ~new_new_n1291__;
  assign new_new_n1294__ = ~new_new_n1292__ & ~new_new_n1293__;
  assign new_new_n1295__ = ~new_new_n1193__ & new_new_n1294__;
  assign new_new_n1296__ = new_new_n1193__ & ~new_new_n1294__;
  assign G6170gat = new_new_n1295__ | new_new_n1296__;
  assign new_new_n1298__ = ~new_new_n1292__ & ~new_new_n1295__;
  assign new_new_n1299__ = ~new_new_n1286__ & ~new_new_n1289__;
  assign new_new_n1300__ = G69gat & G528gat;
  assign new_new_n1301__ = ~new_new_n1280__ & ~new_new_n1283__;
  assign new_new_n1302__ = G86gat & G511gat;
  assign new_new_n1303__ = ~new_new_n1274__ & ~new_new_n1277__;
  assign new_new_n1304__ = G103gat & G494gat;
  assign new_new_n1305__ = ~new_new_n1268__ & ~new_new_n1271__;
  assign new_new_n1306__ = G120gat & G477gat;
  assign new_new_n1307__ = ~new_new_n1262__ & ~new_new_n1265__;
  assign new_new_n1308__ = G137gat & G460gat;
  assign new_new_n1309__ = ~new_new_n1256__ & ~new_new_n1259__;
  assign new_new_n1310__ = G154gat & G443gat;
  assign new_new_n1311__ = ~new_new_n1250__ & ~new_new_n1253__;
  assign new_new_n1312__ = G171gat & G426gat;
  assign new_new_n1313__ = ~new_new_n1244__ & ~new_new_n1247__;
  assign new_new_n1314__ = G188gat & G409gat;
  assign new_new_n1315__ = ~new_new_n1238__ & ~new_new_n1241__;
  assign new_new_n1316__ = G205gat & G392gat;
  assign new_new_n1317__ = ~new_new_n1232__ & ~new_new_n1235__;
  assign new_new_n1318__ = G222gat & G375gat;
  assign new_new_n1319__ = ~new_new_n1226__ & ~new_new_n1229__;
  assign new_new_n1320__ = G239gat & G358gat;
  assign new_new_n1321__ = G256gat & G341gat;
  assign new_new_n1322__ = ~new_new_n1220__ & ~new_new_n1223__;
  assign new_new_n1323__ = ~new_new_n1321__ & ~new_new_n1322__;
  assign new_new_n1324__ = new_new_n1321__ & new_new_n1322__;
  assign new_new_n1325__ = ~new_new_n1323__ & ~new_new_n1324__;
  assign new_new_n1326__ = ~new_new_n1320__ & new_new_n1325__;
  assign new_new_n1327__ = new_new_n1320__ & ~new_new_n1325__;
  assign new_new_n1328__ = ~new_new_n1326__ & ~new_new_n1327__;
  assign new_new_n1329__ = ~new_new_n1319__ & new_new_n1328__;
  assign new_new_n1330__ = new_new_n1319__ & ~new_new_n1328__;
  assign new_new_n1331__ = ~new_new_n1329__ & ~new_new_n1330__;
  assign new_new_n1332__ = ~new_new_n1318__ & new_new_n1331__;
  assign new_new_n1333__ = new_new_n1318__ & ~new_new_n1331__;
  assign new_new_n1334__ = ~new_new_n1332__ & ~new_new_n1333__;
  assign new_new_n1335__ = ~new_new_n1317__ & new_new_n1334__;
  assign new_new_n1336__ = new_new_n1317__ & ~new_new_n1334__;
  assign new_new_n1337__ = ~new_new_n1335__ & ~new_new_n1336__;
  assign new_new_n1338__ = ~new_new_n1316__ & new_new_n1337__;
  assign new_new_n1339__ = new_new_n1316__ & ~new_new_n1337__;
  assign new_new_n1340__ = ~new_new_n1338__ & ~new_new_n1339__;
  assign new_new_n1341__ = ~new_new_n1315__ & new_new_n1340__;
  assign new_new_n1342__ = new_new_n1315__ & ~new_new_n1340__;
  assign new_new_n1343__ = ~new_new_n1341__ & ~new_new_n1342__;
  assign new_new_n1344__ = ~new_new_n1314__ & new_new_n1343__;
  assign new_new_n1345__ = new_new_n1314__ & ~new_new_n1343__;
  assign new_new_n1346__ = ~new_new_n1344__ & ~new_new_n1345__;
  assign new_new_n1347__ = ~new_new_n1313__ & new_new_n1346__;
  assign new_new_n1348__ = new_new_n1313__ & ~new_new_n1346__;
  assign new_new_n1349__ = ~new_new_n1347__ & ~new_new_n1348__;
  assign new_new_n1350__ = ~new_new_n1312__ & new_new_n1349__;
  assign new_new_n1351__ = new_new_n1312__ & ~new_new_n1349__;
  assign new_new_n1352__ = ~new_new_n1350__ & ~new_new_n1351__;
  assign new_new_n1353__ = ~new_new_n1311__ & new_new_n1352__;
  assign new_new_n1354__ = new_new_n1311__ & ~new_new_n1352__;
  assign new_new_n1355__ = ~new_new_n1353__ & ~new_new_n1354__;
  assign new_new_n1356__ = ~new_new_n1310__ & new_new_n1355__;
  assign new_new_n1357__ = new_new_n1310__ & ~new_new_n1355__;
  assign new_new_n1358__ = ~new_new_n1356__ & ~new_new_n1357__;
  assign new_new_n1359__ = ~new_new_n1309__ & new_new_n1358__;
  assign new_new_n1360__ = new_new_n1309__ & ~new_new_n1358__;
  assign new_new_n1361__ = ~new_new_n1359__ & ~new_new_n1360__;
  assign new_new_n1362__ = ~new_new_n1308__ & new_new_n1361__;
  assign new_new_n1363__ = new_new_n1308__ & ~new_new_n1361__;
  assign new_new_n1364__ = ~new_new_n1362__ & ~new_new_n1363__;
  assign new_new_n1365__ = ~new_new_n1307__ & new_new_n1364__;
  assign new_new_n1366__ = new_new_n1307__ & ~new_new_n1364__;
  assign new_new_n1367__ = ~new_new_n1365__ & ~new_new_n1366__;
  assign new_new_n1368__ = ~new_new_n1306__ & new_new_n1367__;
  assign new_new_n1369__ = new_new_n1306__ & ~new_new_n1367__;
  assign new_new_n1370__ = ~new_new_n1368__ & ~new_new_n1369__;
  assign new_new_n1371__ = ~new_new_n1305__ & new_new_n1370__;
  assign new_new_n1372__ = new_new_n1305__ & ~new_new_n1370__;
  assign new_new_n1373__ = ~new_new_n1371__ & ~new_new_n1372__;
  assign new_new_n1374__ = ~new_new_n1304__ & new_new_n1373__;
  assign new_new_n1375__ = new_new_n1304__ & ~new_new_n1373__;
  assign new_new_n1376__ = ~new_new_n1374__ & ~new_new_n1375__;
  assign new_new_n1377__ = ~new_new_n1303__ & new_new_n1376__;
  assign new_new_n1378__ = new_new_n1303__ & ~new_new_n1376__;
  assign new_new_n1379__ = ~new_new_n1377__ & ~new_new_n1378__;
  assign new_new_n1380__ = ~new_new_n1302__ & new_new_n1379__;
  assign new_new_n1381__ = new_new_n1302__ & ~new_new_n1379__;
  assign new_new_n1382__ = ~new_new_n1380__ & ~new_new_n1381__;
  assign new_new_n1383__ = ~new_new_n1301__ & new_new_n1382__;
  assign new_new_n1384__ = new_new_n1301__ & ~new_new_n1382__;
  assign new_new_n1385__ = ~new_new_n1383__ & ~new_new_n1384__;
  assign new_new_n1386__ = ~new_new_n1300__ & new_new_n1385__;
  assign new_new_n1387__ = new_new_n1300__ & ~new_new_n1385__;
  assign new_new_n1388__ = ~new_new_n1386__ & ~new_new_n1387__;
  assign new_new_n1389__ = ~new_new_n1299__ & new_new_n1388__;
  assign new_new_n1390__ = new_new_n1299__ & ~new_new_n1388__;
  assign new_new_n1391__ = ~new_new_n1389__ & ~new_new_n1390__;
  assign new_new_n1392__ = ~new_new_n1298__ & new_new_n1391__;
  assign new_new_n1393__ = new_new_n1298__ & ~new_new_n1391__;
  assign G6180gat = new_new_n1392__ | new_new_n1393__;
  assign new_new_n1395__ = ~new_new_n1389__ & ~new_new_n1392__;
  assign new_new_n1396__ = ~new_new_n1383__ & ~new_new_n1386__;
  assign new_new_n1397__ = G86gat & G528gat;
  assign new_new_n1398__ = ~new_new_n1377__ & ~new_new_n1380__;
  assign new_new_n1399__ = G103gat & G511gat;
  assign new_new_n1400__ = ~new_new_n1371__ & ~new_new_n1374__;
  assign new_new_n1401__ = G120gat & G494gat;
  assign new_new_n1402__ = ~new_new_n1365__ & ~new_new_n1368__;
  assign new_new_n1403__ = G137gat & G477gat;
  assign new_new_n1404__ = ~new_new_n1359__ & ~new_new_n1362__;
  assign new_new_n1405__ = G154gat & G460gat;
  assign new_new_n1406__ = ~new_new_n1353__ & ~new_new_n1356__;
  assign new_new_n1407__ = G171gat & G443gat;
  assign new_new_n1408__ = ~new_new_n1347__ & ~new_new_n1350__;
  assign new_new_n1409__ = G188gat & G426gat;
  assign new_new_n1410__ = ~new_new_n1341__ & ~new_new_n1344__;
  assign new_new_n1411__ = G205gat & G409gat;
  assign new_new_n1412__ = ~new_new_n1335__ & ~new_new_n1338__;
  assign new_new_n1413__ = G222gat & G392gat;
  assign new_new_n1414__ = ~new_new_n1329__ & ~new_new_n1332__;
  assign new_new_n1415__ = G239gat & G375gat;
  assign new_new_n1416__ = G256gat & G358gat;
  assign new_new_n1417__ = ~new_new_n1323__ & ~new_new_n1326__;
  assign new_new_n1418__ = ~new_new_n1416__ & ~new_new_n1417__;
  assign new_new_n1419__ = new_new_n1416__ & new_new_n1417__;
  assign new_new_n1420__ = ~new_new_n1418__ & ~new_new_n1419__;
  assign new_new_n1421__ = ~new_new_n1415__ & new_new_n1420__;
  assign new_new_n1422__ = new_new_n1415__ & ~new_new_n1420__;
  assign new_new_n1423__ = ~new_new_n1421__ & ~new_new_n1422__;
  assign new_new_n1424__ = ~new_new_n1414__ & new_new_n1423__;
  assign new_new_n1425__ = new_new_n1414__ & ~new_new_n1423__;
  assign new_new_n1426__ = ~new_new_n1424__ & ~new_new_n1425__;
  assign new_new_n1427__ = ~new_new_n1413__ & new_new_n1426__;
  assign new_new_n1428__ = new_new_n1413__ & ~new_new_n1426__;
  assign new_new_n1429__ = ~new_new_n1427__ & ~new_new_n1428__;
  assign new_new_n1430__ = ~new_new_n1412__ & new_new_n1429__;
  assign new_new_n1431__ = new_new_n1412__ & ~new_new_n1429__;
  assign new_new_n1432__ = ~new_new_n1430__ & ~new_new_n1431__;
  assign new_new_n1433__ = ~new_new_n1411__ & new_new_n1432__;
  assign new_new_n1434__ = new_new_n1411__ & ~new_new_n1432__;
  assign new_new_n1435__ = ~new_new_n1433__ & ~new_new_n1434__;
  assign new_new_n1436__ = ~new_new_n1410__ & new_new_n1435__;
  assign new_new_n1437__ = new_new_n1410__ & ~new_new_n1435__;
  assign new_new_n1438__ = ~new_new_n1436__ & ~new_new_n1437__;
  assign new_new_n1439__ = ~new_new_n1409__ & new_new_n1438__;
  assign new_new_n1440__ = new_new_n1409__ & ~new_new_n1438__;
  assign new_new_n1441__ = ~new_new_n1439__ & ~new_new_n1440__;
  assign new_new_n1442__ = ~new_new_n1408__ & new_new_n1441__;
  assign new_new_n1443__ = new_new_n1408__ & ~new_new_n1441__;
  assign new_new_n1444__ = ~new_new_n1442__ & ~new_new_n1443__;
  assign new_new_n1445__ = ~new_new_n1407__ & new_new_n1444__;
  assign new_new_n1446__ = new_new_n1407__ & ~new_new_n1444__;
  assign new_new_n1447__ = ~new_new_n1445__ & ~new_new_n1446__;
  assign new_new_n1448__ = ~new_new_n1406__ & new_new_n1447__;
  assign new_new_n1449__ = new_new_n1406__ & ~new_new_n1447__;
  assign new_new_n1450__ = ~new_new_n1448__ & ~new_new_n1449__;
  assign new_new_n1451__ = ~new_new_n1405__ & new_new_n1450__;
  assign new_new_n1452__ = new_new_n1405__ & ~new_new_n1450__;
  assign new_new_n1453__ = ~new_new_n1451__ & ~new_new_n1452__;
  assign new_new_n1454__ = ~new_new_n1404__ & new_new_n1453__;
  assign new_new_n1455__ = new_new_n1404__ & ~new_new_n1453__;
  assign new_new_n1456__ = ~new_new_n1454__ & ~new_new_n1455__;
  assign new_new_n1457__ = ~new_new_n1403__ & new_new_n1456__;
  assign new_new_n1458__ = new_new_n1403__ & ~new_new_n1456__;
  assign new_new_n1459__ = ~new_new_n1457__ & ~new_new_n1458__;
  assign new_new_n1460__ = ~new_new_n1402__ & new_new_n1459__;
  assign new_new_n1461__ = new_new_n1402__ & ~new_new_n1459__;
  assign new_new_n1462__ = ~new_new_n1460__ & ~new_new_n1461__;
  assign new_new_n1463__ = ~new_new_n1401__ & new_new_n1462__;
  assign new_new_n1464__ = new_new_n1401__ & ~new_new_n1462__;
  assign new_new_n1465__ = ~new_new_n1463__ & ~new_new_n1464__;
  assign new_new_n1466__ = ~new_new_n1400__ & new_new_n1465__;
  assign new_new_n1467__ = new_new_n1400__ & ~new_new_n1465__;
  assign new_new_n1468__ = ~new_new_n1466__ & ~new_new_n1467__;
  assign new_new_n1469__ = ~new_new_n1399__ & new_new_n1468__;
  assign new_new_n1470__ = new_new_n1399__ & ~new_new_n1468__;
  assign new_new_n1471__ = ~new_new_n1469__ & ~new_new_n1470__;
  assign new_new_n1472__ = ~new_new_n1398__ & new_new_n1471__;
  assign new_new_n1473__ = new_new_n1398__ & ~new_new_n1471__;
  assign new_new_n1474__ = ~new_new_n1472__ & ~new_new_n1473__;
  assign new_new_n1475__ = ~new_new_n1397__ & new_new_n1474__;
  assign new_new_n1476__ = new_new_n1397__ & ~new_new_n1474__;
  assign new_new_n1477__ = ~new_new_n1475__ & ~new_new_n1476__;
  assign new_new_n1478__ = ~new_new_n1396__ & new_new_n1477__;
  assign new_new_n1479__ = new_new_n1396__ & ~new_new_n1477__;
  assign new_new_n1480__ = ~new_new_n1478__ & ~new_new_n1479__;
  assign new_new_n1481__ = ~new_new_n1395__ & new_new_n1480__;
  assign new_new_n1482__ = new_new_n1395__ & ~new_new_n1480__;
  assign G6190gat = new_new_n1481__ | new_new_n1482__;
  assign new_new_n1484__ = ~new_new_n1478__ & ~new_new_n1481__;
  assign new_new_n1485__ = ~new_new_n1472__ & ~new_new_n1475__;
  assign new_new_n1486__ = G103gat & G528gat;
  assign new_new_n1487__ = ~new_new_n1466__ & ~new_new_n1469__;
  assign new_new_n1488__ = G120gat & G511gat;
  assign new_new_n1489__ = ~new_new_n1460__ & ~new_new_n1463__;
  assign new_new_n1490__ = G137gat & G494gat;
  assign new_new_n1491__ = ~new_new_n1454__ & ~new_new_n1457__;
  assign new_new_n1492__ = G154gat & G477gat;
  assign new_new_n1493__ = ~new_new_n1448__ & ~new_new_n1451__;
  assign new_new_n1494__ = G171gat & G460gat;
  assign new_new_n1495__ = ~new_new_n1442__ & ~new_new_n1445__;
  assign new_new_n1496__ = G188gat & G443gat;
  assign new_new_n1497__ = ~new_new_n1436__ & ~new_new_n1439__;
  assign new_new_n1498__ = G205gat & G426gat;
  assign new_new_n1499__ = ~new_new_n1430__ & ~new_new_n1433__;
  assign new_new_n1500__ = G222gat & G409gat;
  assign new_new_n1501__ = ~new_new_n1424__ & ~new_new_n1427__;
  assign new_new_n1502__ = G239gat & G392gat;
  assign new_new_n1503__ = G256gat & G375gat;
  assign new_new_n1504__ = ~new_new_n1418__ & ~new_new_n1421__;
  assign new_new_n1505__ = ~new_new_n1503__ & ~new_new_n1504__;
  assign new_new_n1506__ = new_new_n1503__ & new_new_n1504__;
  assign new_new_n1507__ = ~new_new_n1505__ & ~new_new_n1506__;
  assign new_new_n1508__ = ~new_new_n1502__ & new_new_n1507__;
  assign new_new_n1509__ = new_new_n1502__ & ~new_new_n1507__;
  assign new_new_n1510__ = ~new_new_n1508__ & ~new_new_n1509__;
  assign new_new_n1511__ = ~new_new_n1501__ & new_new_n1510__;
  assign new_new_n1512__ = new_new_n1501__ & ~new_new_n1510__;
  assign new_new_n1513__ = ~new_new_n1511__ & ~new_new_n1512__;
  assign new_new_n1514__ = ~new_new_n1500__ & new_new_n1513__;
  assign new_new_n1515__ = new_new_n1500__ & ~new_new_n1513__;
  assign new_new_n1516__ = ~new_new_n1514__ & ~new_new_n1515__;
  assign new_new_n1517__ = ~new_new_n1499__ & new_new_n1516__;
  assign new_new_n1518__ = new_new_n1499__ & ~new_new_n1516__;
  assign new_new_n1519__ = ~new_new_n1517__ & ~new_new_n1518__;
  assign new_new_n1520__ = ~new_new_n1498__ & new_new_n1519__;
  assign new_new_n1521__ = new_new_n1498__ & ~new_new_n1519__;
  assign new_new_n1522__ = ~new_new_n1520__ & ~new_new_n1521__;
  assign new_new_n1523__ = ~new_new_n1497__ & new_new_n1522__;
  assign new_new_n1524__ = new_new_n1497__ & ~new_new_n1522__;
  assign new_new_n1525__ = ~new_new_n1523__ & ~new_new_n1524__;
  assign new_new_n1526__ = ~new_new_n1496__ & new_new_n1525__;
  assign new_new_n1527__ = new_new_n1496__ & ~new_new_n1525__;
  assign new_new_n1528__ = ~new_new_n1526__ & ~new_new_n1527__;
  assign new_new_n1529__ = ~new_new_n1495__ & new_new_n1528__;
  assign new_new_n1530__ = new_new_n1495__ & ~new_new_n1528__;
  assign new_new_n1531__ = ~new_new_n1529__ & ~new_new_n1530__;
  assign new_new_n1532__ = ~new_new_n1494__ & new_new_n1531__;
  assign new_new_n1533__ = new_new_n1494__ & ~new_new_n1531__;
  assign new_new_n1534__ = ~new_new_n1532__ & ~new_new_n1533__;
  assign new_new_n1535__ = ~new_new_n1493__ & new_new_n1534__;
  assign new_new_n1536__ = new_new_n1493__ & ~new_new_n1534__;
  assign new_new_n1537__ = ~new_new_n1535__ & ~new_new_n1536__;
  assign new_new_n1538__ = ~new_new_n1492__ & new_new_n1537__;
  assign new_new_n1539__ = new_new_n1492__ & ~new_new_n1537__;
  assign new_new_n1540__ = ~new_new_n1538__ & ~new_new_n1539__;
  assign new_new_n1541__ = ~new_new_n1491__ & new_new_n1540__;
  assign new_new_n1542__ = new_new_n1491__ & ~new_new_n1540__;
  assign new_new_n1543__ = ~new_new_n1541__ & ~new_new_n1542__;
  assign new_new_n1544__ = ~new_new_n1490__ & new_new_n1543__;
  assign new_new_n1545__ = new_new_n1490__ & ~new_new_n1543__;
  assign new_new_n1546__ = ~new_new_n1544__ & ~new_new_n1545__;
  assign new_new_n1547__ = ~new_new_n1489__ & new_new_n1546__;
  assign new_new_n1548__ = new_new_n1489__ & ~new_new_n1546__;
  assign new_new_n1549__ = ~new_new_n1547__ & ~new_new_n1548__;
  assign new_new_n1550__ = ~new_new_n1488__ & new_new_n1549__;
  assign new_new_n1551__ = new_new_n1488__ & ~new_new_n1549__;
  assign new_new_n1552__ = ~new_new_n1550__ & ~new_new_n1551__;
  assign new_new_n1553__ = ~new_new_n1487__ & new_new_n1552__;
  assign new_new_n1554__ = new_new_n1487__ & ~new_new_n1552__;
  assign new_new_n1555__ = ~new_new_n1553__ & ~new_new_n1554__;
  assign new_new_n1556__ = ~new_new_n1486__ & new_new_n1555__;
  assign new_new_n1557__ = new_new_n1486__ & ~new_new_n1555__;
  assign new_new_n1558__ = ~new_new_n1556__ & ~new_new_n1557__;
  assign new_new_n1559__ = ~new_new_n1485__ & new_new_n1558__;
  assign new_new_n1560__ = new_new_n1485__ & ~new_new_n1558__;
  assign new_new_n1561__ = ~new_new_n1559__ & ~new_new_n1560__;
  assign new_new_n1562__ = ~new_new_n1484__ & new_new_n1561__;
  assign new_new_n1563__ = new_new_n1484__ & ~new_new_n1561__;
  assign G6200gat = new_new_n1562__ | new_new_n1563__;
  assign new_new_n1565__ = ~new_new_n1559__ & ~new_new_n1562__;
  assign new_new_n1566__ = ~new_new_n1553__ & ~new_new_n1556__;
  assign new_new_n1567__ = G120gat & G528gat;
  assign new_new_n1568__ = ~new_new_n1547__ & ~new_new_n1550__;
  assign new_new_n1569__ = G137gat & G511gat;
  assign new_new_n1570__ = ~new_new_n1541__ & ~new_new_n1544__;
  assign new_new_n1571__ = G154gat & G494gat;
  assign new_new_n1572__ = ~new_new_n1535__ & ~new_new_n1538__;
  assign new_new_n1573__ = G171gat & G477gat;
  assign new_new_n1574__ = ~new_new_n1529__ & ~new_new_n1532__;
  assign new_new_n1575__ = G188gat & G460gat;
  assign new_new_n1576__ = ~new_new_n1523__ & ~new_new_n1526__;
  assign new_new_n1577__ = G205gat & G443gat;
  assign new_new_n1578__ = ~new_new_n1517__ & ~new_new_n1520__;
  assign new_new_n1579__ = G222gat & G426gat;
  assign new_new_n1580__ = ~new_new_n1511__ & ~new_new_n1514__;
  assign new_new_n1581__ = G239gat & G409gat;
  assign new_new_n1582__ = G256gat & G392gat;
  assign new_new_n1583__ = ~new_new_n1505__ & ~new_new_n1508__;
  assign new_new_n1584__ = ~new_new_n1582__ & ~new_new_n1583__;
  assign new_new_n1585__ = new_new_n1582__ & new_new_n1583__;
  assign new_new_n1586__ = ~new_new_n1584__ & ~new_new_n1585__;
  assign new_new_n1587__ = ~new_new_n1581__ & new_new_n1586__;
  assign new_new_n1588__ = new_new_n1581__ & ~new_new_n1586__;
  assign new_new_n1589__ = ~new_new_n1587__ & ~new_new_n1588__;
  assign new_new_n1590__ = ~new_new_n1580__ & new_new_n1589__;
  assign new_new_n1591__ = new_new_n1580__ & ~new_new_n1589__;
  assign new_new_n1592__ = ~new_new_n1590__ & ~new_new_n1591__;
  assign new_new_n1593__ = ~new_new_n1579__ & new_new_n1592__;
  assign new_new_n1594__ = new_new_n1579__ & ~new_new_n1592__;
  assign new_new_n1595__ = ~new_new_n1593__ & ~new_new_n1594__;
  assign new_new_n1596__ = ~new_new_n1578__ & new_new_n1595__;
  assign new_new_n1597__ = new_new_n1578__ & ~new_new_n1595__;
  assign new_new_n1598__ = ~new_new_n1596__ & ~new_new_n1597__;
  assign new_new_n1599__ = ~new_new_n1577__ & new_new_n1598__;
  assign new_new_n1600__ = new_new_n1577__ & ~new_new_n1598__;
  assign new_new_n1601__ = ~new_new_n1599__ & ~new_new_n1600__;
  assign new_new_n1602__ = ~new_new_n1576__ & new_new_n1601__;
  assign new_new_n1603__ = new_new_n1576__ & ~new_new_n1601__;
  assign new_new_n1604__ = ~new_new_n1602__ & ~new_new_n1603__;
  assign new_new_n1605__ = ~new_new_n1575__ & new_new_n1604__;
  assign new_new_n1606__ = new_new_n1575__ & ~new_new_n1604__;
  assign new_new_n1607__ = ~new_new_n1605__ & ~new_new_n1606__;
  assign new_new_n1608__ = ~new_new_n1574__ & new_new_n1607__;
  assign new_new_n1609__ = new_new_n1574__ & ~new_new_n1607__;
  assign new_new_n1610__ = ~new_new_n1608__ & ~new_new_n1609__;
  assign new_new_n1611__ = ~new_new_n1573__ & new_new_n1610__;
  assign new_new_n1612__ = new_new_n1573__ & ~new_new_n1610__;
  assign new_new_n1613__ = ~new_new_n1611__ & ~new_new_n1612__;
  assign new_new_n1614__ = ~new_new_n1572__ & new_new_n1613__;
  assign new_new_n1615__ = new_new_n1572__ & ~new_new_n1613__;
  assign new_new_n1616__ = ~new_new_n1614__ & ~new_new_n1615__;
  assign new_new_n1617__ = ~new_new_n1571__ & new_new_n1616__;
  assign new_new_n1618__ = new_new_n1571__ & ~new_new_n1616__;
  assign new_new_n1619__ = ~new_new_n1617__ & ~new_new_n1618__;
  assign new_new_n1620__ = ~new_new_n1570__ & new_new_n1619__;
  assign new_new_n1621__ = new_new_n1570__ & ~new_new_n1619__;
  assign new_new_n1622__ = ~new_new_n1620__ & ~new_new_n1621__;
  assign new_new_n1623__ = ~new_new_n1569__ & new_new_n1622__;
  assign new_new_n1624__ = new_new_n1569__ & ~new_new_n1622__;
  assign new_new_n1625__ = ~new_new_n1623__ & ~new_new_n1624__;
  assign new_new_n1626__ = ~new_new_n1568__ & new_new_n1625__;
  assign new_new_n1627__ = new_new_n1568__ & ~new_new_n1625__;
  assign new_new_n1628__ = ~new_new_n1626__ & ~new_new_n1627__;
  assign new_new_n1629__ = ~new_new_n1567__ & new_new_n1628__;
  assign new_new_n1630__ = new_new_n1567__ & ~new_new_n1628__;
  assign new_new_n1631__ = ~new_new_n1629__ & ~new_new_n1630__;
  assign new_new_n1632__ = ~new_new_n1566__ & new_new_n1631__;
  assign new_new_n1633__ = new_new_n1566__ & ~new_new_n1631__;
  assign new_new_n1634__ = ~new_new_n1632__ & ~new_new_n1633__;
  assign new_new_n1635__ = ~new_new_n1565__ & new_new_n1634__;
  assign new_new_n1636__ = new_new_n1565__ & ~new_new_n1634__;
  assign G6210gat = new_new_n1635__ | new_new_n1636__;
  assign new_new_n1638__ = ~new_new_n1632__ & ~new_new_n1635__;
  assign new_new_n1639__ = ~new_new_n1626__ & ~new_new_n1629__;
  assign new_new_n1640__ = G137gat & G528gat;
  assign new_new_n1641__ = ~new_new_n1620__ & ~new_new_n1623__;
  assign new_new_n1642__ = G154gat & G511gat;
  assign new_new_n1643__ = ~new_new_n1614__ & ~new_new_n1617__;
  assign new_new_n1644__ = G171gat & G494gat;
  assign new_new_n1645__ = ~new_new_n1608__ & ~new_new_n1611__;
  assign new_new_n1646__ = G188gat & G477gat;
  assign new_new_n1647__ = ~new_new_n1602__ & ~new_new_n1605__;
  assign new_new_n1648__ = G205gat & G460gat;
  assign new_new_n1649__ = ~new_new_n1596__ & ~new_new_n1599__;
  assign new_new_n1650__ = G222gat & G443gat;
  assign new_new_n1651__ = ~new_new_n1590__ & ~new_new_n1593__;
  assign new_new_n1652__ = G239gat & G426gat;
  assign new_new_n1653__ = G256gat & G409gat;
  assign new_new_n1654__ = ~new_new_n1584__ & ~new_new_n1587__;
  assign new_new_n1655__ = ~new_new_n1653__ & ~new_new_n1654__;
  assign new_new_n1656__ = new_new_n1653__ & new_new_n1654__;
  assign new_new_n1657__ = ~new_new_n1655__ & ~new_new_n1656__;
  assign new_new_n1658__ = ~new_new_n1652__ & new_new_n1657__;
  assign new_new_n1659__ = new_new_n1652__ & ~new_new_n1657__;
  assign new_new_n1660__ = ~new_new_n1658__ & ~new_new_n1659__;
  assign new_new_n1661__ = ~new_new_n1651__ & new_new_n1660__;
  assign new_new_n1662__ = new_new_n1651__ & ~new_new_n1660__;
  assign new_new_n1663__ = ~new_new_n1661__ & ~new_new_n1662__;
  assign new_new_n1664__ = ~new_new_n1650__ & new_new_n1663__;
  assign new_new_n1665__ = new_new_n1650__ & ~new_new_n1663__;
  assign new_new_n1666__ = ~new_new_n1664__ & ~new_new_n1665__;
  assign new_new_n1667__ = ~new_new_n1649__ & new_new_n1666__;
  assign new_new_n1668__ = new_new_n1649__ & ~new_new_n1666__;
  assign new_new_n1669__ = ~new_new_n1667__ & ~new_new_n1668__;
  assign new_new_n1670__ = ~new_new_n1648__ & new_new_n1669__;
  assign new_new_n1671__ = new_new_n1648__ & ~new_new_n1669__;
  assign new_new_n1672__ = ~new_new_n1670__ & ~new_new_n1671__;
  assign new_new_n1673__ = ~new_new_n1647__ & new_new_n1672__;
  assign new_new_n1674__ = new_new_n1647__ & ~new_new_n1672__;
  assign new_new_n1675__ = ~new_new_n1673__ & ~new_new_n1674__;
  assign new_new_n1676__ = ~new_new_n1646__ & new_new_n1675__;
  assign new_new_n1677__ = new_new_n1646__ & ~new_new_n1675__;
  assign new_new_n1678__ = ~new_new_n1676__ & ~new_new_n1677__;
  assign new_new_n1679__ = ~new_new_n1645__ & new_new_n1678__;
  assign new_new_n1680__ = new_new_n1645__ & ~new_new_n1678__;
  assign new_new_n1681__ = ~new_new_n1679__ & ~new_new_n1680__;
  assign new_new_n1682__ = ~new_new_n1644__ & new_new_n1681__;
  assign new_new_n1683__ = new_new_n1644__ & ~new_new_n1681__;
  assign new_new_n1684__ = ~new_new_n1682__ & ~new_new_n1683__;
  assign new_new_n1685__ = ~new_new_n1643__ & new_new_n1684__;
  assign new_new_n1686__ = new_new_n1643__ & ~new_new_n1684__;
  assign new_new_n1687__ = ~new_new_n1685__ & ~new_new_n1686__;
  assign new_new_n1688__ = ~new_new_n1642__ & new_new_n1687__;
  assign new_new_n1689__ = new_new_n1642__ & ~new_new_n1687__;
  assign new_new_n1690__ = ~new_new_n1688__ & ~new_new_n1689__;
  assign new_new_n1691__ = ~new_new_n1641__ & new_new_n1690__;
  assign new_new_n1692__ = new_new_n1641__ & ~new_new_n1690__;
  assign new_new_n1693__ = ~new_new_n1691__ & ~new_new_n1692__;
  assign new_new_n1694__ = ~new_new_n1640__ & new_new_n1693__;
  assign new_new_n1695__ = new_new_n1640__ & ~new_new_n1693__;
  assign new_new_n1696__ = ~new_new_n1694__ & ~new_new_n1695__;
  assign new_new_n1697__ = ~new_new_n1639__ & new_new_n1696__;
  assign new_new_n1698__ = new_new_n1639__ & ~new_new_n1696__;
  assign new_new_n1699__ = ~new_new_n1697__ & ~new_new_n1698__;
  assign new_new_n1700__ = ~new_new_n1638__ & new_new_n1699__;
  assign new_new_n1701__ = new_new_n1638__ & ~new_new_n1699__;
  assign G6220gat = new_new_n1700__ | new_new_n1701__;
  assign new_new_n1703__ = ~new_new_n1697__ & ~new_new_n1700__;
  assign new_new_n1704__ = ~new_new_n1691__ & ~new_new_n1694__;
  assign new_new_n1705__ = G154gat & G528gat;
  assign new_new_n1706__ = ~new_new_n1685__ & ~new_new_n1688__;
  assign new_new_n1707__ = G171gat & G511gat;
  assign new_new_n1708__ = ~new_new_n1679__ & ~new_new_n1682__;
  assign new_new_n1709__ = G188gat & G494gat;
  assign new_new_n1710__ = ~new_new_n1673__ & ~new_new_n1676__;
  assign new_new_n1711__ = G205gat & G477gat;
  assign new_new_n1712__ = ~new_new_n1667__ & ~new_new_n1670__;
  assign new_new_n1713__ = G222gat & G460gat;
  assign new_new_n1714__ = ~new_new_n1661__ & ~new_new_n1664__;
  assign new_new_n1715__ = G239gat & G443gat;
  assign new_new_n1716__ = G256gat & G426gat;
  assign new_new_n1717__ = ~new_new_n1655__ & ~new_new_n1658__;
  assign new_new_n1718__ = ~new_new_n1716__ & ~new_new_n1717__;
  assign new_new_n1719__ = new_new_n1716__ & new_new_n1717__;
  assign new_new_n1720__ = ~new_new_n1718__ & ~new_new_n1719__;
  assign new_new_n1721__ = ~new_new_n1715__ & new_new_n1720__;
  assign new_new_n1722__ = new_new_n1715__ & ~new_new_n1720__;
  assign new_new_n1723__ = ~new_new_n1721__ & ~new_new_n1722__;
  assign new_new_n1724__ = ~new_new_n1714__ & new_new_n1723__;
  assign new_new_n1725__ = new_new_n1714__ & ~new_new_n1723__;
  assign new_new_n1726__ = ~new_new_n1724__ & ~new_new_n1725__;
  assign new_new_n1727__ = ~new_new_n1713__ & new_new_n1726__;
  assign new_new_n1728__ = new_new_n1713__ & ~new_new_n1726__;
  assign new_new_n1729__ = ~new_new_n1727__ & ~new_new_n1728__;
  assign new_new_n1730__ = ~new_new_n1712__ & new_new_n1729__;
  assign new_new_n1731__ = new_new_n1712__ & ~new_new_n1729__;
  assign new_new_n1732__ = ~new_new_n1730__ & ~new_new_n1731__;
  assign new_new_n1733__ = ~new_new_n1711__ & new_new_n1732__;
  assign new_new_n1734__ = new_new_n1711__ & ~new_new_n1732__;
  assign new_new_n1735__ = ~new_new_n1733__ & ~new_new_n1734__;
  assign new_new_n1736__ = ~new_new_n1710__ & new_new_n1735__;
  assign new_new_n1737__ = new_new_n1710__ & ~new_new_n1735__;
  assign new_new_n1738__ = ~new_new_n1736__ & ~new_new_n1737__;
  assign new_new_n1739__ = ~new_new_n1709__ & new_new_n1738__;
  assign new_new_n1740__ = new_new_n1709__ & ~new_new_n1738__;
  assign new_new_n1741__ = ~new_new_n1739__ & ~new_new_n1740__;
  assign new_new_n1742__ = ~new_new_n1708__ & new_new_n1741__;
  assign new_new_n1743__ = new_new_n1708__ & ~new_new_n1741__;
  assign new_new_n1744__ = ~new_new_n1742__ & ~new_new_n1743__;
  assign new_new_n1745__ = ~new_new_n1707__ & new_new_n1744__;
  assign new_new_n1746__ = new_new_n1707__ & ~new_new_n1744__;
  assign new_new_n1747__ = ~new_new_n1745__ & ~new_new_n1746__;
  assign new_new_n1748__ = ~new_new_n1706__ & new_new_n1747__;
  assign new_new_n1749__ = new_new_n1706__ & ~new_new_n1747__;
  assign new_new_n1750__ = ~new_new_n1748__ & ~new_new_n1749__;
  assign new_new_n1751__ = ~new_new_n1705__ & new_new_n1750__;
  assign new_new_n1752__ = new_new_n1705__ & ~new_new_n1750__;
  assign new_new_n1753__ = ~new_new_n1751__ & ~new_new_n1752__;
  assign new_new_n1754__ = ~new_new_n1704__ & new_new_n1753__;
  assign new_new_n1755__ = new_new_n1704__ & ~new_new_n1753__;
  assign new_new_n1756__ = ~new_new_n1754__ & ~new_new_n1755__;
  assign new_new_n1757__ = ~new_new_n1703__ & new_new_n1756__;
  assign new_new_n1758__ = new_new_n1703__ & ~new_new_n1756__;
  assign G6230gat = new_new_n1757__ | new_new_n1758__;
  assign new_new_n1760__ = ~new_new_n1754__ & ~new_new_n1757__;
  assign new_new_n1761__ = ~new_new_n1748__ & ~new_new_n1751__;
  assign new_new_n1762__ = G171gat & G528gat;
  assign new_new_n1763__ = ~new_new_n1742__ & ~new_new_n1745__;
  assign new_new_n1764__ = G188gat & G511gat;
  assign new_new_n1765__ = ~new_new_n1736__ & ~new_new_n1739__;
  assign new_new_n1766__ = G205gat & G494gat;
  assign new_new_n1767__ = ~new_new_n1730__ & ~new_new_n1733__;
  assign new_new_n1768__ = G222gat & G477gat;
  assign new_new_n1769__ = ~new_new_n1724__ & ~new_new_n1727__;
  assign new_new_n1770__ = G239gat & G460gat;
  assign new_new_n1771__ = G256gat & G443gat;
  assign new_new_n1772__ = ~new_new_n1718__ & ~new_new_n1721__;
  assign new_new_n1773__ = ~new_new_n1771__ & ~new_new_n1772__;
  assign new_new_n1774__ = new_new_n1771__ & new_new_n1772__;
  assign new_new_n1775__ = ~new_new_n1773__ & ~new_new_n1774__;
  assign new_new_n1776__ = ~new_new_n1770__ & new_new_n1775__;
  assign new_new_n1777__ = new_new_n1770__ & ~new_new_n1775__;
  assign new_new_n1778__ = ~new_new_n1776__ & ~new_new_n1777__;
  assign new_new_n1779__ = ~new_new_n1769__ & new_new_n1778__;
  assign new_new_n1780__ = new_new_n1769__ & ~new_new_n1778__;
  assign new_new_n1781__ = ~new_new_n1779__ & ~new_new_n1780__;
  assign new_new_n1782__ = ~new_new_n1768__ & new_new_n1781__;
  assign new_new_n1783__ = new_new_n1768__ & ~new_new_n1781__;
  assign new_new_n1784__ = ~new_new_n1782__ & ~new_new_n1783__;
  assign new_new_n1785__ = ~new_new_n1767__ & new_new_n1784__;
  assign new_new_n1786__ = new_new_n1767__ & ~new_new_n1784__;
  assign new_new_n1787__ = ~new_new_n1785__ & ~new_new_n1786__;
  assign new_new_n1788__ = ~new_new_n1766__ & new_new_n1787__;
  assign new_new_n1789__ = new_new_n1766__ & ~new_new_n1787__;
  assign new_new_n1790__ = ~new_new_n1788__ & ~new_new_n1789__;
  assign new_new_n1791__ = ~new_new_n1765__ & new_new_n1790__;
  assign new_new_n1792__ = new_new_n1765__ & ~new_new_n1790__;
  assign new_new_n1793__ = ~new_new_n1791__ & ~new_new_n1792__;
  assign new_new_n1794__ = ~new_new_n1764__ & new_new_n1793__;
  assign new_new_n1795__ = new_new_n1764__ & ~new_new_n1793__;
  assign new_new_n1796__ = ~new_new_n1794__ & ~new_new_n1795__;
  assign new_new_n1797__ = ~new_new_n1763__ & new_new_n1796__;
  assign new_new_n1798__ = new_new_n1763__ & ~new_new_n1796__;
  assign new_new_n1799__ = ~new_new_n1797__ & ~new_new_n1798__;
  assign new_new_n1800__ = ~new_new_n1762__ & new_new_n1799__;
  assign new_new_n1801__ = new_new_n1762__ & ~new_new_n1799__;
  assign new_new_n1802__ = ~new_new_n1800__ & ~new_new_n1801__;
  assign new_new_n1803__ = ~new_new_n1761__ & new_new_n1802__;
  assign new_new_n1804__ = new_new_n1761__ & ~new_new_n1802__;
  assign new_new_n1805__ = ~new_new_n1803__ & ~new_new_n1804__;
  assign new_new_n1806__ = ~new_new_n1760__ & new_new_n1805__;
  assign new_new_n1807__ = new_new_n1760__ & ~new_new_n1805__;
  assign G6240gat = new_new_n1806__ | new_new_n1807__;
  assign new_new_n1809__ = ~new_new_n1803__ & ~new_new_n1806__;
  assign new_new_n1810__ = ~new_new_n1797__ & ~new_new_n1800__;
  assign new_new_n1811__ = G188gat & G528gat;
  assign new_new_n1812__ = ~new_new_n1791__ & ~new_new_n1794__;
  assign new_new_n1813__ = G205gat & G511gat;
  assign new_new_n1814__ = ~new_new_n1785__ & ~new_new_n1788__;
  assign new_new_n1815__ = G222gat & G494gat;
  assign new_new_n1816__ = ~new_new_n1779__ & ~new_new_n1782__;
  assign new_new_n1817__ = G239gat & G477gat;
  assign new_new_n1818__ = G256gat & G460gat;
  assign new_new_n1819__ = ~new_new_n1773__ & ~new_new_n1776__;
  assign new_new_n1820__ = ~new_new_n1818__ & ~new_new_n1819__;
  assign new_new_n1821__ = new_new_n1818__ & new_new_n1819__;
  assign new_new_n1822__ = ~new_new_n1820__ & ~new_new_n1821__;
  assign new_new_n1823__ = ~new_new_n1817__ & new_new_n1822__;
  assign new_new_n1824__ = new_new_n1817__ & ~new_new_n1822__;
  assign new_new_n1825__ = ~new_new_n1823__ & ~new_new_n1824__;
  assign new_new_n1826__ = ~new_new_n1816__ & new_new_n1825__;
  assign new_new_n1827__ = new_new_n1816__ & ~new_new_n1825__;
  assign new_new_n1828__ = ~new_new_n1826__ & ~new_new_n1827__;
  assign new_new_n1829__ = ~new_new_n1815__ & new_new_n1828__;
  assign new_new_n1830__ = new_new_n1815__ & ~new_new_n1828__;
  assign new_new_n1831__ = ~new_new_n1829__ & ~new_new_n1830__;
  assign new_new_n1832__ = ~new_new_n1814__ & new_new_n1831__;
  assign new_new_n1833__ = new_new_n1814__ & ~new_new_n1831__;
  assign new_new_n1834__ = ~new_new_n1832__ & ~new_new_n1833__;
  assign new_new_n1835__ = ~new_new_n1813__ & new_new_n1834__;
  assign new_new_n1836__ = new_new_n1813__ & ~new_new_n1834__;
  assign new_new_n1837__ = ~new_new_n1835__ & ~new_new_n1836__;
  assign new_new_n1838__ = ~new_new_n1812__ & new_new_n1837__;
  assign new_new_n1839__ = new_new_n1812__ & ~new_new_n1837__;
  assign new_new_n1840__ = ~new_new_n1838__ & ~new_new_n1839__;
  assign new_new_n1841__ = ~new_new_n1811__ & new_new_n1840__;
  assign new_new_n1842__ = new_new_n1811__ & ~new_new_n1840__;
  assign new_new_n1843__ = ~new_new_n1841__ & ~new_new_n1842__;
  assign new_new_n1844__ = ~new_new_n1810__ & new_new_n1843__;
  assign new_new_n1845__ = new_new_n1810__ & ~new_new_n1843__;
  assign new_new_n1846__ = ~new_new_n1844__ & ~new_new_n1845__;
  assign new_new_n1847__ = ~new_new_n1809__ & new_new_n1846__;
  assign new_new_n1848__ = new_new_n1809__ & ~new_new_n1846__;
  assign G6250gat = new_new_n1847__ | new_new_n1848__;
  assign new_new_n1850__ = ~new_new_n1844__ & ~new_new_n1847__;
  assign new_new_n1851__ = ~new_new_n1838__ & ~new_new_n1841__;
  assign new_new_n1852__ = G205gat & G528gat;
  assign new_new_n1853__ = ~new_new_n1832__ & ~new_new_n1835__;
  assign new_new_n1854__ = G222gat & G511gat;
  assign new_new_n1855__ = ~new_new_n1826__ & ~new_new_n1829__;
  assign new_new_n1856__ = G239gat & G494gat;
  assign new_new_n1857__ = G256gat & G477gat;
  assign new_new_n1858__ = ~new_new_n1820__ & ~new_new_n1823__;
  assign new_new_n1859__ = ~new_new_n1857__ & ~new_new_n1858__;
  assign new_new_n1860__ = new_new_n1857__ & new_new_n1858__;
  assign new_new_n1861__ = ~new_new_n1859__ & ~new_new_n1860__;
  assign new_new_n1862__ = ~new_new_n1856__ & new_new_n1861__;
  assign new_new_n1863__ = new_new_n1856__ & ~new_new_n1861__;
  assign new_new_n1864__ = ~new_new_n1862__ & ~new_new_n1863__;
  assign new_new_n1865__ = ~new_new_n1855__ & new_new_n1864__;
  assign new_new_n1866__ = new_new_n1855__ & ~new_new_n1864__;
  assign new_new_n1867__ = ~new_new_n1865__ & ~new_new_n1866__;
  assign new_new_n1868__ = ~new_new_n1854__ & new_new_n1867__;
  assign new_new_n1869__ = new_new_n1854__ & ~new_new_n1867__;
  assign new_new_n1870__ = ~new_new_n1868__ & ~new_new_n1869__;
  assign new_new_n1871__ = ~new_new_n1853__ & new_new_n1870__;
  assign new_new_n1872__ = new_new_n1853__ & ~new_new_n1870__;
  assign new_new_n1873__ = ~new_new_n1871__ & ~new_new_n1872__;
  assign new_new_n1874__ = ~new_new_n1852__ & new_new_n1873__;
  assign new_new_n1875__ = new_new_n1852__ & ~new_new_n1873__;
  assign new_new_n1876__ = ~new_new_n1874__ & ~new_new_n1875__;
  assign new_new_n1877__ = ~new_new_n1851__ & new_new_n1876__;
  assign new_new_n1878__ = new_new_n1851__ & ~new_new_n1876__;
  assign new_new_n1879__ = ~new_new_n1877__ & ~new_new_n1878__;
  assign new_new_n1880__ = ~new_new_n1850__ & new_new_n1879__;
  assign new_new_n1881__ = new_new_n1850__ & ~new_new_n1879__;
  assign G6260gat = new_new_n1880__ | new_new_n1881__;
  assign new_new_n1883__ = ~new_new_n1877__ & ~new_new_n1880__;
  assign new_new_n1884__ = ~new_new_n1871__ & ~new_new_n1874__;
  assign new_new_n1885__ = G222gat & G528gat;
  assign new_new_n1886__ = ~new_new_n1865__ & ~new_new_n1868__;
  assign new_new_n1887__ = G239gat & G511gat;
  assign new_new_n1888__ = G256gat & G494gat;
  assign new_new_n1889__ = ~new_new_n1859__ & ~new_new_n1862__;
  assign new_new_n1890__ = ~new_new_n1888__ & ~new_new_n1889__;
  assign new_new_n1891__ = new_new_n1888__ & new_new_n1889__;
  assign new_new_n1892__ = ~new_new_n1890__ & ~new_new_n1891__;
  assign new_new_n1893__ = ~new_new_n1887__ & new_new_n1892__;
  assign new_new_n1894__ = new_new_n1887__ & ~new_new_n1892__;
  assign new_new_n1895__ = ~new_new_n1893__ & ~new_new_n1894__;
  assign new_new_n1896__ = ~new_new_n1886__ & new_new_n1895__;
  assign new_new_n1897__ = new_new_n1886__ & ~new_new_n1895__;
  assign new_new_n1898__ = ~new_new_n1896__ & ~new_new_n1897__;
  assign new_new_n1899__ = ~new_new_n1885__ & new_new_n1898__;
  assign new_new_n1900__ = new_new_n1885__ & ~new_new_n1898__;
  assign new_new_n1901__ = ~new_new_n1899__ & ~new_new_n1900__;
  assign new_new_n1902__ = ~new_new_n1884__ & new_new_n1901__;
  assign new_new_n1903__ = new_new_n1884__ & ~new_new_n1901__;
  assign new_new_n1904__ = ~new_new_n1902__ & ~new_new_n1903__;
  assign new_new_n1905__ = ~new_new_n1883__ & new_new_n1904__;
  assign new_new_n1906__ = new_new_n1883__ & ~new_new_n1904__;
  assign G6270gat = new_new_n1905__ | new_new_n1906__;
  assign new_new_n1908__ = ~new_new_n1902__ & ~new_new_n1905__;
  assign new_new_n1909__ = ~new_new_n1896__ & ~new_new_n1899__;
  assign new_new_n1910__ = G239gat & G528gat;
  assign new_new_n1911__ = G256gat & G511gat;
  assign new_new_n1912__ = ~new_new_n1890__ & ~new_new_n1893__;
  assign new_new_n1913__ = ~new_new_n1911__ & ~new_new_n1912__;
  assign new_new_n1914__ = new_new_n1911__ & new_new_n1912__;
  assign new_new_n1915__ = ~new_new_n1913__ & ~new_new_n1914__;
  assign new_new_n1916__ = ~new_new_n1910__ & new_new_n1915__;
  assign new_new_n1917__ = new_new_n1910__ & ~new_new_n1915__;
  assign new_new_n1918__ = ~new_new_n1916__ & ~new_new_n1917__;
  assign new_new_n1919__ = ~new_new_n1909__ & new_new_n1918__;
  assign new_new_n1920__ = new_new_n1909__ & ~new_new_n1918__;
  assign new_new_n1921__ = ~new_new_n1919__ & ~new_new_n1920__;
  assign new_new_n1922__ = ~new_new_n1908__ & new_new_n1921__;
  assign new_new_n1923__ = new_new_n1908__ & ~new_new_n1921__;
  assign G6280gat = new_new_n1922__ | new_new_n1923__;
  assign new_new_n1925__ = G256gat & G528gat;
  assign new_new_n1926__ = ~new_new_n1913__ & ~new_new_n1916__;
  assign new_new_n1927__ = ~new_new_n1925__ & ~new_new_n1926__;
  assign new_new_n1928__ = ~new_new_n1919__ & ~new_new_n1922__;
  assign new_new_n1929__ = new_new_n1925__ & new_new_n1926__;
  assign new_new_n1930__ = ~new_new_n1927__ & ~new_new_n1929__;
  assign new_new_n1931__ = ~new_new_n1928__ & new_new_n1930__;
  assign G6287gat = ~new_new_n1927__ & ~new_new_n1931__;
  assign new_new_n1933__ = new_new_n1928__ & ~new_new_n1930__;
  assign G6288gat = new_new_n1931__ | new_new_n1933__;
endmodule


