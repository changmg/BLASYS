module max_3_2_tb;
reg [9:0] pi;
wire [4:0] po;
max_3_2 dut(pi[9], pi[8], pi[7], pi[6], pi[5], pi[4], pi[3], pi[2], pi[1], pi[0], po[4], po[3], po[2], po[1], po[0]);
initial
begin
# 1  pi=10'b0000000000;
#1 $display("%b", po);
# 1  pi=10'b0000000001;
#1 $display("%b", po);
# 1  pi=10'b0000000010;
#1 $display("%b", po);
# 1  pi=10'b0000000011;
#1 $display("%b", po);
# 1  pi=10'b0000000100;
#1 $display("%b", po);
# 1  pi=10'b0000000101;
#1 $display("%b", po);
# 1  pi=10'b0000000110;
#1 $display("%b", po);
# 1  pi=10'b0000000111;
#1 $display("%b", po);
# 1  pi=10'b0000001000;
#1 $display("%b", po);
# 1  pi=10'b0000001001;
#1 $display("%b", po);
# 1  pi=10'b0000001010;
#1 $display("%b", po);
# 1  pi=10'b0000001011;
#1 $display("%b", po);
# 1  pi=10'b0000001100;
#1 $display("%b", po);
# 1  pi=10'b0000001101;
#1 $display("%b", po);
# 1  pi=10'b0000001110;
#1 $display("%b", po);
# 1  pi=10'b0000001111;
#1 $display("%b", po);
# 1  pi=10'b0000010000;
#1 $display("%b", po);
# 1  pi=10'b0000010001;
#1 $display("%b", po);
# 1  pi=10'b0000010010;
#1 $display("%b", po);
# 1  pi=10'b0000010011;
#1 $display("%b", po);
# 1  pi=10'b0000010100;
#1 $display("%b", po);
# 1  pi=10'b0000010101;
#1 $display("%b", po);
# 1  pi=10'b0000010110;
#1 $display("%b", po);
# 1  pi=10'b0000010111;
#1 $display("%b", po);
# 1  pi=10'b0000011000;
#1 $display("%b", po);
# 1  pi=10'b0000011001;
#1 $display("%b", po);
# 1  pi=10'b0000011010;
#1 $display("%b", po);
# 1  pi=10'b0000011011;
#1 $display("%b", po);
# 1  pi=10'b0000011100;
#1 $display("%b", po);
# 1  pi=10'b0000011101;
#1 $display("%b", po);
# 1  pi=10'b0000011110;
#1 $display("%b", po);
# 1  pi=10'b0000011111;
#1 $display("%b", po);
# 1  pi=10'b0000100000;
#1 $display("%b", po);
# 1  pi=10'b0000100001;
#1 $display("%b", po);
# 1  pi=10'b0000100010;
#1 $display("%b", po);
# 1  pi=10'b0000100011;
#1 $display("%b", po);
# 1  pi=10'b0000100100;
#1 $display("%b", po);
# 1  pi=10'b0000100101;
#1 $display("%b", po);
# 1  pi=10'b0000100110;
#1 $display("%b", po);
# 1  pi=10'b0000100111;
#1 $display("%b", po);
# 1  pi=10'b0000101000;
#1 $display("%b", po);
# 1  pi=10'b0000101001;
#1 $display("%b", po);
# 1  pi=10'b0000101010;
#1 $display("%b", po);
# 1  pi=10'b0000101011;
#1 $display("%b", po);
# 1  pi=10'b0000101100;
#1 $display("%b", po);
# 1  pi=10'b0000101101;
#1 $display("%b", po);
# 1  pi=10'b0000101110;
#1 $display("%b", po);
# 1  pi=10'b0000101111;
#1 $display("%b", po);
# 1  pi=10'b0000110000;
#1 $display("%b", po);
# 1  pi=10'b0000110001;
#1 $display("%b", po);
# 1  pi=10'b0000110010;
#1 $display("%b", po);
# 1  pi=10'b0000110011;
#1 $display("%b", po);
# 1  pi=10'b0000110100;
#1 $display("%b", po);
# 1  pi=10'b0000110101;
#1 $display("%b", po);
# 1  pi=10'b0000110110;
#1 $display("%b", po);
# 1  pi=10'b0000110111;
#1 $display("%b", po);
# 1  pi=10'b0000111000;
#1 $display("%b", po);
# 1  pi=10'b0000111001;
#1 $display("%b", po);
# 1  pi=10'b0000111010;
#1 $display("%b", po);
# 1  pi=10'b0000111011;
#1 $display("%b", po);
# 1  pi=10'b0000111100;
#1 $display("%b", po);
# 1  pi=10'b0000111101;
#1 $display("%b", po);
# 1  pi=10'b0000111110;
#1 $display("%b", po);
# 1  pi=10'b0000111111;
#1 $display("%b", po);
# 1  pi=10'b0001000000;
#1 $display("%b", po);
# 1  pi=10'b0001000001;
#1 $display("%b", po);
# 1  pi=10'b0001000010;
#1 $display("%b", po);
# 1  pi=10'b0001000011;
#1 $display("%b", po);
# 1  pi=10'b0001000100;
#1 $display("%b", po);
# 1  pi=10'b0001000101;
#1 $display("%b", po);
# 1  pi=10'b0001000110;
#1 $display("%b", po);
# 1  pi=10'b0001000111;
#1 $display("%b", po);
# 1  pi=10'b0001001000;
#1 $display("%b", po);
# 1  pi=10'b0001001001;
#1 $display("%b", po);
# 1  pi=10'b0001001010;
#1 $display("%b", po);
# 1  pi=10'b0001001011;
#1 $display("%b", po);
# 1  pi=10'b0001001100;
#1 $display("%b", po);
# 1  pi=10'b0001001101;
#1 $display("%b", po);
# 1  pi=10'b0001001110;
#1 $display("%b", po);
# 1  pi=10'b0001001111;
#1 $display("%b", po);
# 1  pi=10'b0001010000;
#1 $display("%b", po);
# 1  pi=10'b0001010001;
#1 $display("%b", po);
# 1  pi=10'b0001010010;
#1 $display("%b", po);
# 1  pi=10'b0001010011;
#1 $display("%b", po);
# 1  pi=10'b0001010100;
#1 $display("%b", po);
# 1  pi=10'b0001010101;
#1 $display("%b", po);
# 1  pi=10'b0001010110;
#1 $display("%b", po);
# 1  pi=10'b0001010111;
#1 $display("%b", po);
# 1  pi=10'b0001011000;
#1 $display("%b", po);
# 1  pi=10'b0001011001;
#1 $display("%b", po);
# 1  pi=10'b0001011010;
#1 $display("%b", po);
# 1  pi=10'b0001011011;
#1 $display("%b", po);
# 1  pi=10'b0001011100;
#1 $display("%b", po);
# 1  pi=10'b0001011101;
#1 $display("%b", po);
# 1  pi=10'b0001011110;
#1 $display("%b", po);
# 1  pi=10'b0001011111;
#1 $display("%b", po);
# 1  pi=10'b0001100000;
#1 $display("%b", po);
# 1  pi=10'b0001100001;
#1 $display("%b", po);
# 1  pi=10'b0001100010;
#1 $display("%b", po);
# 1  pi=10'b0001100011;
#1 $display("%b", po);
# 1  pi=10'b0001100100;
#1 $display("%b", po);
# 1  pi=10'b0001100101;
#1 $display("%b", po);
# 1  pi=10'b0001100110;
#1 $display("%b", po);
# 1  pi=10'b0001100111;
#1 $display("%b", po);
# 1  pi=10'b0001101000;
#1 $display("%b", po);
# 1  pi=10'b0001101001;
#1 $display("%b", po);
# 1  pi=10'b0001101010;
#1 $display("%b", po);
# 1  pi=10'b0001101011;
#1 $display("%b", po);
# 1  pi=10'b0001101100;
#1 $display("%b", po);
# 1  pi=10'b0001101101;
#1 $display("%b", po);
# 1  pi=10'b0001101110;
#1 $display("%b", po);
# 1  pi=10'b0001101111;
#1 $display("%b", po);
# 1  pi=10'b0001110000;
#1 $display("%b", po);
# 1  pi=10'b0001110001;
#1 $display("%b", po);
# 1  pi=10'b0001110010;
#1 $display("%b", po);
# 1  pi=10'b0001110011;
#1 $display("%b", po);
# 1  pi=10'b0001110100;
#1 $display("%b", po);
# 1  pi=10'b0001110101;
#1 $display("%b", po);
# 1  pi=10'b0001110110;
#1 $display("%b", po);
# 1  pi=10'b0001110111;
#1 $display("%b", po);
# 1  pi=10'b0001111000;
#1 $display("%b", po);
# 1  pi=10'b0001111001;
#1 $display("%b", po);
# 1  pi=10'b0001111010;
#1 $display("%b", po);
# 1  pi=10'b0001111011;
#1 $display("%b", po);
# 1  pi=10'b0001111100;
#1 $display("%b", po);
# 1  pi=10'b0001111101;
#1 $display("%b", po);
# 1  pi=10'b0001111110;
#1 $display("%b", po);
# 1  pi=10'b0001111111;
#1 $display("%b", po);
# 1  pi=10'b0010000000;
#1 $display("%b", po);
# 1  pi=10'b0010000001;
#1 $display("%b", po);
# 1  pi=10'b0010000010;
#1 $display("%b", po);
# 1  pi=10'b0010000011;
#1 $display("%b", po);
# 1  pi=10'b0010000100;
#1 $display("%b", po);
# 1  pi=10'b0010000101;
#1 $display("%b", po);
# 1  pi=10'b0010000110;
#1 $display("%b", po);
# 1  pi=10'b0010000111;
#1 $display("%b", po);
# 1  pi=10'b0010001000;
#1 $display("%b", po);
# 1  pi=10'b0010001001;
#1 $display("%b", po);
# 1  pi=10'b0010001010;
#1 $display("%b", po);
# 1  pi=10'b0010001011;
#1 $display("%b", po);
# 1  pi=10'b0010001100;
#1 $display("%b", po);
# 1  pi=10'b0010001101;
#1 $display("%b", po);
# 1  pi=10'b0010001110;
#1 $display("%b", po);
# 1  pi=10'b0010001111;
#1 $display("%b", po);
# 1  pi=10'b0010010000;
#1 $display("%b", po);
# 1  pi=10'b0010010001;
#1 $display("%b", po);
# 1  pi=10'b0010010010;
#1 $display("%b", po);
# 1  pi=10'b0010010011;
#1 $display("%b", po);
# 1  pi=10'b0010010100;
#1 $display("%b", po);
# 1  pi=10'b0010010101;
#1 $display("%b", po);
# 1  pi=10'b0010010110;
#1 $display("%b", po);
# 1  pi=10'b0010010111;
#1 $display("%b", po);
# 1  pi=10'b0010011000;
#1 $display("%b", po);
# 1  pi=10'b0010011001;
#1 $display("%b", po);
# 1  pi=10'b0010011010;
#1 $display("%b", po);
# 1  pi=10'b0010011011;
#1 $display("%b", po);
# 1  pi=10'b0010011100;
#1 $display("%b", po);
# 1  pi=10'b0010011101;
#1 $display("%b", po);
# 1  pi=10'b0010011110;
#1 $display("%b", po);
# 1  pi=10'b0010011111;
#1 $display("%b", po);
# 1  pi=10'b0010100000;
#1 $display("%b", po);
# 1  pi=10'b0010100001;
#1 $display("%b", po);
# 1  pi=10'b0010100010;
#1 $display("%b", po);
# 1  pi=10'b0010100011;
#1 $display("%b", po);
# 1  pi=10'b0010100100;
#1 $display("%b", po);
# 1  pi=10'b0010100101;
#1 $display("%b", po);
# 1  pi=10'b0010100110;
#1 $display("%b", po);
# 1  pi=10'b0010100111;
#1 $display("%b", po);
# 1  pi=10'b0010101000;
#1 $display("%b", po);
# 1  pi=10'b0010101001;
#1 $display("%b", po);
# 1  pi=10'b0010101010;
#1 $display("%b", po);
# 1  pi=10'b0010101011;
#1 $display("%b", po);
# 1  pi=10'b0010101100;
#1 $display("%b", po);
# 1  pi=10'b0010101101;
#1 $display("%b", po);
# 1  pi=10'b0010101110;
#1 $display("%b", po);
# 1  pi=10'b0010101111;
#1 $display("%b", po);
# 1  pi=10'b0010110000;
#1 $display("%b", po);
# 1  pi=10'b0010110001;
#1 $display("%b", po);
# 1  pi=10'b0010110010;
#1 $display("%b", po);
# 1  pi=10'b0010110011;
#1 $display("%b", po);
# 1  pi=10'b0010110100;
#1 $display("%b", po);
# 1  pi=10'b0010110101;
#1 $display("%b", po);
# 1  pi=10'b0010110110;
#1 $display("%b", po);
# 1  pi=10'b0010110111;
#1 $display("%b", po);
# 1  pi=10'b0010111000;
#1 $display("%b", po);
# 1  pi=10'b0010111001;
#1 $display("%b", po);
# 1  pi=10'b0010111010;
#1 $display("%b", po);
# 1  pi=10'b0010111011;
#1 $display("%b", po);
# 1  pi=10'b0010111100;
#1 $display("%b", po);
# 1  pi=10'b0010111101;
#1 $display("%b", po);
# 1  pi=10'b0010111110;
#1 $display("%b", po);
# 1  pi=10'b0010111111;
#1 $display("%b", po);
# 1  pi=10'b0011000000;
#1 $display("%b", po);
# 1  pi=10'b0011000001;
#1 $display("%b", po);
# 1  pi=10'b0011000010;
#1 $display("%b", po);
# 1  pi=10'b0011000011;
#1 $display("%b", po);
# 1  pi=10'b0011000100;
#1 $display("%b", po);
# 1  pi=10'b0011000101;
#1 $display("%b", po);
# 1  pi=10'b0011000110;
#1 $display("%b", po);
# 1  pi=10'b0011000111;
#1 $display("%b", po);
# 1  pi=10'b0011001000;
#1 $display("%b", po);
# 1  pi=10'b0011001001;
#1 $display("%b", po);
# 1  pi=10'b0011001010;
#1 $display("%b", po);
# 1  pi=10'b0011001011;
#1 $display("%b", po);
# 1  pi=10'b0011001100;
#1 $display("%b", po);
# 1  pi=10'b0011001101;
#1 $display("%b", po);
# 1  pi=10'b0011001110;
#1 $display("%b", po);
# 1  pi=10'b0011001111;
#1 $display("%b", po);
# 1  pi=10'b0011010000;
#1 $display("%b", po);
# 1  pi=10'b0011010001;
#1 $display("%b", po);
# 1  pi=10'b0011010010;
#1 $display("%b", po);
# 1  pi=10'b0011010011;
#1 $display("%b", po);
# 1  pi=10'b0011010100;
#1 $display("%b", po);
# 1  pi=10'b0011010101;
#1 $display("%b", po);
# 1  pi=10'b0011010110;
#1 $display("%b", po);
# 1  pi=10'b0011010111;
#1 $display("%b", po);
# 1  pi=10'b0011011000;
#1 $display("%b", po);
# 1  pi=10'b0011011001;
#1 $display("%b", po);
# 1  pi=10'b0011011010;
#1 $display("%b", po);
# 1  pi=10'b0011011011;
#1 $display("%b", po);
# 1  pi=10'b0011011100;
#1 $display("%b", po);
# 1  pi=10'b0011011101;
#1 $display("%b", po);
# 1  pi=10'b0011011110;
#1 $display("%b", po);
# 1  pi=10'b0011011111;
#1 $display("%b", po);
# 1  pi=10'b0011100000;
#1 $display("%b", po);
# 1  pi=10'b0011100001;
#1 $display("%b", po);
# 1  pi=10'b0011100010;
#1 $display("%b", po);
# 1  pi=10'b0011100011;
#1 $display("%b", po);
# 1  pi=10'b0011100100;
#1 $display("%b", po);
# 1  pi=10'b0011100101;
#1 $display("%b", po);
# 1  pi=10'b0011100110;
#1 $display("%b", po);
# 1  pi=10'b0011100111;
#1 $display("%b", po);
# 1  pi=10'b0011101000;
#1 $display("%b", po);
# 1  pi=10'b0011101001;
#1 $display("%b", po);
# 1  pi=10'b0011101010;
#1 $display("%b", po);
# 1  pi=10'b0011101011;
#1 $display("%b", po);
# 1  pi=10'b0011101100;
#1 $display("%b", po);
# 1  pi=10'b0011101101;
#1 $display("%b", po);
# 1  pi=10'b0011101110;
#1 $display("%b", po);
# 1  pi=10'b0011101111;
#1 $display("%b", po);
# 1  pi=10'b0011110000;
#1 $display("%b", po);
# 1  pi=10'b0011110001;
#1 $display("%b", po);
# 1  pi=10'b0011110010;
#1 $display("%b", po);
# 1  pi=10'b0011110011;
#1 $display("%b", po);
# 1  pi=10'b0011110100;
#1 $display("%b", po);
# 1  pi=10'b0011110101;
#1 $display("%b", po);
# 1  pi=10'b0011110110;
#1 $display("%b", po);
# 1  pi=10'b0011110111;
#1 $display("%b", po);
# 1  pi=10'b0011111000;
#1 $display("%b", po);
# 1  pi=10'b0011111001;
#1 $display("%b", po);
# 1  pi=10'b0011111010;
#1 $display("%b", po);
# 1  pi=10'b0011111011;
#1 $display("%b", po);
# 1  pi=10'b0011111100;
#1 $display("%b", po);
# 1  pi=10'b0011111101;
#1 $display("%b", po);
# 1  pi=10'b0011111110;
#1 $display("%b", po);
# 1  pi=10'b0011111111;
#1 $display("%b", po);
# 1  pi=10'b0100000000;
#1 $display("%b", po);
# 1  pi=10'b0100000001;
#1 $display("%b", po);
# 1  pi=10'b0100000010;
#1 $display("%b", po);
# 1  pi=10'b0100000011;
#1 $display("%b", po);
# 1  pi=10'b0100000100;
#1 $display("%b", po);
# 1  pi=10'b0100000101;
#1 $display("%b", po);
# 1  pi=10'b0100000110;
#1 $display("%b", po);
# 1  pi=10'b0100000111;
#1 $display("%b", po);
# 1  pi=10'b0100001000;
#1 $display("%b", po);
# 1  pi=10'b0100001001;
#1 $display("%b", po);
# 1  pi=10'b0100001010;
#1 $display("%b", po);
# 1  pi=10'b0100001011;
#1 $display("%b", po);
# 1  pi=10'b0100001100;
#1 $display("%b", po);
# 1  pi=10'b0100001101;
#1 $display("%b", po);
# 1  pi=10'b0100001110;
#1 $display("%b", po);
# 1  pi=10'b0100001111;
#1 $display("%b", po);
# 1  pi=10'b0100010000;
#1 $display("%b", po);
# 1  pi=10'b0100010001;
#1 $display("%b", po);
# 1  pi=10'b0100010010;
#1 $display("%b", po);
# 1  pi=10'b0100010011;
#1 $display("%b", po);
# 1  pi=10'b0100010100;
#1 $display("%b", po);
# 1  pi=10'b0100010101;
#1 $display("%b", po);
# 1  pi=10'b0100010110;
#1 $display("%b", po);
# 1  pi=10'b0100010111;
#1 $display("%b", po);
# 1  pi=10'b0100011000;
#1 $display("%b", po);
# 1  pi=10'b0100011001;
#1 $display("%b", po);
# 1  pi=10'b0100011010;
#1 $display("%b", po);
# 1  pi=10'b0100011011;
#1 $display("%b", po);
# 1  pi=10'b0100011100;
#1 $display("%b", po);
# 1  pi=10'b0100011101;
#1 $display("%b", po);
# 1  pi=10'b0100011110;
#1 $display("%b", po);
# 1  pi=10'b0100011111;
#1 $display("%b", po);
# 1  pi=10'b0100100000;
#1 $display("%b", po);
# 1  pi=10'b0100100001;
#1 $display("%b", po);
# 1  pi=10'b0100100010;
#1 $display("%b", po);
# 1  pi=10'b0100100011;
#1 $display("%b", po);
# 1  pi=10'b0100100100;
#1 $display("%b", po);
# 1  pi=10'b0100100101;
#1 $display("%b", po);
# 1  pi=10'b0100100110;
#1 $display("%b", po);
# 1  pi=10'b0100100111;
#1 $display("%b", po);
# 1  pi=10'b0100101000;
#1 $display("%b", po);
# 1  pi=10'b0100101001;
#1 $display("%b", po);
# 1  pi=10'b0100101010;
#1 $display("%b", po);
# 1  pi=10'b0100101011;
#1 $display("%b", po);
# 1  pi=10'b0100101100;
#1 $display("%b", po);
# 1  pi=10'b0100101101;
#1 $display("%b", po);
# 1  pi=10'b0100101110;
#1 $display("%b", po);
# 1  pi=10'b0100101111;
#1 $display("%b", po);
# 1  pi=10'b0100110000;
#1 $display("%b", po);
# 1  pi=10'b0100110001;
#1 $display("%b", po);
# 1  pi=10'b0100110010;
#1 $display("%b", po);
# 1  pi=10'b0100110011;
#1 $display("%b", po);
# 1  pi=10'b0100110100;
#1 $display("%b", po);
# 1  pi=10'b0100110101;
#1 $display("%b", po);
# 1  pi=10'b0100110110;
#1 $display("%b", po);
# 1  pi=10'b0100110111;
#1 $display("%b", po);
# 1  pi=10'b0100111000;
#1 $display("%b", po);
# 1  pi=10'b0100111001;
#1 $display("%b", po);
# 1  pi=10'b0100111010;
#1 $display("%b", po);
# 1  pi=10'b0100111011;
#1 $display("%b", po);
# 1  pi=10'b0100111100;
#1 $display("%b", po);
# 1  pi=10'b0100111101;
#1 $display("%b", po);
# 1  pi=10'b0100111110;
#1 $display("%b", po);
# 1  pi=10'b0100111111;
#1 $display("%b", po);
# 1  pi=10'b0101000000;
#1 $display("%b", po);
# 1  pi=10'b0101000001;
#1 $display("%b", po);
# 1  pi=10'b0101000010;
#1 $display("%b", po);
# 1  pi=10'b0101000011;
#1 $display("%b", po);
# 1  pi=10'b0101000100;
#1 $display("%b", po);
# 1  pi=10'b0101000101;
#1 $display("%b", po);
# 1  pi=10'b0101000110;
#1 $display("%b", po);
# 1  pi=10'b0101000111;
#1 $display("%b", po);
# 1  pi=10'b0101001000;
#1 $display("%b", po);
# 1  pi=10'b0101001001;
#1 $display("%b", po);
# 1  pi=10'b0101001010;
#1 $display("%b", po);
# 1  pi=10'b0101001011;
#1 $display("%b", po);
# 1  pi=10'b0101001100;
#1 $display("%b", po);
# 1  pi=10'b0101001101;
#1 $display("%b", po);
# 1  pi=10'b0101001110;
#1 $display("%b", po);
# 1  pi=10'b0101001111;
#1 $display("%b", po);
# 1  pi=10'b0101010000;
#1 $display("%b", po);
# 1  pi=10'b0101010001;
#1 $display("%b", po);
# 1  pi=10'b0101010010;
#1 $display("%b", po);
# 1  pi=10'b0101010011;
#1 $display("%b", po);
# 1  pi=10'b0101010100;
#1 $display("%b", po);
# 1  pi=10'b0101010101;
#1 $display("%b", po);
# 1  pi=10'b0101010110;
#1 $display("%b", po);
# 1  pi=10'b0101010111;
#1 $display("%b", po);
# 1  pi=10'b0101011000;
#1 $display("%b", po);
# 1  pi=10'b0101011001;
#1 $display("%b", po);
# 1  pi=10'b0101011010;
#1 $display("%b", po);
# 1  pi=10'b0101011011;
#1 $display("%b", po);
# 1  pi=10'b0101011100;
#1 $display("%b", po);
# 1  pi=10'b0101011101;
#1 $display("%b", po);
# 1  pi=10'b0101011110;
#1 $display("%b", po);
# 1  pi=10'b0101011111;
#1 $display("%b", po);
# 1  pi=10'b0101100000;
#1 $display("%b", po);
# 1  pi=10'b0101100001;
#1 $display("%b", po);
# 1  pi=10'b0101100010;
#1 $display("%b", po);
# 1  pi=10'b0101100011;
#1 $display("%b", po);
# 1  pi=10'b0101100100;
#1 $display("%b", po);
# 1  pi=10'b0101100101;
#1 $display("%b", po);
# 1  pi=10'b0101100110;
#1 $display("%b", po);
# 1  pi=10'b0101100111;
#1 $display("%b", po);
# 1  pi=10'b0101101000;
#1 $display("%b", po);
# 1  pi=10'b0101101001;
#1 $display("%b", po);
# 1  pi=10'b0101101010;
#1 $display("%b", po);
# 1  pi=10'b0101101011;
#1 $display("%b", po);
# 1  pi=10'b0101101100;
#1 $display("%b", po);
# 1  pi=10'b0101101101;
#1 $display("%b", po);
# 1  pi=10'b0101101110;
#1 $display("%b", po);
# 1  pi=10'b0101101111;
#1 $display("%b", po);
# 1  pi=10'b0101110000;
#1 $display("%b", po);
# 1  pi=10'b0101110001;
#1 $display("%b", po);
# 1  pi=10'b0101110010;
#1 $display("%b", po);
# 1  pi=10'b0101110011;
#1 $display("%b", po);
# 1  pi=10'b0101110100;
#1 $display("%b", po);
# 1  pi=10'b0101110101;
#1 $display("%b", po);
# 1  pi=10'b0101110110;
#1 $display("%b", po);
# 1  pi=10'b0101110111;
#1 $display("%b", po);
# 1  pi=10'b0101111000;
#1 $display("%b", po);
# 1  pi=10'b0101111001;
#1 $display("%b", po);
# 1  pi=10'b0101111010;
#1 $display("%b", po);
# 1  pi=10'b0101111011;
#1 $display("%b", po);
# 1  pi=10'b0101111100;
#1 $display("%b", po);
# 1  pi=10'b0101111101;
#1 $display("%b", po);
# 1  pi=10'b0101111110;
#1 $display("%b", po);
# 1  pi=10'b0101111111;
#1 $display("%b", po);
# 1  pi=10'b0110000000;
#1 $display("%b", po);
# 1  pi=10'b0110000001;
#1 $display("%b", po);
# 1  pi=10'b0110000010;
#1 $display("%b", po);
# 1  pi=10'b0110000011;
#1 $display("%b", po);
# 1  pi=10'b0110000100;
#1 $display("%b", po);
# 1  pi=10'b0110000101;
#1 $display("%b", po);
# 1  pi=10'b0110000110;
#1 $display("%b", po);
# 1  pi=10'b0110000111;
#1 $display("%b", po);
# 1  pi=10'b0110001000;
#1 $display("%b", po);
# 1  pi=10'b0110001001;
#1 $display("%b", po);
# 1  pi=10'b0110001010;
#1 $display("%b", po);
# 1  pi=10'b0110001011;
#1 $display("%b", po);
# 1  pi=10'b0110001100;
#1 $display("%b", po);
# 1  pi=10'b0110001101;
#1 $display("%b", po);
# 1  pi=10'b0110001110;
#1 $display("%b", po);
# 1  pi=10'b0110001111;
#1 $display("%b", po);
# 1  pi=10'b0110010000;
#1 $display("%b", po);
# 1  pi=10'b0110010001;
#1 $display("%b", po);
# 1  pi=10'b0110010010;
#1 $display("%b", po);
# 1  pi=10'b0110010011;
#1 $display("%b", po);
# 1  pi=10'b0110010100;
#1 $display("%b", po);
# 1  pi=10'b0110010101;
#1 $display("%b", po);
# 1  pi=10'b0110010110;
#1 $display("%b", po);
# 1  pi=10'b0110010111;
#1 $display("%b", po);
# 1  pi=10'b0110011000;
#1 $display("%b", po);
# 1  pi=10'b0110011001;
#1 $display("%b", po);
# 1  pi=10'b0110011010;
#1 $display("%b", po);
# 1  pi=10'b0110011011;
#1 $display("%b", po);
# 1  pi=10'b0110011100;
#1 $display("%b", po);
# 1  pi=10'b0110011101;
#1 $display("%b", po);
# 1  pi=10'b0110011110;
#1 $display("%b", po);
# 1  pi=10'b0110011111;
#1 $display("%b", po);
# 1  pi=10'b0110100000;
#1 $display("%b", po);
# 1  pi=10'b0110100001;
#1 $display("%b", po);
# 1  pi=10'b0110100010;
#1 $display("%b", po);
# 1  pi=10'b0110100011;
#1 $display("%b", po);
# 1  pi=10'b0110100100;
#1 $display("%b", po);
# 1  pi=10'b0110100101;
#1 $display("%b", po);
# 1  pi=10'b0110100110;
#1 $display("%b", po);
# 1  pi=10'b0110100111;
#1 $display("%b", po);
# 1  pi=10'b0110101000;
#1 $display("%b", po);
# 1  pi=10'b0110101001;
#1 $display("%b", po);
# 1  pi=10'b0110101010;
#1 $display("%b", po);
# 1  pi=10'b0110101011;
#1 $display("%b", po);
# 1  pi=10'b0110101100;
#1 $display("%b", po);
# 1  pi=10'b0110101101;
#1 $display("%b", po);
# 1  pi=10'b0110101110;
#1 $display("%b", po);
# 1  pi=10'b0110101111;
#1 $display("%b", po);
# 1  pi=10'b0110110000;
#1 $display("%b", po);
# 1  pi=10'b0110110001;
#1 $display("%b", po);
# 1  pi=10'b0110110010;
#1 $display("%b", po);
# 1  pi=10'b0110110011;
#1 $display("%b", po);
# 1  pi=10'b0110110100;
#1 $display("%b", po);
# 1  pi=10'b0110110101;
#1 $display("%b", po);
# 1  pi=10'b0110110110;
#1 $display("%b", po);
# 1  pi=10'b0110110111;
#1 $display("%b", po);
# 1  pi=10'b0110111000;
#1 $display("%b", po);
# 1  pi=10'b0110111001;
#1 $display("%b", po);
# 1  pi=10'b0110111010;
#1 $display("%b", po);
# 1  pi=10'b0110111011;
#1 $display("%b", po);
# 1  pi=10'b0110111100;
#1 $display("%b", po);
# 1  pi=10'b0110111101;
#1 $display("%b", po);
# 1  pi=10'b0110111110;
#1 $display("%b", po);
# 1  pi=10'b0110111111;
#1 $display("%b", po);
# 1  pi=10'b0111000000;
#1 $display("%b", po);
# 1  pi=10'b0111000001;
#1 $display("%b", po);
# 1  pi=10'b0111000010;
#1 $display("%b", po);
# 1  pi=10'b0111000011;
#1 $display("%b", po);
# 1  pi=10'b0111000100;
#1 $display("%b", po);
# 1  pi=10'b0111000101;
#1 $display("%b", po);
# 1  pi=10'b0111000110;
#1 $display("%b", po);
# 1  pi=10'b0111000111;
#1 $display("%b", po);
# 1  pi=10'b0111001000;
#1 $display("%b", po);
# 1  pi=10'b0111001001;
#1 $display("%b", po);
# 1  pi=10'b0111001010;
#1 $display("%b", po);
# 1  pi=10'b0111001011;
#1 $display("%b", po);
# 1  pi=10'b0111001100;
#1 $display("%b", po);
# 1  pi=10'b0111001101;
#1 $display("%b", po);
# 1  pi=10'b0111001110;
#1 $display("%b", po);
# 1  pi=10'b0111001111;
#1 $display("%b", po);
# 1  pi=10'b0111010000;
#1 $display("%b", po);
# 1  pi=10'b0111010001;
#1 $display("%b", po);
# 1  pi=10'b0111010010;
#1 $display("%b", po);
# 1  pi=10'b0111010011;
#1 $display("%b", po);
# 1  pi=10'b0111010100;
#1 $display("%b", po);
# 1  pi=10'b0111010101;
#1 $display("%b", po);
# 1  pi=10'b0111010110;
#1 $display("%b", po);
# 1  pi=10'b0111010111;
#1 $display("%b", po);
# 1  pi=10'b0111011000;
#1 $display("%b", po);
# 1  pi=10'b0111011001;
#1 $display("%b", po);
# 1  pi=10'b0111011010;
#1 $display("%b", po);
# 1  pi=10'b0111011011;
#1 $display("%b", po);
# 1  pi=10'b0111011100;
#1 $display("%b", po);
# 1  pi=10'b0111011101;
#1 $display("%b", po);
# 1  pi=10'b0111011110;
#1 $display("%b", po);
# 1  pi=10'b0111011111;
#1 $display("%b", po);
# 1  pi=10'b0111100000;
#1 $display("%b", po);
# 1  pi=10'b0111100001;
#1 $display("%b", po);
# 1  pi=10'b0111100010;
#1 $display("%b", po);
# 1  pi=10'b0111100011;
#1 $display("%b", po);
# 1  pi=10'b0111100100;
#1 $display("%b", po);
# 1  pi=10'b0111100101;
#1 $display("%b", po);
# 1  pi=10'b0111100110;
#1 $display("%b", po);
# 1  pi=10'b0111100111;
#1 $display("%b", po);
# 1  pi=10'b0111101000;
#1 $display("%b", po);
# 1  pi=10'b0111101001;
#1 $display("%b", po);
# 1  pi=10'b0111101010;
#1 $display("%b", po);
# 1  pi=10'b0111101011;
#1 $display("%b", po);
# 1  pi=10'b0111101100;
#1 $display("%b", po);
# 1  pi=10'b0111101101;
#1 $display("%b", po);
# 1  pi=10'b0111101110;
#1 $display("%b", po);
# 1  pi=10'b0111101111;
#1 $display("%b", po);
# 1  pi=10'b0111110000;
#1 $display("%b", po);
# 1  pi=10'b0111110001;
#1 $display("%b", po);
# 1  pi=10'b0111110010;
#1 $display("%b", po);
# 1  pi=10'b0111110011;
#1 $display("%b", po);
# 1  pi=10'b0111110100;
#1 $display("%b", po);
# 1  pi=10'b0111110101;
#1 $display("%b", po);
# 1  pi=10'b0111110110;
#1 $display("%b", po);
# 1  pi=10'b0111110111;
#1 $display("%b", po);
# 1  pi=10'b0111111000;
#1 $display("%b", po);
# 1  pi=10'b0111111001;
#1 $display("%b", po);
# 1  pi=10'b0111111010;
#1 $display("%b", po);
# 1  pi=10'b0111111011;
#1 $display("%b", po);
# 1  pi=10'b0111111100;
#1 $display("%b", po);
# 1  pi=10'b0111111101;
#1 $display("%b", po);
# 1  pi=10'b0111111110;
#1 $display("%b", po);
# 1  pi=10'b0111111111;
#1 $display("%b", po);
# 1  pi=10'b1000000000;
#1 $display("%b", po);
# 1  pi=10'b1000000001;
#1 $display("%b", po);
# 1  pi=10'b1000000010;
#1 $display("%b", po);
# 1  pi=10'b1000000011;
#1 $display("%b", po);
# 1  pi=10'b1000000100;
#1 $display("%b", po);
# 1  pi=10'b1000000101;
#1 $display("%b", po);
# 1  pi=10'b1000000110;
#1 $display("%b", po);
# 1  pi=10'b1000000111;
#1 $display("%b", po);
# 1  pi=10'b1000001000;
#1 $display("%b", po);
# 1  pi=10'b1000001001;
#1 $display("%b", po);
# 1  pi=10'b1000001010;
#1 $display("%b", po);
# 1  pi=10'b1000001011;
#1 $display("%b", po);
# 1  pi=10'b1000001100;
#1 $display("%b", po);
# 1  pi=10'b1000001101;
#1 $display("%b", po);
# 1  pi=10'b1000001110;
#1 $display("%b", po);
# 1  pi=10'b1000001111;
#1 $display("%b", po);
# 1  pi=10'b1000010000;
#1 $display("%b", po);
# 1  pi=10'b1000010001;
#1 $display("%b", po);
# 1  pi=10'b1000010010;
#1 $display("%b", po);
# 1  pi=10'b1000010011;
#1 $display("%b", po);
# 1  pi=10'b1000010100;
#1 $display("%b", po);
# 1  pi=10'b1000010101;
#1 $display("%b", po);
# 1  pi=10'b1000010110;
#1 $display("%b", po);
# 1  pi=10'b1000010111;
#1 $display("%b", po);
# 1  pi=10'b1000011000;
#1 $display("%b", po);
# 1  pi=10'b1000011001;
#1 $display("%b", po);
# 1  pi=10'b1000011010;
#1 $display("%b", po);
# 1  pi=10'b1000011011;
#1 $display("%b", po);
# 1  pi=10'b1000011100;
#1 $display("%b", po);
# 1  pi=10'b1000011101;
#1 $display("%b", po);
# 1  pi=10'b1000011110;
#1 $display("%b", po);
# 1  pi=10'b1000011111;
#1 $display("%b", po);
# 1  pi=10'b1000100000;
#1 $display("%b", po);
# 1  pi=10'b1000100001;
#1 $display("%b", po);
# 1  pi=10'b1000100010;
#1 $display("%b", po);
# 1  pi=10'b1000100011;
#1 $display("%b", po);
# 1  pi=10'b1000100100;
#1 $display("%b", po);
# 1  pi=10'b1000100101;
#1 $display("%b", po);
# 1  pi=10'b1000100110;
#1 $display("%b", po);
# 1  pi=10'b1000100111;
#1 $display("%b", po);
# 1  pi=10'b1000101000;
#1 $display("%b", po);
# 1  pi=10'b1000101001;
#1 $display("%b", po);
# 1  pi=10'b1000101010;
#1 $display("%b", po);
# 1  pi=10'b1000101011;
#1 $display("%b", po);
# 1  pi=10'b1000101100;
#1 $display("%b", po);
# 1  pi=10'b1000101101;
#1 $display("%b", po);
# 1  pi=10'b1000101110;
#1 $display("%b", po);
# 1  pi=10'b1000101111;
#1 $display("%b", po);
# 1  pi=10'b1000110000;
#1 $display("%b", po);
# 1  pi=10'b1000110001;
#1 $display("%b", po);
# 1  pi=10'b1000110010;
#1 $display("%b", po);
# 1  pi=10'b1000110011;
#1 $display("%b", po);
# 1  pi=10'b1000110100;
#1 $display("%b", po);
# 1  pi=10'b1000110101;
#1 $display("%b", po);
# 1  pi=10'b1000110110;
#1 $display("%b", po);
# 1  pi=10'b1000110111;
#1 $display("%b", po);
# 1  pi=10'b1000111000;
#1 $display("%b", po);
# 1  pi=10'b1000111001;
#1 $display("%b", po);
# 1  pi=10'b1000111010;
#1 $display("%b", po);
# 1  pi=10'b1000111011;
#1 $display("%b", po);
# 1  pi=10'b1000111100;
#1 $display("%b", po);
# 1  pi=10'b1000111101;
#1 $display("%b", po);
# 1  pi=10'b1000111110;
#1 $display("%b", po);
# 1  pi=10'b1000111111;
#1 $display("%b", po);
# 1  pi=10'b1001000000;
#1 $display("%b", po);
# 1  pi=10'b1001000001;
#1 $display("%b", po);
# 1  pi=10'b1001000010;
#1 $display("%b", po);
# 1  pi=10'b1001000011;
#1 $display("%b", po);
# 1  pi=10'b1001000100;
#1 $display("%b", po);
# 1  pi=10'b1001000101;
#1 $display("%b", po);
# 1  pi=10'b1001000110;
#1 $display("%b", po);
# 1  pi=10'b1001000111;
#1 $display("%b", po);
# 1  pi=10'b1001001000;
#1 $display("%b", po);
# 1  pi=10'b1001001001;
#1 $display("%b", po);
# 1  pi=10'b1001001010;
#1 $display("%b", po);
# 1  pi=10'b1001001011;
#1 $display("%b", po);
# 1  pi=10'b1001001100;
#1 $display("%b", po);
# 1  pi=10'b1001001101;
#1 $display("%b", po);
# 1  pi=10'b1001001110;
#1 $display("%b", po);
# 1  pi=10'b1001001111;
#1 $display("%b", po);
# 1  pi=10'b1001010000;
#1 $display("%b", po);
# 1  pi=10'b1001010001;
#1 $display("%b", po);
# 1  pi=10'b1001010010;
#1 $display("%b", po);
# 1  pi=10'b1001010011;
#1 $display("%b", po);
# 1  pi=10'b1001010100;
#1 $display("%b", po);
# 1  pi=10'b1001010101;
#1 $display("%b", po);
# 1  pi=10'b1001010110;
#1 $display("%b", po);
# 1  pi=10'b1001010111;
#1 $display("%b", po);
# 1  pi=10'b1001011000;
#1 $display("%b", po);
# 1  pi=10'b1001011001;
#1 $display("%b", po);
# 1  pi=10'b1001011010;
#1 $display("%b", po);
# 1  pi=10'b1001011011;
#1 $display("%b", po);
# 1  pi=10'b1001011100;
#1 $display("%b", po);
# 1  pi=10'b1001011101;
#1 $display("%b", po);
# 1  pi=10'b1001011110;
#1 $display("%b", po);
# 1  pi=10'b1001011111;
#1 $display("%b", po);
# 1  pi=10'b1001100000;
#1 $display("%b", po);
# 1  pi=10'b1001100001;
#1 $display("%b", po);
# 1  pi=10'b1001100010;
#1 $display("%b", po);
# 1  pi=10'b1001100011;
#1 $display("%b", po);
# 1  pi=10'b1001100100;
#1 $display("%b", po);
# 1  pi=10'b1001100101;
#1 $display("%b", po);
# 1  pi=10'b1001100110;
#1 $display("%b", po);
# 1  pi=10'b1001100111;
#1 $display("%b", po);
# 1  pi=10'b1001101000;
#1 $display("%b", po);
# 1  pi=10'b1001101001;
#1 $display("%b", po);
# 1  pi=10'b1001101010;
#1 $display("%b", po);
# 1  pi=10'b1001101011;
#1 $display("%b", po);
# 1  pi=10'b1001101100;
#1 $display("%b", po);
# 1  pi=10'b1001101101;
#1 $display("%b", po);
# 1  pi=10'b1001101110;
#1 $display("%b", po);
# 1  pi=10'b1001101111;
#1 $display("%b", po);
# 1  pi=10'b1001110000;
#1 $display("%b", po);
# 1  pi=10'b1001110001;
#1 $display("%b", po);
# 1  pi=10'b1001110010;
#1 $display("%b", po);
# 1  pi=10'b1001110011;
#1 $display("%b", po);
# 1  pi=10'b1001110100;
#1 $display("%b", po);
# 1  pi=10'b1001110101;
#1 $display("%b", po);
# 1  pi=10'b1001110110;
#1 $display("%b", po);
# 1  pi=10'b1001110111;
#1 $display("%b", po);
# 1  pi=10'b1001111000;
#1 $display("%b", po);
# 1  pi=10'b1001111001;
#1 $display("%b", po);
# 1  pi=10'b1001111010;
#1 $display("%b", po);
# 1  pi=10'b1001111011;
#1 $display("%b", po);
# 1  pi=10'b1001111100;
#1 $display("%b", po);
# 1  pi=10'b1001111101;
#1 $display("%b", po);
# 1  pi=10'b1001111110;
#1 $display("%b", po);
# 1  pi=10'b1001111111;
#1 $display("%b", po);
# 1  pi=10'b1010000000;
#1 $display("%b", po);
# 1  pi=10'b1010000001;
#1 $display("%b", po);
# 1  pi=10'b1010000010;
#1 $display("%b", po);
# 1  pi=10'b1010000011;
#1 $display("%b", po);
# 1  pi=10'b1010000100;
#1 $display("%b", po);
# 1  pi=10'b1010000101;
#1 $display("%b", po);
# 1  pi=10'b1010000110;
#1 $display("%b", po);
# 1  pi=10'b1010000111;
#1 $display("%b", po);
# 1  pi=10'b1010001000;
#1 $display("%b", po);
# 1  pi=10'b1010001001;
#1 $display("%b", po);
# 1  pi=10'b1010001010;
#1 $display("%b", po);
# 1  pi=10'b1010001011;
#1 $display("%b", po);
# 1  pi=10'b1010001100;
#1 $display("%b", po);
# 1  pi=10'b1010001101;
#1 $display("%b", po);
# 1  pi=10'b1010001110;
#1 $display("%b", po);
# 1  pi=10'b1010001111;
#1 $display("%b", po);
# 1  pi=10'b1010010000;
#1 $display("%b", po);
# 1  pi=10'b1010010001;
#1 $display("%b", po);
# 1  pi=10'b1010010010;
#1 $display("%b", po);
# 1  pi=10'b1010010011;
#1 $display("%b", po);
# 1  pi=10'b1010010100;
#1 $display("%b", po);
# 1  pi=10'b1010010101;
#1 $display("%b", po);
# 1  pi=10'b1010010110;
#1 $display("%b", po);
# 1  pi=10'b1010010111;
#1 $display("%b", po);
# 1  pi=10'b1010011000;
#1 $display("%b", po);
# 1  pi=10'b1010011001;
#1 $display("%b", po);
# 1  pi=10'b1010011010;
#1 $display("%b", po);
# 1  pi=10'b1010011011;
#1 $display("%b", po);
# 1  pi=10'b1010011100;
#1 $display("%b", po);
# 1  pi=10'b1010011101;
#1 $display("%b", po);
# 1  pi=10'b1010011110;
#1 $display("%b", po);
# 1  pi=10'b1010011111;
#1 $display("%b", po);
# 1  pi=10'b1010100000;
#1 $display("%b", po);
# 1  pi=10'b1010100001;
#1 $display("%b", po);
# 1  pi=10'b1010100010;
#1 $display("%b", po);
# 1  pi=10'b1010100011;
#1 $display("%b", po);
# 1  pi=10'b1010100100;
#1 $display("%b", po);
# 1  pi=10'b1010100101;
#1 $display("%b", po);
# 1  pi=10'b1010100110;
#1 $display("%b", po);
# 1  pi=10'b1010100111;
#1 $display("%b", po);
# 1  pi=10'b1010101000;
#1 $display("%b", po);
# 1  pi=10'b1010101001;
#1 $display("%b", po);
# 1  pi=10'b1010101010;
#1 $display("%b", po);
# 1  pi=10'b1010101011;
#1 $display("%b", po);
# 1  pi=10'b1010101100;
#1 $display("%b", po);
# 1  pi=10'b1010101101;
#1 $display("%b", po);
# 1  pi=10'b1010101110;
#1 $display("%b", po);
# 1  pi=10'b1010101111;
#1 $display("%b", po);
# 1  pi=10'b1010110000;
#1 $display("%b", po);
# 1  pi=10'b1010110001;
#1 $display("%b", po);
# 1  pi=10'b1010110010;
#1 $display("%b", po);
# 1  pi=10'b1010110011;
#1 $display("%b", po);
# 1  pi=10'b1010110100;
#1 $display("%b", po);
# 1  pi=10'b1010110101;
#1 $display("%b", po);
# 1  pi=10'b1010110110;
#1 $display("%b", po);
# 1  pi=10'b1010110111;
#1 $display("%b", po);
# 1  pi=10'b1010111000;
#1 $display("%b", po);
# 1  pi=10'b1010111001;
#1 $display("%b", po);
# 1  pi=10'b1010111010;
#1 $display("%b", po);
# 1  pi=10'b1010111011;
#1 $display("%b", po);
# 1  pi=10'b1010111100;
#1 $display("%b", po);
# 1  pi=10'b1010111101;
#1 $display("%b", po);
# 1  pi=10'b1010111110;
#1 $display("%b", po);
# 1  pi=10'b1010111111;
#1 $display("%b", po);
# 1  pi=10'b1011000000;
#1 $display("%b", po);
# 1  pi=10'b1011000001;
#1 $display("%b", po);
# 1  pi=10'b1011000010;
#1 $display("%b", po);
# 1  pi=10'b1011000011;
#1 $display("%b", po);
# 1  pi=10'b1011000100;
#1 $display("%b", po);
# 1  pi=10'b1011000101;
#1 $display("%b", po);
# 1  pi=10'b1011000110;
#1 $display("%b", po);
# 1  pi=10'b1011000111;
#1 $display("%b", po);
# 1  pi=10'b1011001000;
#1 $display("%b", po);
# 1  pi=10'b1011001001;
#1 $display("%b", po);
# 1  pi=10'b1011001010;
#1 $display("%b", po);
# 1  pi=10'b1011001011;
#1 $display("%b", po);
# 1  pi=10'b1011001100;
#1 $display("%b", po);
# 1  pi=10'b1011001101;
#1 $display("%b", po);
# 1  pi=10'b1011001110;
#1 $display("%b", po);
# 1  pi=10'b1011001111;
#1 $display("%b", po);
# 1  pi=10'b1011010000;
#1 $display("%b", po);
# 1  pi=10'b1011010001;
#1 $display("%b", po);
# 1  pi=10'b1011010010;
#1 $display("%b", po);
# 1  pi=10'b1011010011;
#1 $display("%b", po);
# 1  pi=10'b1011010100;
#1 $display("%b", po);
# 1  pi=10'b1011010101;
#1 $display("%b", po);
# 1  pi=10'b1011010110;
#1 $display("%b", po);
# 1  pi=10'b1011010111;
#1 $display("%b", po);
# 1  pi=10'b1011011000;
#1 $display("%b", po);
# 1  pi=10'b1011011001;
#1 $display("%b", po);
# 1  pi=10'b1011011010;
#1 $display("%b", po);
# 1  pi=10'b1011011011;
#1 $display("%b", po);
# 1  pi=10'b1011011100;
#1 $display("%b", po);
# 1  pi=10'b1011011101;
#1 $display("%b", po);
# 1  pi=10'b1011011110;
#1 $display("%b", po);
# 1  pi=10'b1011011111;
#1 $display("%b", po);
# 1  pi=10'b1011100000;
#1 $display("%b", po);
# 1  pi=10'b1011100001;
#1 $display("%b", po);
# 1  pi=10'b1011100010;
#1 $display("%b", po);
# 1  pi=10'b1011100011;
#1 $display("%b", po);
# 1  pi=10'b1011100100;
#1 $display("%b", po);
# 1  pi=10'b1011100101;
#1 $display("%b", po);
# 1  pi=10'b1011100110;
#1 $display("%b", po);
# 1  pi=10'b1011100111;
#1 $display("%b", po);
# 1  pi=10'b1011101000;
#1 $display("%b", po);
# 1  pi=10'b1011101001;
#1 $display("%b", po);
# 1  pi=10'b1011101010;
#1 $display("%b", po);
# 1  pi=10'b1011101011;
#1 $display("%b", po);
# 1  pi=10'b1011101100;
#1 $display("%b", po);
# 1  pi=10'b1011101101;
#1 $display("%b", po);
# 1  pi=10'b1011101110;
#1 $display("%b", po);
# 1  pi=10'b1011101111;
#1 $display("%b", po);
# 1  pi=10'b1011110000;
#1 $display("%b", po);
# 1  pi=10'b1011110001;
#1 $display("%b", po);
# 1  pi=10'b1011110010;
#1 $display("%b", po);
# 1  pi=10'b1011110011;
#1 $display("%b", po);
# 1  pi=10'b1011110100;
#1 $display("%b", po);
# 1  pi=10'b1011110101;
#1 $display("%b", po);
# 1  pi=10'b1011110110;
#1 $display("%b", po);
# 1  pi=10'b1011110111;
#1 $display("%b", po);
# 1  pi=10'b1011111000;
#1 $display("%b", po);
# 1  pi=10'b1011111001;
#1 $display("%b", po);
# 1  pi=10'b1011111010;
#1 $display("%b", po);
# 1  pi=10'b1011111011;
#1 $display("%b", po);
# 1  pi=10'b1011111100;
#1 $display("%b", po);
# 1  pi=10'b1011111101;
#1 $display("%b", po);
# 1  pi=10'b1011111110;
#1 $display("%b", po);
# 1  pi=10'b1011111111;
#1 $display("%b", po);
# 1  pi=10'b1100000000;
#1 $display("%b", po);
# 1  pi=10'b1100000001;
#1 $display("%b", po);
# 1  pi=10'b1100000010;
#1 $display("%b", po);
# 1  pi=10'b1100000011;
#1 $display("%b", po);
# 1  pi=10'b1100000100;
#1 $display("%b", po);
# 1  pi=10'b1100000101;
#1 $display("%b", po);
# 1  pi=10'b1100000110;
#1 $display("%b", po);
# 1  pi=10'b1100000111;
#1 $display("%b", po);
# 1  pi=10'b1100001000;
#1 $display("%b", po);
# 1  pi=10'b1100001001;
#1 $display("%b", po);
# 1  pi=10'b1100001010;
#1 $display("%b", po);
# 1  pi=10'b1100001011;
#1 $display("%b", po);
# 1  pi=10'b1100001100;
#1 $display("%b", po);
# 1  pi=10'b1100001101;
#1 $display("%b", po);
# 1  pi=10'b1100001110;
#1 $display("%b", po);
# 1  pi=10'b1100001111;
#1 $display("%b", po);
# 1  pi=10'b1100010000;
#1 $display("%b", po);
# 1  pi=10'b1100010001;
#1 $display("%b", po);
# 1  pi=10'b1100010010;
#1 $display("%b", po);
# 1  pi=10'b1100010011;
#1 $display("%b", po);
# 1  pi=10'b1100010100;
#1 $display("%b", po);
# 1  pi=10'b1100010101;
#1 $display("%b", po);
# 1  pi=10'b1100010110;
#1 $display("%b", po);
# 1  pi=10'b1100010111;
#1 $display("%b", po);
# 1  pi=10'b1100011000;
#1 $display("%b", po);
# 1  pi=10'b1100011001;
#1 $display("%b", po);
# 1  pi=10'b1100011010;
#1 $display("%b", po);
# 1  pi=10'b1100011011;
#1 $display("%b", po);
# 1  pi=10'b1100011100;
#1 $display("%b", po);
# 1  pi=10'b1100011101;
#1 $display("%b", po);
# 1  pi=10'b1100011110;
#1 $display("%b", po);
# 1  pi=10'b1100011111;
#1 $display("%b", po);
# 1  pi=10'b1100100000;
#1 $display("%b", po);
# 1  pi=10'b1100100001;
#1 $display("%b", po);
# 1  pi=10'b1100100010;
#1 $display("%b", po);
# 1  pi=10'b1100100011;
#1 $display("%b", po);
# 1  pi=10'b1100100100;
#1 $display("%b", po);
# 1  pi=10'b1100100101;
#1 $display("%b", po);
# 1  pi=10'b1100100110;
#1 $display("%b", po);
# 1  pi=10'b1100100111;
#1 $display("%b", po);
# 1  pi=10'b1100101000;
#1 $display("%b", po);
# 1  pi=10'b1100101001;
#1 $display("%b", po);
# 1  pi=10'b1100101010;
#1 $display("%b", po);
# 1  pi=10'b1100101011;
#1 $display("%b", po);
# 1  pi=10'b1100101100;
#1 $display("%b", po);
# 1  pi=10'b1100101101;
#1 $display("%b", po);
# 1  pi=10'b1100101110;
#1 $display("%b", po);
# 1  pi=10'b1100101111;
#1 $display("%b", po);
# 1  pi=10'b1100110000;
#1 $display("%b", po);
# 1  pi=10'b1100110001;
#1 $display("%b", po);
# 1  pi=10'b1100110010;
#1 $display("%b", po);
# 1  pi=10'b1100110011;
#1 $display("%b", po);
# 1  pi=10'b1100110100;
#1 $display("%b", po);
# 1  pi=10'b1100110101;
#1 $display("%b", po);
# 1  pi=10'b1100110110;
#1 $display("%b", po);
# 1  pi=10'b1100110111;
#1 $display("%b", po);
# 1  pi=10'b1100111000;
#1 $display("%b", po);
# 1  pi=10'b1100111001;
#1 $display("%b", po);
# 1  pi=10'b1100111010;
#1 $display("%b", po);
# 1  pi=10'b1100111011;
#1 $display("%b", po);
# 1  pi=10'b1100111100;
#1 $display("%b", po);
# 1  pi=10'b1100111101;
#1 $display("%b", po);
# 1  pi=10'b1100111110;
#1 $display("%b", po);
# 1  pi=10'b1100111111;
#1 $display("%b", po);
# 1  pi=10'b1101000000;
#1 $display("%b", po);
# 1  pi=10'b1101000001;
#1 $display("%b", po);
# 1  pi=10'b1101000010;
#1 $display("%b", po);
# 1  pi=10'b1101000011;
#1 $display("%b", po);
# 1  pi=10'b1101000100;
#1 $display("%b", po);
# 1  pi=10'b1101000101;
#1 $display("%b", po);
# 1  pi=10'b1101000110;
#1 $display("%b", po);
# 1  pi=10'b1101000111;
#1 $display("%b", po);
# 1  pi=10'b1101001000;
#1 $display("%b", po);
# 1  pi=10'b1101001001;
#1 $display("%b", po);
# 1  pi=10'b1101001010;
#1 $display("%b", po);
# 1  pi=10'b1101001011;
#1 $display("%b", po);
# 1  pi=10'b1101001100;
#1 $display("%b", po);
# 1  pi=10'b1101001101;
#1 $display("%b", po);
# 1  pi=10'b1101001110;
#1 $display("%b", po);
# 1  pi=10'b1101001111;
#1 $display("%b", po);
# 1  pi=10'b1101010000;
#1 $display("%b", po);
# 1  pi=10'b1101010001;
#1 $display("%b", po);
# 1  pi=10'b1101010010;
#1 $display("%b", po);
# 1  pi=10'b1101010011;
#1 $display("%b", po);
# 1  pi=10'b1101010100;
#1 $display("%b", po);
# 1  pi=10'b1101010101;
#1 $display("%b", po);
# 1  pi=10'b1101010110;
#1 $display("%b", po);
# 1  pi=10'b1101010111;
#1 $display("%b", po);
# 1  pi=10'b1101011000;
#1 $display("%b", po);
# 1  pi=10'b1101011001;
#1 $display("%b", po);
# 1  pi=10'b1101011010;
#1 $display("%b", po);
# 1  pi=10'b1101011011;
#1 $display("%b", po);
# 1  pi=10'b1101011100;
#1 $display("%b", po);
# 1  pi=10'b1101011101;
#1 $display("%b", po);
# 1  pi=10'b1101011110;
#1 $display("%b", po);
# 1  pi=10'b1101011111;
#1 $display("%b", po);
# 1  pi=10'b1101100000;
#1 $display("%b", po);
# 1  pi=10'b1101100001;
#1 $display("%b", po);
# 1  pi=10'b1101100010;
#1 $display("%b", po);
# 1  pi=10'b1101100011;
#1 $display("%b", po);
# 1  pi=10'b1101100100;
#1 $display("%b", po);
# 1  pi=10'b1101100101;
#1 $display("%b", po);
# 1  pi=10'b1101100110;
#1 $display("%b", po);
# 1  pi=10'b1101100111;
#1 $display("%b", po);
# 1  pi=10'b1101101000;
#1 $display("%b", po);
# 1  pi=10'b1101101001;
#1 $display("%b", po);
# 1  pi=10'b1101101010;
#1 $display("%b", po);
# 1  pi=10'b1101101011;
#1 $display("%b", po);
# 1  pi=10'b1101101100;
#1 $display("%b", po);
# 1  pi=10'b1101101101;
#1 $display("%b", po);
# 1  pi=10'b1101101110;
#1 $display("%b", po);
# 1  pi=10'b1101101111;
#1 $display("%b", po);
# 1  pi=10'b1101110000;
#1 $display("%b", po);
# 1  pi=10'b1101110001;
#1 $display("%b", po);
# 1  pi=10'b1101110010;
#1 $display("%b", po);
# 1  pi=10'b1101110011;
#1 $display("%b", po);
# 1  pi=10'b1101110100;
#1 $display("%b", po);
# 1  pi=10'b1101110101;
#1 $display("%b", po);
# 1  pi=10'b1101110110;
#1 $display("%b", po);
# 1  pi=10'b1101110111;
#1 $display("%b", po);
# 1  pi=10'b1101111000;
#1 $display("%b", po);
# 1  pi=10'b1101111001;
#1 $display("%b", po);
# 1  pi=10'b1101111010;
#1 $display("%b", po);
# 1  pi=10'b1101111011;
#1 $display("%b", po);
# 1  pi=10'b1101111100;
#1 $display("%b", po);
# 1  pi=10'b1101111101;
#1 $display("%b", po);
# 1  pi=10'b1101111110;
#1 $display("%b", po);
# 1  pi=10'b1101111111;
#1 $display("%b", po);
# 1  pi=10'b1110000000;
#1 $display("%b", po);
# 1  pi=10'b1110000001;
#1 $display("%b", po);
# 1  pi=10'b1110000010;
#1 $display("%b", po);
# 1  pi=10'b1110000011;
#1 $display("%b", po);
# 1  pi=10'b1110000100;
#1 $display("%b", po);
# 1  pi=10'b1110000101;
#1 $display("%b", po);
# 1  pi=10'b1110000110;
#1 $display("%b", po);
# 1  pi=10'b1110000111;
#1 $display("%b", po);
# 1  pi=10'b1110001000;
#1 $display("%b", po);
# 1  pi=10'b1110001001;
#1 $display("%b", po);
# 1  pi=10'b1110001010;
#1 $display("%b", po);
# 1  pi=10'b1110001011;
#1 $display("%b", po);
# 1  pi=10'b1110001100;
#1 $display("%b", po);
# 1  pi=10'b1110001101;
#1 $display("%b", po);
# 1  pi=10'b1110001110;
#1 $display("%b", po);
# 1  pi=10'b1110001111;
#1 $display("%b", po);
# 1  pi=10'b1110010000;
#1 $display("%b", po);
# 1  pi=10'b1110010001;
#1 $display("%b", po);
# 1  pi=10'b1110010010;
#1 $display("%b", po);
# 1  pi=10'b1110010011;
#1 $display("%b", po);
# 1  pi=10'b1110010100;
#1 $display("%b", po);
# 1  pi=10'b1110010101;
#1 $display("%b", po);
# 1  pi=10'b1110010110;
#1 $display("%b", po);
# 1  pi=10'b1110010111;
#1 $display("%b", po);
# 1  pi=10'b1110011000;
#1 $display("%b", po);
# 1  pi=10'b1110011001;
#1 $display("%b", po);
# 1  pi=10'b1110011010;
#1 $display("%b", po);
# 1  pi=10'b1110011011;
#1 $display("%b", po);
# 1  pi=10'b1110011100;
#1 $display("%b", po);
# 1  pi=10'b1110011101;
#1 $display("%b", po);
# 1  pi=10'b1110011110;
#1 $display("%b", po);
# 1  pi=10'b1110011111;
#1 $display("%b", po);
# 1  pi=10'b1110100000;
#1 $display("%b", po);
# 1  pi=10'b1110100001;
#1 $display("%b", po);
# 1  pi=10'b1110100010;
#1 $display("%b", po);
# 1  pi=10'b1110100011;
#1 $display("%b", po);
# 1  pi=10'b1110100100;
#1 $display("%b", po);
# 1  pi=10'b1110100101;
#1 $display("%b", po);
# 1  pi=10'b1110100110;
#1 $display("%b", po);
# 1  pi=10'b1110100111;
#1 $display("%b", po);
# 1  pi=10'b1110101000;
#1 $display("%b", po);
# 1  pi=10'b1110101001;
#1 $display("%b", po);
# 1  pi=10'b1110101010;
#1 $display("%b", po);
# 1  pi=10'b1110101011;
#1 $display("%b", po);
# 1  pi=10'b1110101100;
#1 $display("%b", po);
# 1  pi=10'b1110101101;
#1 $display("%b", po);
# 1  pi=10'b1110101110;
#1 $display("%b", po);
# 1  pi=10'b1110101111;
#1 $display("%b", po);
# 1  pi=10'b1110110000;
#1 $display("%b", po);
# 1  pi=10'b1110110001;
#1 $display("%b", po);
# 1  pi=10'b1110110010;
#1 $display("%b", po);
# 1  pi=10'b1110110011;
#1 $display("%b", po);
# 1  pi=10'b1110110100;
#1 $display("%b", po);
# 1  pi=10'b1110110101;
#1 $display("%b", po);
# 1  pi=10'b1110110110;
#1 $display("%b", po);
# 1  pi=10'b1110110111;
#1 $display("%b", po);
# 1  pi=10'b1110111000;
#1 $display("%b", po);
# 1  pi=10'b1110111001;
#1 $display("%b", po);
# 1  pi=10'b1110111010;
#1 $display("%b", po);
# 1  pi=10'b1110111011;
#1 $display("%b", po);
# 1  pi=10'b1110111100;
#1 $display("%b", po);
# 1  pi=10'b1110111101;
#1 $display("%b", po);
# 1  pi=10'b1110111110;
#1 $display("%b", po);
# 1  pi=10'b1110111111;
#1 $display("%b", po);
# 1  pi=10'b1111000000;
#1 $display("%b", po);
# 1  pi=10'b1111000001;
#1 $display("%b", po);
# 1  pi=10'b1111000010;
#1 $display("%b", po);
# 1  pi=10'b1111000011;
#1 $display("%b", po);
# 1  pi=10'b1111000100;
#1 $display("%b", po);
# 1  pi=10'b1111000101;
#1 $display("%b", po);
# 1  pi=10'b1111000110;
#1 $display("%b", po);
# 1  pi=10'b1111000111;
#1 $display("%b", po);
# 1  pi=10'b1111001000;
#1 $display("%b", po);
# 1  pi=10'b1111001001;
#1 $display("%b", po);
# 1  pi=10'b1111001010;
#1 $display("%b", po);
# 1  pi=10'b1111001011;
#1 $display("%b", po);
# 1  pi=10'b1111001100;
#1 $display("%b", po);
# 1  pi=10'b1111001101;
#1 $display("%b", po);
# 1  pi=10'b1111001110;
#1 $display("%b", po);
# 1  pi=10'b1111001111;
#1 $display("%b", po);
# 1  pi=10'b1111010000;
#1 $display("%b", po);
# 1  pi=10'b1111010001;
#1 $display("%b", po);
# 1  pi=10'b1111010010;
#1 $display("%b", po);
# 1  pi=10'b1111010011;
#1 $display("%b", po);
# 1  pi=10'b1111010100;
#1 $display("%b", po);
# 1  pi=10'b1111010101;
#1 $display("%b", po);
# 1  pi=10'b1111010110;
#1 $display("%b", po);
# 1  pi=10'b1111010111;
#1 $display("%b", po);
# 1  pi=10'b1111011000;
#1 $display("%b", po);
# 1  pi=10'b1111011001;
#1 $display("%b", po);
# 1  pi=10'b1111011010;
#1 $display("%b", po);
# 1  pi=10'b1111011011;
#1 $display("%b", po);
# 1  pi=10'b1111011100;
#1 $display("%b", po);
# 1  pi=10'b1111011101;
#1 $display("%b", po);
# 1  pi=10'b1111011110;
#1 $display("%b", po);
# 1  pi=10'b1111011111;
#1 $display("%b", po);
# 1  pi=10'b1111100000;
#1 $display("%b", po);
# 1  pi=10'b1111100001;
#1 $display("%b", po);
# 1  pi=10'b1111100010;
#1 $display("%b", po);
# 1  pi=10'b1111100011;
#1 $display("%b", po);
# 1  pi=10'b1111100100;
#1 $display("%b", po);
# 1  pi=10'b1111100101;
#1 $display("%b", po);
# 1  pi=10'b1111100110;
#1 $display("%b", po);
# 1  pi=10'b1111100111;
#1 $display("%b", po);
# 1  pi=10'b1111101000;
#1 $display("%b", po);
# 1  pi=10'b1111101001;
#1 $display("%b", po);
# 1  pi=10'b1111101010;
#1 $display("%b", po);
# 1  pi=10'b1111101011;
#1 $display("%b", po);
# 1  pi=10'b1111101100;
#1 $display("%b", po);
# 1  pi=10'b1111101101;
#1 $display("%b", po);
# 1  pi=10'b1111101110;
#1 $display("%b", po);
# 1  pi=10'b1111101111;
#1 $display("%b", po);
# 1  pi=10'b1111110000;
#1 $display("%b", po);
# 1  pi=10'b1111110001;
#1 $display("%b", po);
# 1  pi=10'b1111110010;
#1 $display("%b", po);
# 1  pi=10'b1111110011;
#1 $display("%b", po);
# 1  pi=10'b1111110100;
#1 $display("%b", po);
# 1  pi=10'b1111110101;
#1 $display("%b", po);
# 1  pi=10'b1111110110;
#1 $display("%b", po);
# 1  pi=10'b1111110111;
#1 $display("%b", po);
# 1  pi=10'b1111111000;
#1 $display("%b", po);
# 1  pi=10'b1111111001;
#1 $display("%b", po);
# 1  pi=10'b1111111010;
#1 $display("%b", po);
# 1  pi=10'b1111111011;
#1 $display("%b", po);
# 1  pi=10'b1111111100;
#1 $display("%b", po);
# 1  pi=10'b1111111101;
#1 $display("%b", po);
# 1  pi=10'b1111111110;
#1 $display("%b", po);
# 1  pi=10'b1111111111;
#1 $display("%b", po);
end
endmodule
