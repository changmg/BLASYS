// Benchmark "ex" written by ABC on Thu Jul 14 00:21:31 2022

module ex ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m,
    F  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m;
  output F;
  assign F = ~f & a;
endmodule


