module mult16(\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] 
, \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \r[0] , \r[1] , \r[2] , \r[3] , \r[4] , \r[5] , \r[6] , \r[7] , \r[8] , \r[9] 
, \r[10] , \r[11] , \r[12] , \r[13] , \r[14] , \r[15] , \r[16] , \r[17] , \r[18] , \r[19] , \r[20] , \r[21] , \r[22] , \r[23] , \r[24] , \r[25] , \r[26] , \r[27] , \r[28] , \r[29] , \r[30] 
, \r[31] );
  input \a[0] ;
  input \a[10] ;
  input \a[11] ;
  input \a[12] ;
  input \a[13] ;
  input \a[14] ;
  input \a[15] ;
  input \a[1] ;
  input \a[2] ;
  input \a[3] ;
  input \a[4] ;
  input \a[5] ;
  input \a[6] ;
  input \a[7] ;
  input \a[8] ;
  input \a[9] ;
  input \b[0] ;
  input \b[10] ;
  input \b[11] ;
  input \b[12] ;
  input \b[13] ;
  input \b[14] ;
  input \b[15] ;
  input \b[1] ;
  input \b[2] ;
  input \b[3] ;
  input \b[4] ;
  input \b[5] ;
  input \b[6] ;
  input \b[7] ;
  input \b[8] ;
  input \b[9] ;
  output \r[0] ;
  output \r[10] ;
  output \r[11] ;
  output \r[12] ;
  output \r[13] ;
  output \r[14] ;
  output \r[15] ;
  output \r[16] ;
  output \r[17] ;
  output \r[18] ;
  output \r[19] ;
  output \r[1] ;
  output \r[20] ;
  output \r[21] ;
  output \r[22] ;
  output \r[23] ;
  output \r[24] ;
  output \r[25] ;
  output \r[26] ;
  output \r[27] ;
  output \r[28] ;
  output \r[29] ;
  output \r[2] ;
  output \r[30] ;
  output \r[31] ;
  output \r[3] ;
  output \r[4] ;
  output \r[5] ;
  output \r[6] ;
  output \r[7] ;
  output \r[8] ;
  output \r[9] ;
  top U0 ( .pi00( \a[0] ) , .pi01( \a[1] ) , .pi02( \a[2] ) , .pi03( \a[3] ) , .pi04( \a[4] ) , .pi05( \a[5] ) , .pi06( \a[6] ) , .pi07( \a[7] ) , .pi08( \a[8] ) , .pi09( \a[9] ) , .pi10( \a[10] ) , .pi11( \a[11] ) , .pi12( \a[12] ) , .pi13( \a[13] ) , .pi14( \a[14] ) , .pi15( \a[15] ) , .pi16( \b[0] ) , .pi17( \b[1] ) , .pi18( \b[2] ) , .pi19( \b[3] ) , .pi20( \b[4] ) , .pi21( \b[5] ) , .pi22( \b[6] ) , .pi23( \b[7] ) , .pi24( \b[8] ) , .pi25( \b[9] ) , .pi26( \b[10] ) , .pi27( \b[11] ) , .pi28( \b[12] ) , .pi29( \b[13] ) , .pi30( \b[14] ) , .pi31( \b[15] ) , .po00( \r[0] ) , .po01( \r[1] ) , .po02( \r[2] ) , .po03( \r[3] ) , .po04( \r[4] ) , .po05( \r[5] ) , .po06( \r[6] ) , .po07( \r[7] ) , .po08( \r[8] ) , .po09( \r[9] ) , .po10( \r[10] ) , .po11( \r[11] ) , .po12( \r[12] ) , .po13( \r[13] ) , .po14( \r[14] ) , .po15( \r[15] ) , .po16( \r[16] ) , .po17( \r[17] ) , .po18( \r[18] ) , .po19( \r[19] ) , .po20( \r[20] ) , .po21( \r[21] ) , .po22( \r[22] ) , .po23( \r[23] ) , .po24( \r[24] ) , .po25( \r[25] ) , .po26( \r[26] ) , .po27( \r[27] ) , .po28( \r[28] ) , .po29( \r[29] ) , .po30( \r[30] ) , .po31( \r[31] ) );
endmodule

module top(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31;
  wire n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, tpo00, tpo01, tpo02, tpo03, tpo04, tpo05, tpo06, tpo07, tpo08, tpo09, tpo10, tpo11, tpo12, tpo13, tpo14, tpo15, tpo16, tpo17, tpo18, tpo19, tpo20, tpo21, tpo22, tpo23, tpo24, tpo25, tpo26, tpo27, tpo28, tpo29, tpo30, tpo31;
  assign po00 = tpo00;
  assign po01 = tpo01;
  assign po02 = tpo02;
  assign po03 = tpo03;
  assign po04 = tpo04;
  assign po05 = tpo05;
  assign po06 = tpo06;
  assign po07 = tpo07;
  assign po08 = tpo08;
  assign po09 = tpo09;
  assign po10 = tpo10;
  assign po11 = ~tpo11;
  assign po12 = tpo12;
  assign po13 = tpo13;
  assign po14 = tpo14;
  assign po15 = tpo15;
  assign po16 = tpo16;
  assign po17 = ~tpo17;
  assign po18 = tpo18;
  assign po19 = ~tpo19;
  assign po20 = tpo20;
  assign po21 = ~tpo21;
  assign po22 = tpo22;
  assign po23 = ~tpo23;
  assign po24 = tpo24;
  assign po25 = ~tpo25;
  assign po26 = tpo26;
  assign po27 = ~tpo27;
  assign po28 = tpo28;
  assign po29 = ~tpo29;
  assign po30 = tpo30;
  assign po31 = ~tpo31;
  mult16_0 U0 ( .pi0( n102 ), .pi1( n103 ), .pi2( n104 ), .pi3( n105 ), .pi4( n107 ), .pi5( n109 ), .pi6( n129 ), .pi7( n131 ), .po0( n110 ), .po1( n111 ), .po2( n132 ), .po3( n133 ), .po4( n142 ) );
  mult16_1 U1 ( .pi00( pi06 ), .pi01( pi07 ), .pi02( pi08 ), .pi03( pi09 ), .pi04( pi10 ), .pi05( pi11 ), .pi06( pi16 ), .pi07( pi17 ), .pi08( pi19 ), .pi09( n22 ), .pi10( n62 ), .pi11( n89 ), .pi12( n91 ), .po00(  ), .po01(  ), .po02(  ), .po03( n45 ), .po04( n59 ), .po05( n63 ), .po06( n75 ), .po07( n76 ), .po08( n77 ), .po09( n78 ), .po10( n92 ), .po11( n103 ), .po12( n104 ) );
  mult16_2 U2 ( .pi0( n75 ), .pi1( n77 ), .pi2( n78 ), .pi3( n79 ), .pi4( n84 ), .pi5( n92 ), .pi6( n94 ), .pi7( n97 ), .po0( n85 ), .po1( n98 ), .po2( n101 ), .po3( n102 ) );
  mult16_3 U3 ( .pi0( pi03 ), .pi1( pi24 ), .pi2( n35 ), .pi3( n60 ), .pi4( n61 ), .pi5( n80 ), .pi6( n82 ), .po0( n62 ), .po1( n83 ), .po2( n84 ), .po3( n95 ) );
  mult16_4 U4 ( .pi00( pi05 ), .pi01( pi06 ), .pi02( pi07 ), .pi03( pi08 ), .pi04( pi09 ), .pi05( pi10 ), .pi06( pi11 ), .pi07( pi18 ), .pi08( pi20 ), .pi09( pi21 ), .pi10( n46 ), .pi11( n81 ), .pi12( n83 ), .pi13( n93 ), .po00(  ), .po01( n60 ), .po02( n61 ), .po03( n79 ), .po04( n90 ), .po05( n91 ), .po06( n94 ), .po07( n106 ), .po08( n107 ), .po09( n108 ), .po10( n113 ), .po11( n130 ) );
  mult16_5 U5 ( .pi00( pi04 ), .pi01( pi05 ), .pi02( pi06 ), .pi03( pi07 ), .pi04( pi08 ), .pi05( pi22 ), .pi06( pi23 ), .pi07( pi24 ), .pi08( n108 ), .pi09( n130 ), .po00(  ), .po01( n65 ), .po02( n81 ), .po03( n82 ), .po04( n93 ), .po05( n109 ), .po06( n131 ), .po07( n134 ), .po08( n149 ), .po09( n152 ) );
  mult16_6 U6 ( .pi0( n100 ), .pi1( n101 ), .pi2( n110 ), .pi3( n111 ), .pi4( n112 ), .pi5( n113 ), .pi6( n119 ), .po0( n120 ), .po1( n121 ), .po2( n139 ), .po3( n140 ) );
  mult16_7 U7 ( .pi00( n162 ), .pi01( n163 ), .pi02( n164 ), .pi03( n176 ), .pi04( n178 ), .pi05( n179 ), .pi06( n180 ), .pi07( n181 ), .pi08( n197 ), .pi09( n213 ), .po0( tpo16 ), .po1( tpo17 ), .po2( tpo18 ), .po3( n214 ) );
  mult16_8 U8 ( .pi00( n117 ), .pi01( n121 ), .pi02( n132 ), .pi03( n133 ), .pi04( n138 ), .pi05( n139 ), .pi06( n140 ), .pi07( n142 ), .pi08( n151 ), .pi09( n158 ), .pi10( n160 ), .pi11( n161 ), .po0( n141 ), .po1( tpo15 ), .po2( n163 ), .po3( n164 ), .po4( n179 ), .po5( n180 ) );
  mult16_9 U9 ( .pi00( n114 ), .pi01( n116 ), .pi02( n118 ), .pi03( n134 ), .pi04( n135 ), .pi05( n136 ), .pi06( n137 ), .pi07( n152 ), .pi08( n154 ), .pi09( n156 ), .po0( n119 ), .po1( n138 ), .po2( n157 ), .po3( n158 ), .po4( n159 ), .po5( n177 ) );
  mult16_10 U10 ( .pi00( pi00 ), .pi01( pi01 ), .pi02( pi02 ), .pi03( pi03 ), .pi04( pi28 ), .pi05( pi29 ), .pi06( pi30 ), .pi07( pi31 ), .pi08( n159 ), .pi09( n177 ), .po00(  ), .po01(  ), .po02(  ), .po03(  ), .po04(  ), .po05(  ), .po06( n96 ), .po07( n117 ), .po08( n118 ), .po09( n137 ), .po10( n155 ), .po11( n156 ), .po12( n160 ), .po13( n162 ), .po14( n178 ), .po15( n181 ) );
  mult16_11 U11 ( .pi00( pi00 ), .pi01( pi01 ), .pi02( pi02 ), .pi03( pi03 ), .pi04( pi25 ), .pi05( pi26 ), .pi06( pi27 ), .pi07( n95 ), .pi08( n96 ), .pi09( n115 ), .po0( n53 ), .po1( n68 ), .po2( n87 ), .po3( n97 ), .po4( n100 ), .po5( n112 ), .po6( n114 ), .po7( n116 ), .po8( n135 ) );
  mult16_12 U12 ( .pi0( pi03 ), .pi1( pi04 ), .pi2( pi05 ), .pi3( pi06 ), .pi4( pi25 ), .pi5( pi26 ), .pi6( pi27 ), .pi7( n157 ), .po00(  ), .po01(  ), .po02(  ), .po03(  ), .po04( n115 ), .po05( n136 ), .po06( n153 ), .po07( n154 ), .po08( n165 ), .po09( n166 ) );
  mult16_13 U13 ( .pi0( n42 ), .pi1( n54 ), .po0( n55 ), .po1( n56 ) );
  mult16_14 U14 ( .pi0( n55 ), .pi1( n57 ), .pi2( n58 ), .pi3( n71 ), .pi4( n88 ), .po0( tpo10 ), .po1( tpo11 ), .po2( n99 ) );
  mult16_15 U15 ( .pi00( n69 ), .pi01( n72 ), .pi02( n73 ), .pi03( n74 ), .pi04( n85 ), .pi05( n86 ), .pi06( n87 ), .pi07( n98 ), .pi08( n99 ), .pi09( n120 ), .pi10( n141 ), .po0( n88 ), .po1( tpo12 ), .po2( tpo13 ), .po3( tpo14 ), .po4( n161 ) );
  mult16_16 U16 ( .pi0( n27 ), .pi1( n34 ), .pi2( n37 ), .pi3( n38 ), .pi4( n39 ), .pi5( n52 ), .pi6( n53 ), .pi7( n70 ), .po0( n40 ), .po1( n54 ), .po2( n71 ), .po3( n72 ) );
  mult16_17 U17 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi02 ), .pi3( pi03 ), .pi4( pi22 ), .pi5( pi23 ), .pi6( pi24 ), .pi7( n50 ), .pi8( n65 ), .po00(  ), .po01(  ), .po02(  ), .po03( n24 ), .po04( n27 ), .po05( n28 ), .po06( n39 ), .po07( n51 ), .po08( n64 ), .po09( n66 ), .po10( n67 ), .po11( n80 ) );
  mult16_18 U18 ( .pi00( n43 ), .pi01( n44 ), .pi02( n45 ), .pi03( n47 ), .pi04( n48 ), .pi05( n49 ), .pi06( n51 ), .pi07( n63 ), .pi08( n64 ), .pi09( n66 ), .pi10( n67 ), .pi11( n68 ), .po0( n52 ), .po1( n69 ), .po2( n70 ), .po3( n73 ), .po4( n74 ), .po5( n86 ) );
  mult16_19 U19 ( .pi0( n26 ), .pi1( n28 ), .pi2( n29 ), .pi3( n32 ), .pi4( n40 ), .po0( n33 ), .po1( n41 ), .po2( n42 ) );
  mult16_20 U20 ( .pi0( n5 ), .pi1( n6 ), .pi2( n8 ), .pi3( n9 ), .pi4( n11 ), .pi5( n12 ), .pi6( n14 ), .pi7( n15 ), .pi8( n16 ), .po0( tpo04 ), .po1( tpo05 ), .po2( n17 ), .po3( n18 ), .po4( n19 ), .po5( n20 ) );
  mult16_21 U21 ( .pi00( n17 ), .pi01( n18 ), .pi02( n19 ), .pi03( n20 ), .pi04( n23 ), .pi05( n24 ), .pi06( n25 ), .pi07( n33 ), .pi08( n41 ), .pi09( n56 ), .po0( tpo06 ), .po1( tpo07 ), .po2( tpo08 ), .po3( n57 ), .po4( tpo09 ), .po5( n58 ) );
  mult16_22 U22 ( .pi00( pi00 ), .pi01( pi01 ), .pi02( pi02 ), .pi03( pi03 ), .pi04( pi04 ), .pi05( pi05 ), .pi06( pi06 ), .pi07( pi07 ), .pi08( pi18 ), .pi09( pi20 ), .pi10( pi21 ), .pi11( n3 ), .po00(  ), .po01(  ), .po02(  ), .po03(  ), .po04( n10 ), .po05( n12 ), .po06( n16 ), .po07( n21 ), .po08( n25 ), .po09( n26 ), .po10( n31 ), .po11( n35 ), .po12( n36 ), .po13( n38 ), .po14( n46 ), .po15( n47 ), .po16( n48 ), .po17( n49 ), .po18( n50 ) );
  mult16_23 U23 ( .pi00( pi00 ), .pi01( pi01 ), .pi02( pi17 ), .pi03( pi18 ), .pi04( tpo00 ), .pi05( n0 ), .pi06( n1 ), .pi07( n2 ), .pi08( n4 ), .pi09( n10 ), .po0(  ), .po1(  ), .po2( tpo01 ), .po3( tpo02 ), .po4( n3 ), .po5( n5 ), .po6( tpo03 ), .po7( n6 ), .po8( n11 ) );
  mult16_24 U24 ( .pi00( pi06 ), .pi01( pi07 ), .pi02( pi08 ), .pi03( pi16 ), .pi04( pi17 ), .pi05( n7 ), .pi06( n13 ), .pi07( n30 ), .pi08( n31 ), .pi09( n36 ), .po0(  ), .po1( n22 ), .po2( n32 ), .po3( n34 ), .po4( n37 ), .po5( n43 ), .po6( n44 ) );
  mult16_25 U25 ( .pi00( pi00 ), .pi01( pi01 ), .pi02( pi02 ), .pi03( pi03 ), .pi04( pi04 ), .pi05( pi05 ), .pi06( pi16 ), .pi07( pi17 ), .pi08( pi19 ), .pi09( n21 ), .pi10( n22 ), .po00(  ), .po01(  ), .po02(  ), .po03( tpo00 ), .po04( n0 ), .po05( n1 ), .po06( n2 ), .po07( n4 ), .po08( n7 ), .po09( n8 ), .po10( n9 ), .po11( n13 ), .po12( n14 ), .po13( n15 ), .po14( n23 ), .po15( n29 ), .po16( n30 ) );
  mult16_26 U26 ( .pi0( n289 ), .pi1( n291 ), .pi2( n292 ), .pi3( n293 ), .pi4( n294 ), .pi5( n302 ), .pi6( n303 ), .pi7( n304 ), .po0( n295 ), .po1( n305 ), .po2( n306 ), .po3( n307 ), .po4( n308 ) );
  mult16_27 U27 ( .pi00( pi10 ), .pi01( pi11 ), .pi02( pi12 ), .pi03( pi13 ), .pi04( pi14 ), .pi05( pi28 ), .pi06( pi29 ), .pi07( pi30 ), .pi08( pi31 ), .pi09( n274 ), .pi10( n299 ), .pi11( n301 ), .po0( n283 ), .po1( n290 ), .po2( n292 ), .po3( n294 ), .po4( n300 ), .po5( n303 ), .po6( n304 ), .po7( n312 ), .po8( n314 ) );
  mult16_28 U28 ( .pi00( pi12 ), .pi01( pi13 ), .pi02( pi14 ), .pi03( pi15 ), .pi04( pi25 ), .pi05( pi26 ), .pi06( pi27 ), .pi07( n283 ), .pi08( n290 ), .pi09( n300 ), .po0( n262 ), .po1( n273 ), .po2( n284 ), .po3( n289 ), .po4( n291 ), .po5( n301 ), .po6( n302 ), .po7( n309 ) );
  mult16_29 U29 ( .pi0( n297 ), .pi1( n298 ), .pi2( n306 ), .pi3( n307 ), .pi4( n313 ), .po0( tpo26 ), .po1( tpo27 ), .po2( n316 ) );
  mult16_30 U30 ( .pi0( pi13 ), .pi1( pi14 ), .pi2( pi15 ), .pi3( pi28 ), .pi4( pi29 ), .pi5( pi30 ), .pi6( pi31 ), .pi7( n311 ), .pi8( n318 ), .po0(  ), .po1(  ), .po2( n299 ), .po3( n310 ), .po4( n315 ), .po5( n317 ), .po6( tpo30 ), .po7( tpo31 ) );
  mult16_31 U31 ( .pi0( n305 ), .pi1( n308 ), .pi2( n309 ), .pi3( n310 ), .pi4( n312 ), .pi5( n314 ), .pi6( n315 ), .pi7( n316 ), .pi8( n317 ), .po0( n311 ), .po1( n313 ), .po2( tpo28 ), .po3( tpo29 ), .po4( n318 ) );
  mult16_32 U32 ( .pi0( n258 ), .pi1( n261 ), .pi2( n264 ), .pi3( n266 ), .pi4( n267 ), .pi5( n268 ), .pi6( n279 ), .po0( n265 ), .po1( n269 ), .po2( n280 ), .po3( n281 ) );
  mult16_33 U33 ( .pi0( pi11 ), .pi1( pi12 ), .pi2( pi13 ), .pi3( pi14 ), .pi4( pi15 ), .pi5( pi22 ), .pi6( pi23 ), .pi7( pi24 ), .po00(  ), .po01(  ), .po02( n208 ), .po03( n225 ), .po04( n233 ), .po05( n234 ), .po06( n250 ), .po07( n251 ), .po08( n259 ), .po09( n260 ), .po10( n261 ), .po11( n270 ) );
  mult16_34 U34 ( .pi0( n222 ), .pi1( n223 ), .pi2( n233 ), .pi3( n234 ), .pi4( n251 ), .pi5( n252 ), .pi6( n254 ), .po0( n235 ), .po1( n255 ), .po2( n258 ), .po3( n267 ) );
  mult16_35 U35 ( .pi0( n265 ), .pi1( n276 ), .pi2( n278 ), .pi3( n281 ), .pi4( n282 ), .pi5( n287 ), .pi6( n288 ), .pi7( n296 ), .po0( n279 ), .po1( tpo24 ), .po2( tpo25 ), .po3( n297 ) );
  mult16_36 U36 ( .pi00( n259 ), .pi01( n260 ), .pi02( n270 ), .pi03( n271 ), .pi04( n272 ), .pi05( n273 ), .pi06( n275 ), .pi07( n284 ), .pi08( n285 ), .pi09( n286 ), .pi10( n295 ), .po0( n276 ), .po1( n287 ), .po2( n293 ), .po3( n296 ), .po4( n298 ) );
  mult16_37 U37 ( .pi00( pi07 ), .pi01( pi08 ), .pi02( pi09 ), .pi03( pi10 ), .pi04( pi11 ), .pi05( pi28 ), .pi06( pi29 ), .pi07( pi30 ), .pi08( pi31 ), .pi09( n277 ), .po00( n253 ), .po01( n263 ), .po02( n266 ), .po03( n268 ), .po04( n274 ), .po05( n275 ), .po06( n278 ), .po07( n282 ), .po08( n285 ), .po09( n286 ) );
  mult16_38 U38 ( .pi00( pi08 ), .pi01( pi09 ), .pi02( pi10 ), .pi03( pi11 ), .pi04( pi12 ), .pi05( pi25 ), .pi06( pi26 ), .pi07( pi27 ), .pi08( n250 ), .pi09( n253 ), .pi10( n262 ), .pi11( n263 ), .po0( n200 ), .po1( n239 ), .po2( n254 ), .po3( n264 ), .po4( n271 ), .po5( n272 ), .po6( n277 ) );
  mult16_39 U39 ( .pi0( n214 ), .pi1( n215 ), .pi2( n216 ), .pi3( n217 ), .pi4( n230 ), .pi5( n243 ), .po0( tpo19 ), .po1( n244 ), .po2( n245 ), .po3( tpo20 ) );
  mult16_40 U40 ( .pi00( n218 ), .pi01( n221 ), .pi02( n227 ), .pi03( n228 ), .pi04( n229 ), .pi05( n231 ), .pi06( n232 ), .pi07( n235 ), .pi08( n240 ), .pi09( n242 ), .po0( n230 ), .po1( n243 ), .po2( n246 ), .po3( n248 ), .po4( n249 ) );
  mult16_41 U41 ( .pi00( n244 ), .pi01( n245 ), .pi02( n246 ), .pi03( n247 ), .pi04( n248 ), .pi05( n249 ), .pi06( n255 ), .pi07( n256 ), .pi08( n257 ), .pi09( n269 ), .pi10( n280 ), .po0( tpo21 ), .po1( tpo22 ), .po2( tpo23 ), .po3( n288 ) );
  mult16_42 U42 ( .pi00( pi06 ), .pi01( pi07 ), .pi02( pi08 ), .pi03( pi09 ), .pi04( pi10 ), .pi05( pi25 ), .pi06( pi26 ), .pi07( pi27 ), .pi08( n200 ), .pi09( n203 ), .pi10( n219 ), .pi11( n220 ), .po0( n167 ), .po1( n168 ), .po2( n184 ), .po3( n201 ), .po4( n221 ), .po5( n236 ), .po6( n238 ), .po7( n241 ) );
  mult16_43 U43 ( .pi00( pi05 ), .pi01( pi06 ), .pi02( pi07 ), .pi03( pi08 ), .pi04( pi28 ), .pi05( pi29 ), .pi06( pi30 ), .pi07( pi31 ), .pi08( n236 ), .pi09( n237 ), .pi10( n238 ), .pi11( n239 ), .pi12( n241 ), .po0( n202 ), .po1( n220 ), .po2( n240 ), .po3( n242 ), .po4( n247 ), .po5( n252 ), .po6( n256 ), .po7( n257 ) );
  mult16_44 U44 ( .pi00( pi02 ), .pi01( pi03 ), .pi02( pi04 ), .pi03( pi05 ), .pi04( pi28 ), .pi05( pi29 ), .pi06( pi30 ), .pi07( pi31 ), .pi08( n155 ), .pi09( n198 ), .pi10( n199 ), .pi11( n201 ), .pi12( n202 ), .pi13( n211 ), .po00( n169 ), .po01( n185 ), .po02( n194 ), .po03( n196 ), .po04( n203 ), .po05( n204 ), .po06( n212 ), .po07( n216 ), .po08( n229 ), .po09( n231 ) );
  mult16_45 U45 ( .pi00( pi05 ), .pi01( pi27 ), .pi02( n153 ), .pi03( n166 ), .pi04( n167 ), .pi05( n168 ), .pi06( n169 ), .pi07( n183 ), .pi08( n184 ), .pi09( n185 ), .po0( n170 ), .po1( n186 ), .po2( n198 ), .po3( n211 ) );
  mult16_46 U46 ( .pi0( n182 ), .pi1( n186 ), .pi2( n187 ), .pi3( n193 ), .pi4( n194 ), .pi5( n195 ), .pi6( n196 ), .pi7( n210 ), .pi8( n212 ), .po0( n197 ), .po1( n213 ), .po2( n215 ), .po3( n217 ) );
  mult16_47 U47 ( .pi00( n90 ), .pi01( n125 ), .pi02( n126 ), .pi03( n127 ), .pi04( n128 ), .pi05( n148 ), .pi06( n149 ), .pi07( n150 ), .pi08( n165 ), .pi09( n170 ), .pi10( n175 ), .po0( n129 ), .po1( n151 ), .po2( n176 ), .po3( n182 ), .po4( n195 ) );
  mult16_48 U48 ( .pi00( n76 ), .pi01( n106 ), .pi02( n122 ), .pi03( n123 ), .pi04( n124 ), .pi05( n144 ), .pi06( n145 ), .pi07( n146 ), .pi08( n147 ), .pi09( n172 ), .pi10( n173 ), .pi11( n174 ), .po0( n125 ), .po1( n148 ), .po2( n175 ), .po3( n183 ), .po4( n187 ) );
  mult16_49 U49 ( .pi00( pi10 ), .pi01( pi11 ), .pi02( pi12 ), .pi03( pi13 ), .pi04( pi14 ), .pi05( pi15 ), .pi06( pi16 ), .pi07( pi17 ), .pi08( pi19 ), .pi09( n59 ), .pi10( n171 ), .pi11( n189 ), .po00( n89 ), .po01( n105 ), .po02( n122 ), .po03( n123 ), .po04( n124 ), .po05( n126 ), .po06( n143 ), .po07( n144 ), .po08( n172 ), .po09( n188 ), .po10( n190 ), .po11( n205 ) );
  mult16_50 U50 ( .pi00( pi11 ), .pi01( pi12 ), .pi02( pi13 ), .pi03( pi14 ), .pi04( pi15 ), .pi05( pi18 ), .pi06( pi20 ), .pi07( pi21 ), .pi08( n143 ), .pi09( n224 ), .pi10( n225 ), .po00( n128 ), .po01( n146 ), .po02( n147 ), .po03( n171 ), .po04( n189 ), .po05( n191 ), .po06( n206 ), .po07( n207 ), .po08( n222 ), .po09( n223 ), .po10( n226 ), .po11( n232 ), .po12( n237 ) );
  mult16_51 U51 ( .pi00( pi07 ), .pi01( pi08 ), .pi02( pi09 ), .pi03( pi10 ), .pi04( pi11 ), .pi05( pi12 ), .pi06( pi21 ), .pi07( pi22 ), .pi08( pi23 ), .pi09( pi24 ), .pi10( n191 ), .pi11( n207 ), .pi12( n208 ), .po00( n127 ), .po01( n145 ), .po02( n150 ), .po03( n173 ), .po04( n174 ), .po05( n192 ), .po06( n199 ), .po07( n209 ), .po08( n219 ), .po09( n224 ) );
  mult16_52 U52 ( .pi0( n188 ), .pi1( n190 ), .pi2( n192 ), .pi3( n204 ), .pi4( n205 ), .pi5( n206 ), .pi6( n209 ), .pi7( n226 ), .po0( n193 ), .po1( n210 ), .po2( n218 ), .po3( n227 ), .po4( n228 ) );
endmodule
