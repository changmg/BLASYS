module c7552_tb;
reg [206:0] pi;
wire [54:0] po;
c7552 dut( pi[0] , pi[1] , pi[2] , pi[3] , pi[4] , pi[5] , pi[6] , pi[7] , pi[8] , pi[9] , pi[10] , pi[11] , pi[12] , pi[13] , pi[14] , pi[15] , pi[16] , pi[17] , pi[18] , pi[19] , pi[20] , pi[21] , pi[22] , pi[23] , pi[24] , pi[25] , pi[26] , pi[27] , pi[28] , pi[29] , pi[30] , pi[31] , pi[32] , pi[33] , pi[34] , pi[35] , pi[36] , pi[37] , pi[38] , pi[39] , pi[40] , pi[41] , pi[42] , pi[43] , pi[44] , pi[45] , pi[46] , pi[47] , pi[48] , pi[49] , pi[50] , pi[51] , pi[52] , pi[53] , pi[54] , pi[55] , pi[56] , pi[57] , pi[58] , pi[59] , pi[60] , pi[61] , pi[62] , pi[63] , pi[64] , pi[65] , pi[66] , pi[67] , pi[68] , pi[69] , pi[70] , pi[71] , pi[72] , pi[73] , pi[74] , pi[75] , pi[76] , pi[77] , pi[78] , pi[79] , pi[80] , pi[81] , pi[82] , pi[83] , pi[84] , pi[85] , pi[86] , pi[87] , pi[88] , pi[89] , pi[90] , pi[91] , pi[92] , pi[93] , pi[94] , pi[95] , pi[96] , pi[97] , pi[98] , pi[99] , pi[100] , pi[101] , pi[102] , pi[103] , pi[104] , pi[105] , pi[106] , pi[107] , pi[108] , pi[109] , pi[110] , pi[111] , pi[112] , pi[113] , pi[114] , pi[115] , pi[116] , pi[117] , pi[118] , pi[119] , pi[120] , pi[121] , pi[122] , pi[123] , pi[124] , pi[125] , pi[126] , pi[127] , pi[128] , pi[129] , pi[130] , pi[131] , pi[132] , pi[133] , pi[134] , pi[135] , pi[136] , pi[137] , pi[138] , pi[139] , pi[140] , pi[141] , pi[142] , pi[143] , pi[144] , pi[145] , pi[146] , pi[147] , pi[148] , pi[149] , pi[150] , pi[151] , pi[152] , pi[153] , pi[154] , pi[155] , pi[156] , pi[157] , pi[158] , pi[159] , pi[160] , pi[161] , pi[162] , pi[163] , pi[164] , pi[165] , pi[166] , pi[167] , pi[168] , pi[169] , pi[170] , pi[171] , pi[172] , pi[173] , pi[174] , pi[175] , pi[176] , pi[177] , pi[178] , pi[179] , pi[180] , pi[181] , pi[182] , pi[183] , pi[184] , pi[185] , pi[186] , pi[187] , pi[188] , pi[189] , pi[190] , pi[191] , pi[192] , pi[193] , pi[194] , pi[195] , pi[196] , pi[197] , pi[198] , pi[199] , pi[200] , pi[201] , pi[202] , pi[203] , pi[204] , pi[205] , pi[206] , po[0] , po[1] , po[2] , po[3] , po[4] , po[5] , po[6] , po[7] , po[8] , po[9] , po[10] , po[11] , po[12] , po[13] , po[14] , po[15] , po[16] , po[17] , po[18] , po[19] , po[20] , po[21] , po[22] , po[23] , po[24] , po[25] , po[26] , po[27] , po[28] , po[29] , po[30] , po[31] , po[32] , po[33] , po[34] , po[35] , po[36] , po[37] , po[38] , po[39] , po[40] , po[41] , po[42] , po[43] , po[44] , po[45] , po[46] , po[47] , po[48] , po[49] , po[50] , po[51] , po[52] , po[53] , po[54] );
initial
begin
# 1  pi=207'b101111101110100000010111001111001000001111001001000101111000100001000110100101110110111111001111110010100001111101010100110110000001110011100101110111111101000011110011000010001111100111100010010010010011001;
#1 $display("%b", po);
# 1  pi=207'b100100100110101001000101111101000011100101001100111101101100110011001001010010001000001111001101011010100100101001110010001100010101101100100000101101101100101011111010111001011000110001111101111010111100110;
#1 $display("%b", po);
# 1  pi=207'b110100110110001111101001111011101111000110011101011011011110010011011001110101101111010110001100100001010110010011111011000011010110001110100001010100001101100011011101111010000011010000001110000010100100010;
#1 $display("%b", po);
# 1  pi=207'b011100111001111001110101101000011101110100101001011000111001010001101011110010011111010110101101101011010110010100111100010011000011110100101110110110100111011000110110111000111010111011000000010101001110001;
#1 $display("%b", po);
# 1  pi=207'b011101001100000101101101011010110001011100001100001110010011110111110000101100110110101110011110011101001100001011101001100000101111001101011110101101000100110010001011001111001101111000111101110011011101101;
#1 $display("%b", po);
# 1  pi=207'b100111101101101000111010110101101000010110011110110010001011110011101111110000100010000111110100011010100100011111011000110101000010001000010000100110111001011101110110110111111111110001110101001101010001000;
#1 $display("%b", po);
# 1  pi=207'b011100010100111010110000101110110111000001100011011001101011011001100001100101110011011101111101111001011100010000011100011010101010001101100000100101011001100001001110000101100010001110100011001001110100000;
#1 $display("%b", po);
# 1  pi=207'b001010101001100001101111000011100111110100011110100000111101001100100100100010110001110011000100011011100000001011101110010000110011011111000011011110001100101100101011101101100011011110001111001000000001001;
#1 $display("%b", po);
# 1  pi=207'b100111000110010101011101000100001001011001110101000000010000100011011010101111011001001000000110100111010011101110010011000110010010001000101110100011011011001011001010110110011001000011000011110100000101011;
#1 $display("%b", po);
# 1  pi=207'b100100111111000110000100000001000010010000110000100100100100101100001101011010100100111110011001011011111011111110111101011111100000000001000000100101100111111001001011001110110111000100011111101100100011000;
#1 $display("%b", po);
# 1  pi=207'b010111111000111110101100001000101011111011010101010011100111001001001100100010010010101010000010110110100101000101101000100101101011000010111001101100010000010010100000101111011110110101100100000111100101101;
#1 $display("%b", po);
# 1  pi=207'b010011001010011110111110111001010110111110000110101100110110011101101111101010100101110111010001011010111110101001100110000110000100100111000011111100110101111011000111101000101010100000000000001110110111111;
#1 $display("%b", po);
# 1  pi=207'b000010110001000011110100110001000100101000001111111010000011001010110001010110001000110111010101101101001000111011110111111100001100001001001111111001011000111101110100100100001000111010111111110100011011100;
#1 $display("%b", po);
# 1  pi=207'b010100111001000011001001011000100010011010100000001010000000111011110010011110001101100100110111100001111011000101111100101001100001111101010101101101011100000010001011010000100110100000001010100110101100111;
#1 $display("%b", po);
# 1  pi=207'b110010001101000101010001001010000101100001101000101110111100011001011010111001100110100011001100010111100000101010010100000100011010111001101001100011110100100110111110111001110000000110110110000011101110111;
#1 $display("%b", po);
# 1  pi=207'b100011101001000011111010001001010001100110101110001101001010011100111100001000110100011111001010111000011011011110101100101000110101000000001000001101011111100100001110101001111001001101101001010111110110101;
#1 $display("%b", po);
# 1  pi=207'b111100011100000110001100001110111100001011000010111010000101111110011101100010110111100110100001101011000110101101100100100000111111011111001000001101100001100011010011011011011010111011001011110110111001001;
#1 $display("%b", po);
# 1  pi=207'b111100000000010001001110100011101010010101000000011010011100001101111110011001000000011100000111100101011100110110111111000011000000000000100010000110110111000011011011110011101001110000101111011011000100010;
#1 $display("%b", po);
# 1  pi=207'b001101011001001000010111011011101011110100101101100001000111110100000111110100111001001111101000110111001010011011010001010001011100110001010101011011101101010001101011111011000101111101101111011010110010011;
#1 $display("%b", po);
# 1  pi=207'b011000111100110000100001011101010110010111110011110101011101110000000100100010101111001100001111110110000111110010011111011010111011111001101110010110000000111100111000000000011000000001111110001101100011100;
#1 $display("%b", po);
# 1  pi=207'b100100011010110111000001010000001100110100000101010110110011000011000010110000011100101110010101000011010111010001101100011010100100101010100100011100101100111101110001111001010010000010111001110010011011100;
#1 $display("%b", po);
# 1  pi=207'b101001100010110010111100011001011111111000100000101010110000101100110111000101101100100101000010111101000111001000101000011010010001101101110010101000101101011111110001110101000100011000000001011111000000111;
#1 $display("%b", po);
# 1  pi=207'b001110110111001010110000111000010001001111010111101111100111100011100111101100010101001111101111010110101110010011111101000011110100010111011110110101100100110000000111010011011110000010010111011101101110100;
#1 $display("%b", po);
# 1  pi=207'b100110000111010101101100100011100100110101010110100000111101011110111011010101001100011001000001000001011011001000000100000001000010000111111010000001010111001011011111010010110110101110101100111011000110010;
#1 $display("%b", po);
# 1  pi=207'b100101000110100010001111011010101100111001001010111001000101011110011001010010000111010101100001000100110010111110111011100011001010010001100101000110000010100101000000000101000100100001010010011000010011010;
#1 $display("%b", po);
# 1  pi=207'b100110111111011010100100010010000000100001000011001001110000111010101000000001000101100001111000100110001011001011001111001110111100110011100010000101010111100001011011110110100111001111110000011110011111011;
#1 $display("%b", po);
# 1  pi=207'b111011100010011001000001000001100000111100100101111010010111110000101100100100011101011110010011010100010101001110111111000100101010011110110000100111011010110000000010010100001101100100110100000011010101011;
#1 $display("%b", po);
# 1  pi=207'b110101100111101010100001101101001010111101001001001111001000010111100001111110111110101101000100110000011011010010100000100010011111011000001111110011100110101000110101011001101100001001001000001010010010011;
#1 $display("%b", po);
# 1  pi=207'b000111111011001000010110000000001100000101010110010110101100100010001100000011011000000011101100100101110011010110010010101011000011011001000110111010001001001111101011010010011010000010110001001101110001100;
#1 $display("%b", po);
# 1  pi=207'b100100110011010011100011001100011111011100101011100110100111100111100011011110001111000100000101011000011011110100111110001101011101011001011001000101110110100101111100100011100100101000011111111100100110001;
#1 $display("%b", po);
# 1  pi=207'b000110110001011111010010111111101100010110111001011011011010010100010001110000001100111010010101010100010110111110010101110000100100100010110110100011010001000010100001110010010111101010101010010001001011100;
#1 $display("%b", po);
# 1  pi=207'b010011010000101011111101110010100000000100101100010010101101000001010110110111000111011101110010110011000010000100110001010001001101110101101110001101110011101001111010111001110101101000000110001000100000010;
#1 $display("%b", po);
# 1  pi=207'b010110000000010100110110010000111110110000001010111110101001100010011000101111111010101010000011110111000110010000011000000000110011111001110010001000101110111111001101111111100101011100111000011010000011010;
#1 $display("%b", po);
# 1  pi=207'b101100100110100001001101101001001110001010101001011110000100001101100011101110100111010010000010010111010110101001100100010101110011001001110110100110100100001100111100011000010001011000101010010010110010100;
#1 $display("%b", po);
# 1  pi=207'b000010101101111001011000011110100110101000110010000111100101011001110001011010110000010111001110100001111000101001011011111001101001001001110100110101010110101111000010001001111001100100110001010011101110001;
#1 $display("%b", po);
# 1  pi=207'b000111110111000101010011001101011000010001001111110000100011011110100110110011111101001010101100111010001011111101011111010100001101000100001100110011011110110111000001100010111101010111011101101001111101011;
#1 $display("%b", po);
# 1  pi=207'b111110100001001111100100011010101011101110111111000001001111111111100100000111000100010101011100110000001111100001010111000010111111111010000111011110000001111110011001110000011010110011100001111110110111110;
#1 $display("%b", po);
# 1  pi=207'b001110000101110000011000100110110011001110011000100000111001111101101010111110101010010000011001001111110111101010000001010100111011010111000110101101011111111010000001110000000110000110011111000111001001111;
#1 $display("%b", po);
# 1  pi=207'b100100000101000111111001011100001011000001101110000010110100011100100011010100000100010111010010011001001010010000111010101111101111001010100100011110011011010100110010001001011011010111001011100000011000101;
#1 $display("%b", po);
# 1  pi=207'b101001001001010001010011101011110101110001111110001010111000101001100000010111001101011010000010010000011001100001010001011101111000101010100011100010010011001100110101010011110010100111001111000000101000111;
#1 $display("%b", po);
# 1  pi=207'b011011100011111101100011111000100001010100110101110000100001110110101101101100111000000001010100111000001111111111001101111011010110111100101001011110011111100000100010010001111001001010100001110110011111101;
#1 $display("%b", po);
# 1  pi=207'b000111100000011110110011111011001000000110001000000100000011000000100010101011001000011101011010011110000001011001100110100001110100010000101100101010110100011110011110010011101010001100110111111000110110000;
#1 $display("%b", po);
# 1  pi=207'b011100010010101010011101010001010010111011010101111011011101010100101110100100110000101110011011111010001000011100110001011011011101100010111110100111110000110100011110010100100111110111001111110010101110000;
#1 $display("%b", po);
# 1  pi=207'b111110100010110110110011101000001010101000001100001010100111000101111001101011100001100110110100001100001111001010100001101001010001110101100010011011010011100001011101111110100000100111001101111001101001001;
#1 $display("%b", po);
# 1  pi=207'b110101001111110001111000011000000110011111100010010001010101001110110001110100001110100100101101011101010000101001111101001010110000111001100011110000100000010101101110100010101100000110100001111100010010100;
#1 $display("%b", po);
# 1  pi=207'b010111010010010011011011010111000101100001100100100001000101110110010110110101010100001110000010001011010000100010111001111111011001100001111101101011101001110110010011001111011110011010110001101011000100000;
#1 $display("%b", po);
# 1  pi=207'b000101000000011111010001000000101001100101100100100000111110111000000010101010100000110010000101110010111011011011111000111010100001010101111101110100011111000110010000110011000111111110100010100000000100110;
#1 $display("%b", po);
# 1  pi=207'b000011011100001100110010101000011000000000110001010011111010111111010101011110101110010110011000010101001111001111111111010011001000110011011111010100011001110110110011011011000011010111011111110101111001000;
#1 $display("%b", po);
# 1  pi=207'b011001111001000000000101100001100011011110001101010101010001001100011001100001001000111011101110000111011001011010110010010110101110111001010010101110010101110011101000001000100101111100111010011011100101001;
#1 $display("%b", po);
# 1  pi=207'b000101000110000011111101110000001100000001111011010111101001111011101011100000100110110010001101001011100011101011010100100100000010111100010100001000010111000111001111110111111011001110100111111110101111100;
#1 $display("%b", po);
# 1  pi=207'b111010100100000000010001110110100111010111111110001011010001100000001100101100011010110010111001001110101101001101011101100000100011000001110010001001001001010110000001110000010110100001110101110111100010110;
#1 $display("%b", po);
# 1  pi=207'b010111001011001110110001110010001101110010001110110100000010101100101010001011010011110101110010010100010010101111110001110111110110110111010101110011000110010011110011010000101110001100010111000001011011111;
#1 $display("%b", po);
# 1  pi=207'b101101101010010101010110110011110001011000000110110110100110000001100111110110001001010000000100010011100101110001001011011010000010110111110011010111000101111010111000101111100010000101010110110000000010100;
#1 $display("%b", po);
# 1  pi=207'b010111001000110101111001000000001100111011000101001001110111111010111100100111010000000001111011100110100101111011000110100000001001000011010010110101110110111101101000101001110101000101000111011110000001111;
#1 $display("%b", po);
# 1  pi=207'b100110110001101000000001100111111011000001010011110000111110001111011101000101011101011001101011110110011110000010110101111011010110111011111110011010001110100000110000000010000100010010010111001001011011110;
#1 $display("%b", po);
# 1  pi=207'b001000100001010110101000111011001101100011110001100010001110001101010001101111011111000111001111001101000010001101111101011011010100000000111001001100101010000010011100100001000101111011100001111100111001000;
#1 $display("%b", po);
# 1  pi=207'b110010001101100100101001110101001001110011010011100001111001000111011011000111110001001100010110000000011110101110000110110010001110001111111101011010001011111001111001111111100110101000111011011101100011101;
#1 $display("%b", po);
# 1  pi=207'b011100101100101101000011110110001010100010011011011100100100000101001010001000011001011110001000011100000010100100100101011100111100001111000010011110011111010000110001110010001001000000110101101001011111000;
#1 $display("%b", po);
# 1  pi=207'b100100000001101100000000011010011110000010011101000010010101011101111111001001100001110011000011111010100101001001101101010101000010010010100011111100100110110010110010101010011010110111100000110000001110010;
#1 $display("%b", po);
# 1  pi=207'b101111100011100011000011100110010010100000000010101011110101100111111000010010110100011000001010011111000011010010101010100101111001110011010100001001100110011001100010101100000001110100110001011111010001011;
#1 $display("%b", po);
# 1  pi=207'b000110101101001101011011101101100011110100010111110100011111101111111001101110110101001111100011001101011111011011100011110010101101111101101011100111110100000110101110000100101001011111011010110001100001011;
#1 $display("%b", po);
# 1  pi=207'b001010011101010010010100110101100111010100101101001011101101011001101111101100111110111011100111000100010010011011010001000111000111100100110010110101111101100100100110001101001010011100011000000000110001001;
#1 $display("%b", po);
# 1  pi=207'b011100100111001001000011011101011001100100101011111101011110000010010010100001110000011000000000010010001010111100011010000101111001101001010111011001111110010100100010001101011011110101011010111001001000011;
#1 $display("%b", po);
# 1  pi=207'b111101000110010000101110011100010111000100000111000001111001100001101011110100100111001011010100111101011000011101100001100100000101001100101000110111101011010101010011010010101001111000111111110100100010001;
#1 $display("%b", po);
# 1  pi=207'b101011101001101011000001110111100110110111000000010011010100000111011010000111101011100110111101110001001011000101011100011000100001110111001110111001110010111100111101100000011011001100100101111100010110110;
#1 $display("%b", po);
# 1  pi=207'b000111001101000011101011011101011000100011111011000011000010000011100101010000111100000000011101001100001011100101111011000001011010011100000101011010100010100000000110100010000010110001010000010100001000011;
#1 $display("%b", po);
# 1  pi=207'b000000010111101101010111101100001100111101110000010010000010101001011001011111101110011110000001111111111001011001101101111011100010100011111011000110110011110001100010100011101001011001100010101000001101110;
#1 $display("%b", po);
# 1  pi=207'b010010100101000010010111011101101001110111100110111110000010101010010000010000100011011011000000001110110100100011001110100001011000101011101010000001110101110101011101101010000011010000111011101010000101010;
#1 $display("%b", po);
# 1  pi=207'b111010100010111101000001100100011111110001111001011000101100001001000100010101000111101011101000001010100101100000111010010011010110011100101110010101001101001000001011110010100111000110011110001001010001111;
#1 $display("%b", po);
# 1  pi=207'b101110000001011010110001011101011010110010001111010000001000010100101000001110001010111100100001010101110110100001011101100111010000110000011110100001100101011010110000111011110110100001111010001011111010101;
#1 $display("%b", po);
# 1  pi=207'b010001011011000000010100011110100100011001101000010110011010101110101110101011011011101010000000001100100101001110000101010011001100100111111100011100001001110011000000001101101011110101100101010110111011001;
#1 $display("%b", po);
# 1  pi=207'b000000000110100001011011101001010010101100110000010000001000010010000101110011001001000011001100011101010000100110001111101110001010000011100101011001100101111011101000111110101011011010000111000110011110101;
#1 $display("%b", po);
# 1  pi=207'b011111001111010100101110001001100111100011011011010011100101110001110111111111101101101101100111000001110011100001010110011100111000001000000000010100010001001111011100011001101101101000111000010101000101010;
#1 $display("%b", po);
# 1  pi=207'b110110011000010011001000100000000110011111110000100110001110001000000101011000010011001101000000001101010100101100111011101010001101001011011111011011010110100000101100010100111110001100001110111101110011011;
#1 $display("%b", po);
# 1  pi=207'b100100101011010100010010010001110011000101111010111100011100111000101000011001011101111000100110100000111000000111000101100011111100001010100011100101010011100001001010010001000110001010001000011101011100100;
#1 $display("%b", po);
# 1  pi=207'b010010011100110011001001000010111110001111010100101010011111011110101110111011011010110010111001010110101101000101100100000100000101110001110000010001100011101010110000101111111011101010101001101010010100000;
#1 $display("%b", po);
# 1  pi=207'b000100010001100000111100101010011111100011010011000100001111011111010100111101110001101010111000011010011001100111100000000011000111110100111101000000111011010011001101111010001110011010101110000001001111111;
#1 $display("%b", po);
# 1  pi=207'b101010111010010010000000010111000100111001011001001100010010001110000111001010110101100010111001011110001110110110100110110100011110000101100001001111100111010100000101001000101010010011110110111011010011000;
#1 $display("%b", po);
# 1  pi=207'b101011001101001001111001101110011111001010111001011100010001010110011101101011011010000100000010101011101001111010001101110110011100001101010101100011110011110001001111010110011101111010001001000000011000001;
#1 $display("%b", po);
# 1  pi=207'b110100100010001010001100000011010011101011101011100110111010010001001101011111110111011100010100101011000101111111000101001111011101000110001110001000100100011101000100101100011101001101001100111011011011100;
#1 $display("%b", po);
# 1  pi=207'b000010001100100100111010100000000011011110110001111001000000101010001011010001100101001101000000010001011000110000101110011001111111000100111000110110110100110100001110101011000111110000001011101010101100010;
#1 $display("%b", po);
# 1  pi=207'b010111010110111010001000110011100000110100101110111010111110001111101100101101111010110111011111100001001111100001101111100011000000101010110011111001111001010101010001000100101000100011000010000110110111001;
#1 $display("%b", po);
# 1  pi=207'b110111010100010000110010110001010010110100110011001001100101010111011000001100001100011010110001101001110001101100100101001000101010000010100010101100110011111101011011000011101100100111101001111011101101110;
#1 $display("%b", po);
# 1  pi=207'b100001110001000001000000110101100100001011110010111000011110100100010110000111101010110110111011100110101101001000000000110010010001110010011011000110000100001111001100001011111011100010100111100001110100010;
#1 $display("%b", po);
# 1  pi=207'b001000010100101100010001101100110101110011010101011111001101011100100000110111000100010110010010111110011010111010000110100100001110111011110111111011000001100011001011111101101101101101110000100100100110100;
#1 $display("%b", po);
# 1  pi=207'b101111000000000111100010000000010101101101110100000101010011101111001111010010110111110111101101011000101111101110001101011101011011100001111110000110001111011100001110010000101001011101000110010110110000000;
#1 $display("%b", po);
# 1  pi=207'b011111111001001100110000011100110001100001001101011001110111010110110101010100011001110110000111111100011110000111111011100000100100011001101010010000010101001000110010111010011011100111110101001001110101000;
#1 $display("%b", po);
# 1  pi=207'b110111011101111101111100001100101000010100111100110101000000010011011101110001101101101011001110011100111011100000011110001010011011010110001010111000011011101010001111000101101110001011111011110110010011010;
#1 $display("%b", po);
# 1  pi=207'b011110000011110111011010100000011011000111101101000010110111011001110010011101111001101101011010100100011111111001001101011100101001010110110010101101111001100001101100101001100011110110110001011011001110101;
#1 $display("%b", po);
# 1  pi=207'b010001110100001111011011110010001010101000100011111110011101101011001110100000001001001111010011100000111101011000010010101001011111000111011000100111110000001000110001101111010111100111100110010010110001011;
#1 $display("%b", po);
# 1  pi=207'b101001000100011001011110011111000111111010100000001000011101011100111011111001100111000100111011001011110011001100101100010000010011110111101010001111101111011001001110001111000100010000000100101111010110100;
#1 $display("%b", po);
# 1  pi=207'b010000111100010010110000010011110111011001011100110111000011110000101111010010011110001100100001001100010000111010001011000101000001010111011101011000110100101001110111111101001111101010010100011101100100001;
#1 $display("%b", po);
# 1  pi=207'b010110010010010111010111111110110011011110011010011010010100011101011000000111111111011011000010110010100100111101110101100100100111011000100101101001100011110001000000010001111101011011011000100100110000001;
#1 $display("%b", po);
# 1  pi=207'b000100000111111100101111010110000011010011101101000110011110010110001011001010000001011010110101011010001111000001111101100011000110000101001111110100010000001100010111001001001111101111000110110000101110110;
#1 $display("%b", po);
# 1  pi=207'b110111110000000001010101001110111000000001011000000000000110100110000111011011110100000000001001111101011111111010011011010011011110001000100010110111101011110100101001100100100000111000100001100001101111010;
#1 $display("%b", po);
# 1  pi=207'b101110100001110010110111110000000101111100100101100001000010011111011011110011101101100100001101110110011000101110101011000001101000000010110111101110110110011001010011011010010111010000000010111000000001010;
#1 $display("%b", po);
# 1  pi=207'b101010110110110110000001011001101001011110001011010001110000000111001100100011000000001010101101110000101001111101001011100001011101110100101101101001000010111010101001010000100011101101111110001110001001001;
#1 $display("%b", po);
# 1  pi=207'b000000100011010011000110000000001111111000111110011001111001010110001001101111110110101001110000110101010000111110111001100000010011101011100111000010101011011101010101110010011110110111001111100110101000111;
#1 $display("%b", po);
# 1  pi=207'b110100001000100111111001011011010110011011110101011111100000011110001000001101111100010101110111110101110110111010001001111010100001111000111100111111110011101101011111110111111111110110001010110000001110100;
#1 $display("%b", po);
# 1  pi=207'b000110000100011111110010000001111011011000011011011110001110100010111110010100000100011011010110001001100111100011000111011000001011001101000101000000100101110100101110010000101111110000100101110110000100011;
#1 $display("%b", po);
# 1  pi=207'b011000000000010100000111011001011000000001011111011001111010000011001001010111101100100101001011101111100111011101111101011101100011011101110100010011011101100000100000011101101001010101011001101101110001100;
#1 $display("%b", po);
# 1  pi=207'b001000001011101101000100100101000000000011100110010100110110111010010101110101101100110011110110010011101111011101000011001000011101110110011000110010001111111101101100010101010000110101100011111101000011101;
#1 $display("%b", po);
# 1  pi=207'b010010110100110001111101100110110000011100000101100100101100001110011101101110111001011100011011001000010101010010010001111111011101101001111110110000011100110001000101101101000011011001110000111101101000111;
#1 $display("%b", po);
# 1  pi=207'b110011000101011001000000101111110010111100000011011011111101111110110000110001010101101110110100010110110110101101111111011110101100100101101101000010101000100101001110111100011111110000001011101010000000111;
#1 $display("%b", po);
# 1  pi=207'b111010011000011001000011001011111100001011110111010000000010000101111100010100100101111110011101001111010001010001010101111011001000111101111100111111010111110110011010101100010101010001100011011011100010011;
#1 $display("%b", po);
# 1  pi=207'b101011101110011011110000000101000110011100001010101110100111000011001011010111011001100001010001101000011111101101011010111001010111000110101100110011110110011110111001101011001000010010110011000001111100010;
#1 $display("%b", po);
# 1  pi=207'b110101011011111100110110101111000001011100100111100100101010111100110100111011111110100101111111110000001101100001000000000000111101001111011100001001111110000111100110011010110101000011001000010111011001001;
#1 $display("%b", po);
# 1  pi=207'b010000001010101110110101000101001011111100111101011001111111110110000001111111011000110010011011110100010001100010101001000010101000001100010010001110100110001111111101100010100101001010001011101010011010011;
#1 $display("%b", po);
# 1  pi=207'b101101111010001010111100111111100101110001010000111011101101000001011010011011110110100001111111001010001101010011000100011111001011101000100000101011001101101111100100100100011100000100110011010000100111000;
#1 $display("%b", po);
# 1  pi=207'b101011001111111101101110101101101001011000101111111010010011001111110011111111110100100011100010011110101101110110011001101101010000111000011101001010111000000111111001101101101110101110100001011000101101101;
#1 $display("%b", po);
# 1  pi=207'b001101000101111110001110110011000100001110000111011110011101101010100010101011111111100011011011110101100001001111100101011100111010010001111001101000110000111010111100111011101100011101100001110111010101110;
#1 $display("%b", po);
# 1  pi=207'b001110100101000010011010111101101100000000000101000100001101011000110100001010011000011001001111010100110101100110100011000000000010000100100000011010101100010010001000101101000010011110110000100111001111111;
#1 $display("%b", po);
# 1  pi=207'b100001001101110010100001100111100010101000010010000101010000111000111110111001110011011000100110001000000100001111010100010100100100110001011010010100101110000001000011011011100011101000101010100111111011110;
#1 $display("%b", po);
# 1  pi=207'b111000101010011111011111101101111111110001000011000100010000101100010101000100110111011100010010001111101010100010110001001100011111000001000111000101101110100001111110100111100110101101010000110001101000000;
#1 $display("%b", po);
# 1  pi=207'b110101010010000011001010010011010100110111001010000000101111001101100111111111100101011110001010110100111011001001011010101011110110001010000011000110000100010011000000011001111001110100011111011010111110010;
#1 $display("%b", po);
# 1  pi=207'b110111000110011000011011011001010001110101011011101011100111010101011000101001100000110011110111111001001110000000101000100100001001011000010010110000100001010110110100101111100110000111101100111011111001001;
#1 $display("%b", po);
# 1  pi=207'b011010010000100011100010101101000101011110000011000000010100110011110101001111100100011000010011101010111101001101001001100101100111001010100101101110111001101111001001101100000001101010101010100101010000110;
#1 $display("%b", po);
# 1  pi=207'b110100000011100011010000110000100100000010111000010100111101011001000010001001011001010101011001100010110011111000101111111100001111000011100000011110101000011011101001100111010110010111100101001111110101111;
#1 $display("%b", po);
# 1  pi=207'b000110101111010010001111000001110101010011010000000111101011000111010000110011100111000000100011110010010010111010111001001100010001011101111010110000110001010111111010001100101011101100100111010110001110110;
#1 $display("%b", po);
# 1  pi=207'b100000111010110101000110111011010001010001010010010101011000111011111111000011001000010101100001011110110000101100111000001110101000001110111000010011011001110101001000010101000111010010010001110001000100001;
#1 $display("%b", po);
# 1  pi=207'b000001111101011111110110111101101100000001101000011001111000001000110000110000000111100011100101010000001111010111101111111000110101101001100100111000110010011001000010100111110111111001010001011000000111111;
#1 $display("%b", po);
# 1  pi=207'b111101011010011000111011111101001110010011000110100101010001100011010000010100001010111100101100100010010010001010011000101101101001010010011010011110010011101001010110111110000011110100101000001001110110110;
#1 $display("%b", po);
# 1  pi=207'b111111111000001100000011100111011110011011010111110111110001101001001001101011010010100000010011100011101011101001100110110110110110110011001000111110000001100101000110010111101101111100011001101001111000111;
#1 $display("%b", po);
# 1  pi=207'b111000010000011000110011001011100110000100011010010011000100000101000100100001111000000000110111100001001010010000100101011111101000001111001000010000111000010111111110011001010100101101010101111001110100000;
#1 $display("%b", po);
# 1  pi=207'b011110011001000001110101100011001101000011000010001011111010010001010010000110110010110000011101111111110111110001001100110101000001000100000110000011000110010100001111110010010000010110101111101010000000010;
#1 $display("%b", po);
# 1  pi=207'b011001001101011101001011001011000101110111111101100000110111010011000100000001010100010011111100101110000101110001100111101011001010100100000100111110111001010110111101101000101111111000010100100010111010111;
#1 $display("%b", po);
# 1  pi=207'b101111111110000001010000101101001111001101101011101101011010010010100001001011001101000101101011011101010111001111001010001101100101011100000101100110110000101010100000010111111001000110100101001111110111011;
#1 $display("%b", po);
# 1  pi=207'b001110110010000010111100100110110100110100110001110000010100011110100011010001001100100101000001011011111100011000100010011000111000111111100110101100010111001100011101010110101101111100011111110011010110100;
#1 $display("%b", po);
# 1  pi=207'b110010100101001000110101100000001000010111110111100001100001110010010101111001111110100100101100000011011111001101000000110110001011101011011101000110001011010011100110011111011001000010100011000011110110111;
#1 $display("%b", po);
# 1  pi=207'b100011010010011101100100010110101011001100001111101001000111111010000000101011111111010100101010100110101101001111001010001111011111011001011000111100000000011000000100000111011111010110111101000111010000100;
#1 $display("%b", po);
# 1  pi=207'b011110111000101011110110000001111110110000010010011110001001111001111101011010100011011110000001100100110110101000100000010000100101110000110010100000011011000111101110001110001011010111011110111010001000111;
#1 $display("%b", po);
# 1  pi=207'b111111101111011011100010111101011010000101111000100100111110000110101110000101100011100101010101010111000111101101110010100101100101011011100001001100110110111011000100010001001110100001100110101011010000010;
#1 $display("%b", po);
# 1  pi=207'b011011111011110110111101001110101100111001111001100111001000000110110011100111001001111000111111001010011100011110010111010111011001010001011010011100001100011101011000001101000101000000010000000110001011001;
#1 $display("%b", po);
# 1  pi=207'b110000100001010011101100001010111001010010010101001010101110000100110110011000000000010100001101100110011111111000010101100011001110001001101000011010111001100101001111010001001001110001111100000001011010001;
#1 $display("%b", po);
# 1  pi=207'b011111010100110101000001100110101001100101111100110110010111010011110111010011000010110101111111000101100000011000100011110110111100100100011011111110100001010001111011101010101010101101110110001010010110101;
#1 $display("%b", po);
# 1  pi=207'b011010101001100111111010111010011101110011100101100101100100101001100010001010100011001010001000110001100110100111110010011110000100110100101011001110101101011010010000101001111010100010110011110111010010001;
#1 $display("%b", po);
# 1  pi=207'b000010011000001001110001110000010100111110010011011110010100101100010000011101101010011000111110111011111101011010001000001011110111001000110000011000101001101111010011100011101111111001000001001111101011000;
#1 $display("%b", po);
# 1  pi=207'b111010010000000110001111011011001010111010000001101100011100010110001001111110000011101110111000010011111110010110010010110111100010010000111100101110101001000011001111000011100010000101001010000000100000111;
#1 $display("%b", po);
# 1  pi=207'b001100010001010001100011000001011011000001111001001101110010110101010101110010111100110011000111010011111110010101101101011101010101001011001001110011011100110111011001000000011001011001011010111011011111101;
#1 $display("%b", po);
# 1  pi=207'b011100011110000111101111001011011010101001101110101101001001010101111000011010110010010110100011110010111001001110110011000010100011100010101010111011110110110001101010100110100100010111011111001000111111110;
#1 $display("%b", po);
# 1  pi=207'b001001110001101011000011111000100010110101001001111000010010000011100000011000110101111011100101101000001000010000011100110010001101100101000010001101111100011010110001100001000101001000001001100110111011001;
#1 $display("%b", po);
# 1  pi=207'b000100110111000111000010000000111110101101000010011000000100101111010101010010010000110000001110011011101100011101111110000001001010100110011101101001001001000001011111011001010100101101001011101001000000111;
#1 $display("%b", po);
# 1  pi=207'b110100111111010010110010110001100100011010000011111000100111111100110010001011001011110101101100100101111001000101011110001111110010110101000110001011010010100100010010110011011110000011100011011010110100010;
#1 $display("%b", po);
# 1  pi=207'b011011011011010000111101110110001110000100101100101111010011001100111011100110100011100011000110010010010100011101000111101110010111000001011010010000100010110010101110010001100001100110110011100001111110100;
#1 $display("%b", po);
# 1  pi=207'b010010010010101010011100001011001111011101101011111111000100101010011000101000100100010010001100100001011001011110111111001101001100101000101111010010100111101111010000000110111110010011110001010110100110011;
#1 $display("%b", po);
# 1  pi=207'b001110100001110111111110110111110010011010101110111001100010111101001111110000101000001100111100110111111010100101111100100001101001100101000100111001000000001011111110001101100110011000110000101110101101111;
#1 $display("%b", po);
# 1  pi=207'b001011000101010100111100010001111100001101010001100110011001010100010001101011111111110101101101110110100011000010100010110101011010100100011001001110001101001111101010001111010100011010000111011101000100110;
#1 $display("%b", po);
# 1  pi=207'b111101101111010001010011010010110110101001000101000111110101111011100000000000010001011011101010110010000101110100110000010101000000110110000011111111000000011110110100111111101000110100001100110011100101100;
#1 $display("%b", po);
# 1  pi=207'b110111010011111001111001100000011011100011101110000110010110010001011001110100101010000111111000100111011000101110001001110001110100111001010011101011001011000110010111010101010010010011100010001001100110001;
#1 $display("%b", po);
# 1  pi=207'b110100110000000111010100010001100011000011100110010101001010000000110011000000000111110011001001101000111001010000110010111111000111000101001010101111110000110010001000001000011011001110001011001001000001000;
#1 $display("%b", po);
# 1  pi=207'b011001110000111010101011000111001011111000000101001100011100000001100100011000101111010011001111001011010010001011110100111111011010111001101111010000010000110001111001101011100001000010010010000111110011101;
#1 $display("%b", po);
# 1  pi=207'b100111011010011000111100111111111110101010111100110111101000111111011000011110100110100010011100010101011111011111001010110000111001100001001011010010011110010011011010000000111111001110100100000010101111001;
#1 $display("%b", po);
# 1  pi=207'b100011111111010001010111000101100100111001111101100010101010010000000001111100100111111100011100010010010010001011101110000101101110100100010001000101100000010001000000101000010111011111111010100110000011011;
#1 $display("%b", po);
# 1  pi=207'b011010101110111100100100010110110100010101110100000100100001100010101101101010110001010000011001011001100110001000011100100111011100100010001001111011001000001010101100100100100010110100011010110100011111001;
#1 $display("%b", po);
# 1  pi=207'b001100011001111101101011011000100001110101011011011001010001000110110001000101010100110110110111100000010101111101000000101110000011111001110010011000001100001100100110010001100100110011010001010010010001111;
#1 $display("%b", po);
# 1  pi=207'b000101100011110001111100001011010111010000110001010101000010100111111100110011110100010000000011101011110101111110111111011110010110010000101111101000011110101110001001100111010011010110000001110111011101100;
#1 $display("%b", po);
# 1  pi=207'b110111100000000011000111101101100001000100111000101101001000000100110011010111100011000100110011011000111001100000111011101011010001111100110100111010100101100001111100011011010001010011000101101101100101010;
#1 $display("%b", po);
# 1  pi=207'b000100000001001100101010001010110110011110101000010011001000001011010111001000111111101000010011100011001010110110110101011111100011101101110101110001001001101100010011011010011000100010101001111111011111101;
#1 $display("%b", po);
# 1  pi=207'b101111111100011110010000011110101011110011100000110010110001110101101001011011110100001101111110000110100001001010111110101101011010101101101001111100101011100111110111011001101001011101111000101101111100011;
#1 $display("%b", po);
# 1  pi=207'b111000011111010000001111110110101011110101110010010010010010101100111111111011010100010101100111001011010100010101111110111110111100011100010111100100110010011011101010111111100000110100000111001011001010001;
#1 $display("%b", po);
# 1  pi=207'b101111110111011101000010100011001111000001010000100111001110101000010011010010101101001010100101100011010100001110111001011101000100010110100000111000011010100111111110001010011010111110100000101001000110010;
#1 $display("%b", po);
# 1  pi=207'b110001011000111110100111111010001101111010010000111010010011101001011100110011100101011010110110111101110110010101001010110101100011100001000100101011001010100001110111111010110000000010100110001011100001100;
#1 $display("%b", po);
# 1  pi=207'b111101101000000110001101011001011001101110110000010111100100101001001001001101110110010110010011110011001110001100110000110010010000110101110010010001011000001101110000010100001010110110110011101000010001000;
#1 $display("%b", po);
# 1  pi=207'b000000110011001000001001011010010101101000011110011111000010000100110101110000010111101000001010000011110100000101011001000000101100010010110110000100010111000000001101010100111000000011011000010111111111010;
#1 $display("%b", po);
# 1  pi=207'b111010110111001101001111100101100000000000000011111111001011001001110011110110100110010001011000010000011110100001100011000111111010000101010101111100001000111110100000010111100101001001000110001111100011101;
#1 $display("%b", po);
# 1  pi=207'b000000111101010011101101100101001101010101001011000000100000100011101011000111000000111001101111111000001000001011000001001010111011001110011110010001011011100110011010011011000100111001001110101010001111111;
#1 $display("%b", po);
# 1  pi=207'b100010100110000000001111010000011101000100010000001011100001101110000110100101100011110100011110101100111000000010010010011011110001110111111111010001010100010101001000101111111011100001101100011100110110000;
#1 $display("%b", po);
# 1  pi=207'b001111000011010001100010000111010101100111010001000110010110011001011111000010101011000000010010011111101111001111011100110110100010111111001001101110101010111010100000011101110110011100101110110011011100101;
#1 $display("%b", po);
# 1  pi=207'b011001000100100100000101101101100100000100010111010111000001101010010110011000000001100000101011111110010111011001111011110100010111010001110111010110011100001000001100110010000111001100001111110100011010010;
#1 $display("%b", po);
# 1  pi=207'b001111100111001001000100001101110011101010000000111011000101000001001001101110110001111000000101111010100100000100011011000011101100111001011000111111101000110100100001011000111100100001010000011011111000110;
#1 $display("%b", po);
# 1  pi=207'b010000000100010111110011010110000111011100001011001000100001011101001100100001010011101011000001100011101111100110111110011001100000110100111101011101111011110011010010110010111100100100001101010001111111010;
#1 $display("%b", po);
# 1  pi=207'b000100110111101110000011010111001001001011100010010011011101001111100101010111001110010111011110000111111010111010101000000011010010111010100000011011001100011110110100111110110011000010010111100100110111110;
#1 $display("%b", po);
# 1  pi=207'b010111011110111100100011100111101000111111010001111010001010110110100110101000011010010001100000010010011100101111100100111010001100011110010100111111010010000111011011010110001000100110001111000011010111100;
#1 $display("%b", po);
# 1  pi=207'b110000101011010100000100110001011110110000111110111110011011001100000101000001011100001001110100001110111001111101101110010010000011001011101000101111101000001001110001111001100101011000010011110110001111010;
#1 $display("%b", po);
# 1  pi=207'b011111101101101010010100000101001100110100110100100000011100110001010100110110010100100010110011110011001101101001001000110011111001110101000101100001001111011010010100111001100111110011110000110100111000001;
#1 $display("%b", po);
# 1  pi=207'b111111101101111100110101110110000010010110101100101110101010101100110110100100010011111011001000011011110111010111000101111001110011010000100000100001010110101010110010110011011011111101000000100110000011000;
#1 $display("%b", po);
# 1  pi=207'b011000101010100000010110011001000110100000110001100011101101110101111111100101111110000100010111011011011011111010111111010100110010010011110111100010100100010010011111111110101000101111001000101111110111011;
#1 $display("%b", po);
# 1  pi=207'b101000100111000101001010101011111110001111010101101001011010011110010000010000110100101110110111111010010010110101110010101100110011000100010111001010110100111011101110100001001101011000111001100000001110011;
#1 $display("%b", po);
# 1  pi=207'b011000000111000101000101000001100001111011000000011110111000010000000000000001110100111011011111100010100000001010010101110010111101010001101100111101011001000000100101001101000111110010101101000001011000110;
#1 $display("%b", po);
# 1  pi=207'b100000101101000010000000100001111000111010101111101111000000110011110000010011010101001011100010010111010001010001100010000010011111010110101101000000000010001111111011110010100110110010100101101001100111110;
#1 $display("%b", po);
# 1  pi=207'b000001110101110100000111101011000111011001011111100001010000010011100100010011001000110001000101010001000000111000100100001011011010100001101001001000111110110111111010111000001111111001101110111010011111100;
#1 $display("%b", po);
# 1  pi=207'b111111110001101100110010011110010010001001010000110011010111001000000100001100110111011100000011100100001111110110010000110110010010001101101100000110111101011110010110110011101010111001001011100100110011001;
#1 $display("%b", po);
# 1  pi=207'b001010100010010101100011110001000111100001000011010000101110101011010000001110100100110001100110101110010111110001001111000101110000111010000011100111010100100000001011011111011111010110000010010100011011001;
#1 $display("%b", po);
# 1  pi=207'b111100101100000010000100110110100001101010011100100110101110000001001001011101101010000000011111100010000010000001011000011000101010010110001110001001011100111110111010100100010110011100010101110111100010010;
#1 $display("%b", po);
# 1  pi=207'b011111100001100111000000110011101001111111000011010101000000110101011010011110111101011110001001110100011010001101101001111101001101010101100001101100000100011100001011110111011111111010001011011100110111010;
#1 $display("%b", po);
# 1  pi=207'b001011010100000111011001011010011111001110111011101001001101011101111011111110001101001111000011100110100000110100010110110000010110111000101000000110101000100011001010011110100111011010001011000111001010101;
#1 $display("%b", po);
# 1  pi=207'b110100001010001011101010110011100111101011100010111100110001000010101000010100011000110010110111000100101010001011001000110000001001111010001110101110011000111000010101101000010010010011011101000100110001100;
#1 $display("%b", po);
# 1  pi=207'b011110011000100101110101100100001010101110100000010110100011100111110111111111111101000111001000111111110000100110100101010110111110011010001101000101000110100010011000000100100000100011001100001000110101111;
#1 $display("%b", po);
# 1  pi=207'b001111011001011110101110100110111110111100111101000110001110111001001101010010111000010011011111101001110100101101010110110001000000011111101101010100110011001111010010000110001011101010000000101101110011001;
#1 $display("%b", po);
# 1  pi=207'b100011110110101001100111100110101101011110111100111100100111110011101110111111111101011010110010000111100001100010110111111010111100011101111011011001101110000000101100001011111001010000111001110001001010000;
#1 $display("%b", po);
# 1  pi=207'b001110000100001100001101101011000000010110101111111110101100111101010010101010000110000110110011011100000000100000000001011110000010010011110010111011001001100100011011010001011010001111111111111101100000011;
#1 $display("%b", po);
# 1  pi=207'b100010010101001010100100100100111101110000011111110101110010001101111000101010101010100110100000001111101001101101011101011111001111011111101100000110111001100010001010000101100011011100000000101011010101010;
#1 $display("%b", po);
# 1  pi=207'b010101001110001100001101000011101011101001101010101000111011000011101011011010000100011000110010001100111101110111010000110101001111110100001001011011111011000100001101110100111010111111000010100000100101011;
#1 $display("%b", po);
# 1  pi=207'b100110101100001100100101010100000011101010001000110011101110101001010001101000100001001111001011111100001100100101010011001010101011110101101100001100001000000111100101010010001111001001100111101001010000001;
#1 $display("%b", po);
# 1  pi=207'b010010011001001011101000001110011100001100001100011011101111000101001011110010000001100001100010111011011110101100111101100011101010110111100111100111101010101000000011111000010111110000100010010101110101110;
#1 $display("%b", po);
# 1  pi=207'b100110101111111100101001101101101000001101010111111100100001100011101100111110110001001000110111010010011001000001100111110111001111101010000001100001111101000000000111100001100110111000101101100011101100100;
#1 $display("%b", po);
# 1  pi=207'b010011010001011101010001100110110101111010000001001001111010000100101010000010011011000010011100010100010101100101110101011110010101000000110000000111010011101000000101111101101110011110000001111100101101000;
#1 $display("%b", po);
# 1  pi=207'b000011010101100001111011100101001001000011001010010110111110001101010111111011001111001100010100001100101111100101000000100101111011011010010101101111001111101100000010010001001011001010110010001010101100000;
#1 $display("%b", po);
# 1  pi=207'b100001001100011011000111100010111010001101010110010100101010101100100010101010000001010010000100101111111001010001001011001111001001100100011011011110111001011000101111011000001101011011100100111000101110001;
#1 $display("%b", po);
# 1  pi=207'b101000100000000010101001011100001000000101110001010000010011010001010111110100001010110001111101111011001100101000011111110011101111011000010010101001001011110010100000101110010100011000101110010100010110000;
#1 $display("%b", po);
# 1  pi=207'b001100110011001101111110100000101011000111101100001101011001110010111011100011011100111010111100000101011101000100011100100000001110010010101100111000010110011010001011101001111000011011011111001101011100111;
#1 $display("%b", po);
# 1  pi=207'b100101110111110111111001011101110110000100100101001001011111011111111111101111110100111010110010010000001001001001100110111111010110001010011001000001110101011010100111101100000001001010111011001110101100000;
#1 $display("%b", po);
# 1  pi=207'b111101001001111011001110100101110001000011010010011101011010010000001111000001000001001110011100011110101000001110010111011000111100000000101100100100101010101101010111110111010001010110111110101111000100001;
#1 $display("%b", po);
# 1  pi=207'b101111101000001100110010100111100110110110110100010010101100111111101100010110100011111110010000110010001100001001000000011001101110001111001110001010100100101110010111001001010000000010110110001011000100111;
#1 $display("%b", po);
# 1  pi=207'b111100010111100001010001111101010101111010001101001000111000111110010010000000110000000011001101010010010101100011100001000001101100100011110111101010011110010101011101011110010110001101101100010100110110010;
#1 $display("%b", po);
# 1  pi=207'b010011010000110101001110001101100000011001000000100110000110101000100000101100100011000110001000000110000011101100001101100110100111110100010000001000011010110001000111010101101111111010100101010001011011110;
#1 $display("%b", po);
# 1  pi=207'b110111001010111011111011111011000100110011000010010110000010001010001001000011000111110011010101000111010111100101111001111010110011011100110010111001010100111001001011100010110001111000110001011110010110110;
#1 $display("%b", po);
# 1  pi=207'b101111001001001100101111010110101001011001111011001011111110011010100011100011000100001001001000111010111111110100110101001011001010101110010110010101111001010000001100101101000010111110011011011110011100111;
#1 $display("%b", po);
# 1  pi=207'b011001001100001101010111011111011011101001010101011111101101100011000110010000101101000000010010010100011010101010011110101001001110000001101000101101011101011111011010110111000011100001011100100000011110001;
#1 $display("%b", po);
# 1  pi=207'b010101011101100000100110100110101011111111000110100000101001101000000110100001000100011011110101000100000011100111000011011110001111111000000101101110010010100010011010011101100101111001101011001000000100100;
#1 $display("%b", po);
# 1  pi=207'b010001011111101110111000101110101111010011101101110110010011101101100100111001011100001011001011010011111100011110011101011101110100000001011001011001101001001111110100110010111101111010010100010011010110010;
#1 $display("%b", po);
# 1  pi=207'b100110001000010110101101000011110110010011110100110101100100110100101110011000101011011111111110010100101011110111111000000111100100100000010011100111101110100100101010101111100000001010111100010001001111100;
#1 $display("%b", po);
# 1  pi=207'b111010000011000111001001100000011000010011100010111011110011001000101001000100100111111011101101010101111000010110100110010010000111000111111010111011100101110110000101111100110011101111111001000111010001001;
#1 $display("%b", po);
# 1  pi=207'b010111001110110001101011110001101001011000101100000000110000101111101011001111101110101110011100010110011101011010100010010010000011100001110000110011011010001011001111110011101100100001010000000110110111110;
#1 $display("%b", po);
# 1  pi=207'b011101011100101110100101010110110001001110010001101011100001000110011011011111001111111111110111010010111010110101101001001001011000101111101101001010010100000010110011000101000101101011011001111001111000010;
#1 $display("%b", po);
# 1  pi=207'b000000101011110111010101011011101001100000101110010001110011000010100111010010100000110011110000111111110110111101001111110010010100011111010101010011101100001110110111000010101000000100101001001111001111000;
#1 $display("%b", po);
# 1  pi=207'b101010110100001110111110111000101111100001001011101101110110010101101101111101100001111111001001010011000101101000101011101100110110010100111101100000101000011001000000000101011111011101001111010110010010101;
#1 $display("%b", po);
# 1  pi=207'b110100101000001101001110101000000100100011101110011001010000100101100111101100001010001100110011110100010010000110011111111001010001101110010110101010111100010010111100011001100000101011100101010000010110101;
#1 $display("%b", po);
# 1  pi=207'b110110101001000100000011110110111010011000101100101010001110110000011101100111111000001001000101010011011011100110111111000011100000110000110110001111101111100011100001000011110011100010100101110100010110110;
#1 $display("%b", po);
# 1  pi=207'b110010100011011011110100000000001111001101000110110100100001111010111100101100100101010001100100010010101011100100101101010110011110111110101100010100101010000010101110001011110011011100111010111111110011011;
#1 $display("%b", po);
# 1  pi=207'b011001100111011010000100101101010110001011011111000011111001001000110001111000111100011011110101111100100110000010001100000010101010100111101011000000111101000010001110001110111110001010111010110011111100000;
#1 $display("%b", po);
# 1  pi=207'b100111000000010011111111111110010100011001011101001101010100110111001011010000011000010100000101001111000110111101110101001001100000101111100101111110101111101011001001100011000010011101111010101111000000011;
#1 $display("%b", po);
# 1  pi=207'b010101010111111111110011001011000110101100001001111001010110000110101011110001011101110010001100010011101011111101110000011001111101000001101011101011110101001011100010111000010110010101000000111111110101111;
#1 $display("%b", po);
# 1  pi=207'b101000101101001110101010010011101010001010110000111100111110111000111100110100000011001101001010011000101001001000001001111011110011010111011000001111000010011100001100011010011100110100110101001001001101000;
#1 $display("%b", po);
# 1  pi=207'b101110101010110010010111010100011100000100110010100111110010010111100110010101010001011101010010011010001010110111110110000101000011100111001110010111111110110101111101100101110100010001111010100101101101110;
#1 $display("%b", po);
# 1  pi=207'b011111011101011100000000110000011000000001011001101101001000000000011000000101001011001110101011011010100101111101100010101101110101100000100001110101010000100011010001011101100011011101010010110100110110100;
#1 $display("%b", po);
# 1  pi=207'b011101110100100111001001111011110001010110100100111000000011100001000111111001000111100111110101100111111111001111010110001110110101000011010100110000011101111101111010101000001101010110101001100110101010011;
#1 $display("%b", po);
# 1  pi=207'b010101001111000010110000111101011101000010010110011111101000101010110000000001000101010111010011011101011100101000100011110011011001011111011000001110110000101011010101000111000011101101100001100110000010110;
#1 $display("%b", po);
# 1  pi=207'b101111001110100010101000001111010000011110101110001001100000111111111010000110011001001101110000000010000110101100100011010110000101111001010010110110101101011011110100001011011001111010111011110101000011100;
#1 $display("%b", po);
# 1  pi=207'b111010001001110111011001101011110110010011110111001001101111011111100100100011011110111101101111001100000100011110011000101100101111011010100000100111001000001110000010000101000001111000100001101001011101101;
#1 $display("%b", po);
# 1  pi=207'b000010110101000100101100001101101001010001110110101110011100100111000110000101101100100111100001111111100000110010011001101101000011000000001011010011000100001000111111110101001111100010111001000000101011101;
#1 $display("%b", po);
# 1  pi=207'b000111100110100001100110001010010111010001010000010100101000011010011101010110011001010101010101110011101000010110011110110001010101010010010111010011000010111001001001100111010100000111110000010001100000111;
#1 $display("%b", po);
# 1  pi=207'b001010110001100001000010100011001011000000111111111111010111000111000110110000011111000010011011010001000000111100000010001101000011111000010001001010011110110111111010001110111100100010011101001111111101101;
#1 $display("%b", po);
# 1  pi=207'b111111000000110010111110101011101010101111010110111000100111101110101001010010011111101011000000100011000111100111100001101110000000111011001011101011101000100001101011000011100111101010111010111110011001001;
#1 $display("%b", po);
# 1  pi=207'b110001011100011111100110100001010011011101001010100010101000100001011111010000010101110000110001100011101000001111101001100010010100010000111010111100011110100111100000100100101001000111011001000010010001010;
#1 $display("%b", po);
# 1  pi=207'b101001011101001111111001010000111101000001011000101000101101100010010111101011000010110111111110101101101000110110011110001001101110100101001111011011100000001000000101110000100101110011010110010101110001001;
#1 $display("%b", po);
# 1  pi=207'b001010111011111000010001100001110001000010000100010010000110010101110001110100100100010001101110010101111001110100001001111011010000111000110111010101111010000000101100001011011110001000101001011100111100110;
#1 $display("%b", po);
# 1  pi=207'b010100000100100111010101011010011101011110010000110011001111010110010000110011111100010110100011001000110001001000101001101001101110100101110010110001011111011001101011001101100111010110100000010101011001010;
#1 $display("%b", po);
# 1  pi=207'b101111010010010010011111110100011011101011000000100001001101010111000111100010111010010001000000100101010010010000000100111100100101000110100001100011110001110111111011000101001111110011001100011011111101101;
#1 $display("%b", po);
# 1  pi=207'b100000010111000010100101011111111001010011110011111101111101101010001010000101100101100100101111100010110111000001111100111111010010111110000101001011000101011100100110101100111000011001100100001111011100111;
#1 $display("%b", po);
# 1  pi=207'b011111101100001011011100010100100011011100111110010110111001000101110011100000001011110001110000001110110000001011111100010110000010110000010011110110110100100001001101001010000000010001100111011110010010100;
#1 $display("%b", po);
# 1  pi=207'b101001000000000001110000111011100011001110101000011110101010001011100111111100111110100011001110011110011111001110001111111111101010101011011000101100110001001111011110000101011111011101111100101001100101010;
#1 $display("%b", po);
# 1  pi=207'b111101010011000100011100001110111111110110101111100101100111000111000011010101111110101101111011010100110011101101001001110011010110011010110010100100010101011001001110101111111110100110000111010000011111000;
#1 $display("%b", po);
# 1  pi=207'b101000101101111100100101000001001101010100110111101001101101001101000101011011000001001010101000010010001101110010110000110010011101101000000111000111011001111000101001010011101001100110100001011101110101100;
#1 $display("%b", po);
# 1  pi=207'b000011011111000101001100110101001101000101000101111101110000111111101010010101001010111111101110100011101110100000011111000001101101100111110010111010001000001100101110111010011011010001111110011011101101000;
#1 $display("%b", po);
# 1  pi=207'b000111111110111001010000010011011010110001111011001001000010111101010011100010110110100111010111100110001101100000011111011110000100111011100000101110110011110011000010111011110000110000000010101000100111101;
#1 $display("%b", po);
# 1  pi=207'b110100100011110111001011111011011011101001010111011111101111001101110110010111110011000010101011010000011110101110001001011010011001000110111010011000010101111111001101000111000010010001010010010100100000011;
#1 $display("%b", po);
# 1  pi=207'b011010000100111111100101000111101001101110100111110001000000011110001010010000100011110001010111000110010000100101010100111100111010110111101100000000010001111110110011101000001111001110101001110100011010101;
#1 $display("%b", po);
# 1  pi=207'b101011011111111000111110011011000110110010001001011111111000011101001111011111001001110011100000101010001011000010101011100111011010010111101001001100101010101111000111100101011011110100101111100000001101110;
#1 $display("%b", po);
# 1  pi=207'b100101011001001111000011010010010001111110100111101110110010001001100100110110101010101110010010001111100010000000101000111111101001100100101000100010010010000110111111011100100110101101100011011011010011101;
#1 $display("%b", po);
# 1  pi=207'b100001101011110000011110101000011001010001001110001011110001111110010000011001111110011010110001110110001111100001110000000000000101110011011110111111100110100110010111100110100111101001111111110101100001100;
#1 $display("%b", po);
# 1  pi=207'b101110111111001011000111100110000111100110010000010011100110011010110001111110111101011111100101001001110110111101010001100011011011100001010011110010010001000001101001110111010110101000000101000000101000101;
#1 $display("%b", po);
# 1  pi=207'b101111011001100010111101001101100100011100001000111000101100001001000100001000101010001011100010100000111011001111100001100100110000110111101100100001100000111000001101100100010001101011100000011001100010001;
#1 $display("%b", po);
# 1  pi=207'b000110000111101000001111000010000111011000010011001010101001100000001110110110111100111100110110101011111010010001011001101111011110110010100100010101100110100111111101000111010110110000111011001110000100100;
#1 $display("%b", po);
# 1  pi=207'b101111011111001000000101001111100110100110011000111001010100010100101000100100001100111101101000011011101111111011101011100110001110001111000111100000001010110010111001001010111110010001101010110111000010101;
#1 $display("%b", po);
# 1  pi=207'b110110100111101101101000001011101011110110100000110111100110010101110011100001100101001000000100000010110110001100001111110000011010001000000001011001110111010001001001000011101100110110010011001110000100001;
#1 $display("%b", po);
# 1  pi=207'b001010010100110101110101000101111010000100111110100111101100010001100100011001111010001000111011001001001101011110001101110101100111011010000101110011111000011101100110101001010100111110000101111001010110110;
#1 $display("%b", po);
# 1  pi=207'b110000110101111110011001010000100011110010011000101011000111011100000001111100101000001011011001100111110011111000110000111101000000110011001101001100011010001101011111100100010101100111010011110111010110001;
#1 $display("%b", po);
# 1  pi=207'b010100011011110001101111110000111011111100101001101100001110001010010100011010100100011011000001101011100111001010110010011101000010110001001001010010001010010001011111110101010111101011110010000001001000001;
#1 $display("%b", po);
# 1  pi=207'b000110111000101011101101001010010011111001111101010110001100110000000001100010100111001000010010001100101011000000010011101110100000011101111011110011010111001100011111100011111110110010110001000001010111000;
#1 $display("%b", po);
# 1  pi=207'b001000000111011011101101110110010110100101000100000000000011100110110010011101111001100101000011001100010100011111101010111000111100010110101100010100111000111011001111100001010101000110001111100111001001100;
#1 $display("%b", po);
# 1  pi=207'b110110011111100101000011001100111011101101000111110111111110101101101100000001110000101000011101011101100010001000110001011101100111110001111111001010111101100101111111100111011000011101001110101001101000100;
#1 $display("%b", po);
# 1  pi=207'b100011111100100110101001001001011101010011111001011001000100101100101100001011110011110000011110010000110000110010100000101110001010100101001010010111011110100000010000000100011011010001010011001101011101011;
#1 $display("%b", po);
# 1  pi=207'b001010000111101011111110011010000001110010001101001101101000010010101111011101110010000101010100111001001101111101101010000010111010110111101011011011101110101011111100101001111011100000000101000001010000101;
#1 $display("%b", po);
# 1  pi=207'b000101011000010000011001001010111001110001110001111101000110011001101110001101101000100001111110100010001000110111011010110000111000000011100001110111011000110100110110001011011101110011010111110000111110111;
#1 $display("%b", po);
# 1  pi=207'b110110101011101000011101101011000100101100000011011110111000100111110111010100111011010001111001110110000110110111001100110100100111100110110110110100100011111111000001010010001011110110001011001001010101011;
#1 $display("%b", po);
# 1  pi=207'b000111010101100011011010000001111010001001010101000110101011100110111001111110011111011001011001000010100001001000111111110110101000111101110011110101000000001010100000011001001100111000101101000000001011001;
#1 $display("%b", po);
# 1  pi=207'b110101101101010111111001001101000000010100110111011001001001100011001011110001000111110100011101011001100010000100110010111000101110011001011001111100001111110000000001001010001001101100010000011100001001010;
#1 $display("%b", po);
# 1  pi=207'b100111001111001100010000000001110110100100101111111001001111010000011101101111001111011110001111101110010000100101100110111000001111000000101010110101001011110011100111111001001111010100010100101000100000001;
#1 $display("%b", po);
# 1  pi=207'b001101110011101000100000000010010100011001000111010011110110001001000100110010001010001000100010101001011101000111011000101110010000101010101111101001101100111111101010111111101000001110111110101110010010111;
#1 $display("%b", po);
# 1  pi=207'b000110010011111101000101110100000100001010111111101000001011011110100111000010111110000100100000011110001001000100011011101101000011110110001101001101101110100101101101010011110001001101010100001101100101000;
#1 $display("%b", po);
# 1  pi=207'b110100010101011111011011111000000110010010001110111001110000000101011011001111011101111110110001010101001100001100100100101110000101011111011010111111010001111100100100011100000110110101110111110001100110010;
#1 $display("%b", po);
# 1  pi=207'b000111011110100001100100010000110001011010010101111001001000100111111001000000111110110000110001100010101111000110011110111101001010000000100011101011001100101101011000000011001110011011111101100011000101000;
#1 $display("%b", po);
# 1  pi=207'b101111011111111000110111111000110111010110001000000100010100001000100110000001101000001111101011101011111010110101001111100101000110000100111101001110011001110110110111001100000100101100101001010000110001010;
#1 $display("%b", po);
# 1  pi=207'b001000000001001101110010011101101010001111110000110111111010001010110100001011100001100111011001100110100111111101101111011001100010110110011010001100000100111111101000000101100001101100011111110001001001011;
#1 $display("%b", po);
# 1  pi=207'b111100100110111110110110101010101101001000000110100001111110110110011101010100000101011110011111010000011100011011010100110110100110110100011001100001111110100100010001101010110110010101010011111110101001111;
#1 $display("%b", po);
# 1  pi=207'b000101110011101010010110100111000000100100110000111110101111001100110101000010100110011001111011000110001010010000010100011001001010011110001100001011001011010110101001101110111000110000010101010000111101110;
#1 $display("%b", po);
# 1  pi=207'b000000001111110001111001111000100101111010010111010100000001110010111010101110011011101101101010000010011111110111100011010001111010001110010100000011000000001111100011000111100010100111011101101010111111100;
#1 $display("%b", po);
# 1  pi=207'b010100101110110110010000000101001011010110001011010000101000111110010100010001011000100010101100101101110001010010011101111010010000111011001101100011010000010001001101010010110011011110101100000101010010101;
#1 $display("%b", po);
# 1  pi=207'b011000110011101100111110001001001001111001101110011001110010110100010001110001000011100010111100100110011101010011000010111110101011000110100011101110110100101110010001101110011110101011110101000100101011000;
#1 $display("%b", po);
# 1  pi=207'b110110100001000100001011011001011110000001001011001101011011110100111001010011100111010101001001010111000011010101000101101111110111000111000010100101101001001010101101000010100110110010010110001001101110010;
#1 $display("%b", po);
# 1  pi=207'b101110101011001000100101000001110000100011001101010100110001001001111100110001100100101111110010111111001011110000111011111110111101111010101001101000111101000011011011011100000110011101000111101010111100011;
#1 $display("%b", po);
# 1  pi=207'b100110100001001001001000011101100000100110001011010101111001010110011010110011000011011111000001110110011000001110111000011010101111100101111110000001000000101000101111010000110101000111111000011011110110010;
#1 $display("%b", po);
# 1  pi=207'b111100001100101110110010110101111110110001011001001111101011001100011000011101001101100101110000001000110001111010010100111010100111001111100101111100000011010001110111011010101110011111111101100001100101010;
#1 $display("%b", po);
# 1  pi=207'b101101111101011100010111110001010011110101111100111010101111101110101011111000001000111011100111010110110101010011101110010101000010010011100010001111010011001101011010011110011111110000011100000011001011001;
#1 $display("%b", po);
# 1  pi=207'b101000010110011011100111010101001101110101010010000111111100010110011001011100011101011000111010000101110000100010110111010101110111100100100010100010110100001011111001000100011101000111101111010001111111011;
#1 $display("%b", po);
# 1  pi=207'b110000101111010111111011111010011101111000000111100011001111000111000101111000100111101000010110000010110001111101011111111101111111010111111000110011111011100011100001110110110000000010101011010101001110110;
#1 $display("%b", po);
# 1  pi=207'b100010010100000010100011011010100111111000110000000010100000000000000010101111101100111101101110001101110011111001110100001001101110001111101111111010100111111110100011010001001000010010001100001010011010000;
#1 $display("%b", po);
# 1  pi=207'b001100000010000101000100001011001011111100101100000100011010110101111100111110100111101011100000011100011001101110101000010011110110101100001111111100000000000100001100001011110100010000000011000001011010100;
#1 $display("%b", po);
# 1  pi=207'b011110100100001110001100100111111100101010011110110100000010001010100101010010110001110000110111010010111110110101011100101100001111111111000001111111000010101101111101000000100010011111110000100000000001011;
#1 $display("%b", po);
# 1  pi=207'b001010100100101111111001011011111011011001110011111010101001000010001000111001001111100100111101011010000010110101111100000100001100101001011010001000000101001010111110100110101011000000010000111011000110001;
#1 $display("%b", po);
# 1  pi=207'b111111111011010001001011001111011111001100010011010010001000100001110001000100000001001101110111110100100100100101000010100101100111101011010111001000000000000111011000001010111111100101001110110111110111101;
#1 $display("%b", po);
# 1  pi=207'b111101001010100101101001101010100100001100001111111001101000111100000011100101111010000001001001111100001101110001000110101011000110110100001100001001111010100011010100001010101110001000010011001100111011101;
#1 $display("%b", po);
# 1  pi=207'b000011010001110011010000110101110010101110000001100000100010110001100001110111010101111111110001100100011111110000000001010111101011101010101111110001000110011000011000001110001110110010110100110001000110100;
#1 $display("%b", po);
# 1  pi=207'b110011111111011110001111001100111001110010110111000101111011111101001000000111000100101101110111100011010001000110011110101001010111011010001001000111110000110010001111010110001101111100001101101100100011101;
#1 $display("%b", po);
# 1  pi=207'b001001011111010011001001101111100001010110100001101000101110110011110010100000000100011011101011010011101110100101001110000001000110111101101000000111011011110000000011100100011111110010011000001000101000001;
#1 $display("%b", po);
# 1  pi=207'b111010110000100001110110100010001101000110101101011001100000001000010111000010011010100110101100100100111110000100100000010110110011011011100001100001111001001101010110001111001101110001001010000011100010011;
#1 $display("%b", po);
# 1  pi=207'b100100100110001101011111101111110001101111001100000100001001101011110110101011000100101010101001101001101000001100111000111100010000100011010000110010001011010110110111011000110000100000110011000110010110011;
#1 $display("%b", po);
# 1  pi=207'b001010011001010010001001001001100110111110101110011011101100111101110110000010010101100100000001011100011011001010010001010100111110111001011011110001011100000101100001001111100001000011010000101110000010100;
#1 $display("%b", po);
# 1  pi=207'b101101011011110010111001100011000011011111010100111000101111011010010111110100101010000001111111110101010000101010010010110000000010011000000011111110000100100001111001110100101110010001111000110010010101100;
#1 $display("%b", po);
# 1  pi=207'b010011010101100101011110000000000011011100001001110011010001011010110001001110101011111000000111010010100100111101111101101111001111100110111100111010011001011011011010011100100010011100011110010111011110000;
#1 $display("%b", po);
# 1  pi=207'b001010110111010111110011010010100010111010101111010111000000001101111010101011100101110110100110111111000000011000010010101001100000111101101111011011110110110001101110110111111000111010111101011111010000010;
#1 $display("%b", po);
# 1  pi=207'b001100100010110011100000101000110110001011101110111101110000011001001011111101101100110111111100011001001110001100001100101101110101000010100001100111101100001010000001001110010110110001101010110010101001011;
#1 $display("%b", po);
# 1  pi=207'b101111111111000011011011010011010101011111000010000000100011011000111011111010011101110100001000110011010101010000010011111000101101010010010001011110110100001010111000111001110011111011011100010110010000011;
#1 $display("%b", po);
# 1  pi=207'b111010110110010111101101010110111111100101111111000110001100110011010100010010100111101110000010100010111000100111101111000111010010011011110110101101111011101100010110110101000110011010010100111001001111000;
#1 $display("%b", po);
# 1  pi=207'b101000000011101111010110111101001110010000101101001101011000001101000001110011011010000111111101101001011100100000100011000111101101110001111100111100010100001010010010011010001100110110000100111000000101110;
#1 $display("%b", po);
# 1  pi=207'b011110001111100111110010001101011001110100001010011010000010110111000111111000001100000000011110101110110101010110110100011111101101000010111110100001011101111100100011110111001011100010001110111101110000010;
#1 $display("%b", po);
# 1  pi=207'b101111010000011010011111100101001111101011110001011001111011110011000001010010001101000100110110101000010011001100110000100111011011101011001001111111011011100100010111111001100110100000111011000100011001111;
#1 $display("%b", po);
# 1  pi=207'b100111011101000110101010100100010100011011001101100001100100101010111010111011101100011110001111101000000011001111011001110101001001110011111010111001110100011101001011111000101011110001100000101101000001110;
#1 $display("%b", po);
# 1  pi=207'b001010010110101100100001010000011100110011101111110110100011001010100101101100000101100100100011100101010111011000011111110000001100001001101110110100111111011101101101110100000101111110100000011001110001101;
#1 $display("%b", po);
# 1  pi=207'b001001101101000111100010010111111000111011100100001000010000111100011100101001010100101111100101010010110000001100100110110101101011100011101110011101001101010010111010101100101111100101100110010000011001100;
#1 $display("%b", po);
# 1  pi=207'b101101001010001111010110111001011101010001010110010110100010011110010110111000010111011001111001100011000110101011011001010000000011111100011010100101101010111000000011110010110110001010010101110110010010111;
#1 $display("%b", po);
# 1  pi=207'b001111001111110000111000110000011000101000011010111010011011110110000110111111001010000110100000101011010110001110101000010010011001010010011101000100101110010001010011111010001100010110010011110110000001110;
#1 $display("%b", po);
# 1  pi=207'b010100100100101100001001101110101100100100010111111000101001010100110001011011001010000011101111000101100001010000011100010110010011101110100011000111011011111010010101011100001010111001001111110010110001000;
#1 $display("%b", po);
# 1  pi=207'b110100001101010001010110010011000010100010001101100001100010010111001010110001101100011010111110011111110100111101010011001110100100000100001001111100011011101101111101110101000111000100111110001001010100100;
#1 $display("%b", po);
# 1  pi=207'b110000111100010111101011011100100101101111001011100100001010110000111111111000111111101101101110101010101111011110001011111011010000010000001010110111000000010110100000010110101001101111111000011011100011011;
#1 $display("%b", po);
# 1  pi=207'b110101010101110000000010101001101100110001001011111000100110010100010010111010101110101011110100100000001110001111011100111101111110100001101110100111110100110000010010111111111011100110001110010010010110111;
#1 $display("%b", po);
# 1  pi=207'b010011100011000001101100001010010101011000100011010000011111111010011100010001010011101000110011011001010111000110000010100001101111101110001100001100101010110000110001001110000110010110000010011101100101100;
#1 $display("%b", po);
# 1  pi=207'b110100100101011110001010101011011100111110001001000001000010101011010000101010000011100100000000001100000110111011100100001001110011000101100111010010001100101111011100011010100001010110101001011101011000011;
#1 $display("%b", po);
# 1  pi=207'b101010111111011001111111100001101000001011100110101011011011010001000111000000110001100110111001001101110000100110101001011110010111111111001001000111111001110011110001001011001000001111110000111000000001001;
#1 $display("%b", po);
# 1  pi=207'b111111100111010001110111001110111010111101111011000000100011001010100100101101011010011010011111000000010001110101001111110110111101111010000100110011001101001101101001011100000010011001110100010101010111100;
#1 $display("%b", po);
# 1  pi=207'b101101010000110110010000011101001000000100001100010010001001111101111111010000100000111001111110100001101000110111011111111110011000010110011111011011111111110100101110111001111010110000001011100111000101110;
#1 $display("%b", po);
# 1  pi=207'b111111001111100010111110010101100111000010101110101100001001111010010110011010111011110010001011001111001110011011000110000101111110111001100010010101010110011110001100010111101101001110010100000000010110000;
#1 $display("%b", po);
# 1  pi=207'b010101001110011110100011011010010010000010100111101100011000001110001011000100111010111111011110101101111010010010001000011100011110101101100111100010000110111110011111100000100111110110010000011010001100011;
#1 $display("%b", po);
# 1  pi=207'b110111011011100111111111000110010010101000000010001010111001010101110000110100010110011010011010010000111000001100011010100100100001001011101110110010111111100010010100000101100011100010101101101111010110010;
#1 $display("%b", po);
# 1  pi=207'b010101001000011100001011011101101110011010001000111111110110100001011010001011011100000001110101110111000100111111110110001000000010001001111001101000101101000101100000111011100101000101110001101110010001010;
#1 $display("%b", po);
# 1  pi=207'b010000011010111100011010010010110010111111000111001001111011010000111110110101100000001001000100010100001001010100010000110110101101101001010011011000000101010110111000010111010001101101001111011000000101111;
#1 $display("%b", po);
# 1  pi=207'b010111111110011001010001111110100010110100111001111100001100111100111010101111011110111100010101110010001111011011000111010100100110000000100110111011111010011110111110101011001000101001001010111011000110110;
#1 $display("%b", po);
# 1  pi=207'b001000011010101110100010100010011011100001110100011011101110110011101100001100010101010010101011100011010101110011101010110011011110011000110000000001011111100111010001011110011010011110011101100100001011001;
#1 $display("%b", po);
# 1  pi=207'b011100011000110101010101111010110100001110110010111101100100001101101100101111101011110101111011000000000011010111011100110010100000011011110101101100011011101000011100001110101011101010011111100000010110101;
#1 $display("%b", po);
# 1  pi=207'b100100111110101001100001111010111100011010100110010011000001101010111000110100111000100101001101001111110010001001001000111110001011010011000111111011000011001110110010000010100101111000010101001001010001100;
#1 $display("%b", po);
# 1  pi=207'b000101100000010110001011001001000100111101010100000011111001011110011000001101010010111101110111111000011011000010001111100100100101001100010010000111010000011110010101001010100011111010101100011100000011011;
#1 $display("%b", po);
# 1  pi=207'b100101110100001000100001011001111010100010010101100111101111011001001111011000010100110000000111011001011101111011100101110010000010000000000000010100011101111010000001011110011011001000010000010111111000111;
#1 $display("%b", po);
# 1  pi=207'b000000110110100110111011111001100011100100110111011111110100100101101101001100001010000011010110000001000110001010011001011100001101001000011111011111111001111101000110010100100100101101011000111010110101100;
#1 $display("%b", po);
# 1  pi=207'b001000011111111110000011111000011000011010011000111011011110011000000010001100101010011101000110010001100100000111110101100000001110001110001111111011110010111001100100101000110101010010110100100100001111111;
#1 $display("%b", po);
# 1  pi=207'b010010100010000000111001101010111010011010110111100000010001011111001101000000010110010000111101110101100100000110100010110010101001100011000010000001101100011000110000010101110001111001011110001111100001111;
#1 $display("%b", po);
# 1  pi=207'b101001100101110100010110101001011011110010110011011011101000010000101100111011011011011010101000010010100111000110110011001011101010100111011100100010111000110100011001000101001101010010000111100000100100111;
#1 $display("%b", po);
# 1  pi=207'b010101001111100101010010010100111011011110010000100110110001111000010110000101010100010010101100110100110100100111111011100000100100111100001101111100100001010100111101011111010110101001011000001101001001011;
#1 $display("%b", po);
# 1  pi=207'b111000111011110011101001110000000101000101001100001010100011001111100110110000001100111001000101101111101001001011100110111011000100001011110010000000101010001011101101011100001011011000000100111110010000100;
#1 $display("%b", po);
# 1  pi=207'b100100100111000100111101110101110100110011101110110101100001000100111100001101111111000000010000110101010111110010100101010010111111001101100010010001110100000100001010011101101101110100011111000001101100110;
#1 $display("%b", po);
# 1  pi=207'b110110110111111010111111001100001001111000101100000111001010100001110110110001010000101010010010111101110111010000011001111001011101101110111111100100101111000010101100100101101000000010110110010001000111010;
#1 $display("%b", po);
# 1  pi=207'b001001110111110101110000110100110011001001000110011101011100111111010011100000011011010100010111010001111100011011000010011101101110111001010111000101101010100001010001101011000001100010111101100011100100011;
#1 $display("%b", po);
# 1  pi=207'b001110010100111010011011110001010010010000001001001000101011011100100011110100101010001010110111011111110010001110100101010010111000000110100100011111010100010010100110001100010000011001111011011101000110100;
#1 $display("%b", po);
# 1  pi=207'b000101100110101110101001111101010010001100111011010011011001000110110011100100110110010010001000011000101001111111010111100000000101110101010001101000011111110100011110000110110010111111010010000101101111000;
#1 $display("%b", po);
# 1  pi=207'b010111110111001010010011110010011101101011100101111100000011101001110001000110010100011101100100001111011110110010010011010010100100100100100111111000101110101001000010010010011001110111001100111011010101011;
#1 $display("%b", po);
# 1  pi=207'b010111011110101100111001000010010001111110110000001011010101110110011010101001011100010100011111011011011010001011001111011101101011101000101100000010111101100110101010100011111111101110001001001110010001011;
#1 $display("%b", po);
# 1  pi=207'b000101100000100111000111100110101000111101101011111010101101100101000000011011010101010010111110101101001111100110010000011000001100100001011000000111010011100011010011100001110110010101000111000000001000111;
#1 $display("%b", po);
# 1  pi=207'b101011101111010001101011000100100001011100110001101100011111110000100100011011110100000010111110011100001101100000101111001100010011001000111010000111101011111110001110001000100101000010100000101010111101000;
#1 $display("%b", po);
# 1  pi=207'b011101000111111110010010100000111000110100000111111111101101010100001010011000100001110010110111010000010111001011001111101010001001111001001001011010000001101011101000110010111101000101101101000111010001101;
#1 $display("%b", po);
# 1  pi=207'b010100001000101101001111101000011010011001110100100010010111101111111010010011011111011110110010111100111010011100001101111100100001101100011110010000111100110100000101100000100100111001000111110010011010011;
#1 $display("%b", po);
# 1  pi=207'b100010001100001101111011111111100010110100100011011000000101001000010001110100110000001101010011111101111110100001100010000000000101001110001001110111011111100111100001000000100100000011101001000110011010110;
#1 $display("%b", po);
# 1  pi=207'b001011101101010100001111001111111011100101001100011101000100100101010011110000011011011010000100001001000100100011010000011111001110011010011011101000010111100010110000011010010011001001111101110110011101011;
#1 $display("%b", po);
# 1  pi=207'b100100110001100000111001111111010011110101100101010010001011110011010011100000100100000011100000111001101001111101110100101111011111011100110100111100000001111110111111111001000100010001001110111110001010010;
#1 $display("%b", po);
# 1  pi=207'b100000110001001001100100101000110011010101001100100000101101011010000110111111011101110011110110011101000111000001111110100111010011010111111111101000110110000100001100100011101100110000100000001010101010100;
#1 $display("%b", po);
# 1  pi=207'b111100101101010100001101010011000111001110000101001100100000000101100011110010100100110011101010000101101111000001111111001111101010000010100000100001010001111000101110010010001001010110011100010001110111111;
#1 $display("%b", po);
# 1  pi=207'b010110111111111001101000001111000001001100011100101110101011010111100111011110111011001111101000000110001100011000111011011110011000101100110010000011000000011011000101110001000101111100110110100101111111100;
#1 $display("%b", po);
# 1  pi=207'b101100000101110111111001001111111110100011010101100100011110010010111000000110100010000001110111000100010011100101011100011111101111110011100001100111001110101000111000100100011110110101010001100100000011110;
#1 $display("%b", po);
# 1  pi=207'b010011101101010101111111000111001101010001111100100001101011110011100010000110010010010111010011000100100101101111100101010000101011010100100110101110011111111100000001101100010011001110101001101101111000100;
#1 $display("%b", po);
# 1  pi=207'b101011010001101010000100101011111101011000111100100100000000001010010010011111010000110010111010101011000001100101111011110110011001001110100100000110000101010000111010011101010000110010000110010100011011001;
#1 $display("%b", po);
# 1  pi=207'b001011110011110110000110001111110111000001111101001100011110110101001111000011000111110000100010111011110100010110100000001001111001100000001101101100001010110101010010001100100001010000010101101111110110000;
#1 $display("%b", po);
# 1  pi=207'b111110100100011010100011011001111110111001100010000100111000001111011011000010101000110110000110000001011011101100000111010100000101000101101101011110000110000000010110000010010011011010111001010001100001100;
#1 $display("%b", po);
# 1  pi=207'b001100000101011000011111011111011101101000111000110010110011101010100100100010000001000100001010001100000011110110001100011101100001110110111010111011101000001011001001011000110010100111110011111111100110110;
#1 $display("%b", po);
# 1  pi=207'b111001111100011111111001000000010001110000100101100001111110110001110011001011101000000000001001001001000001110111011111100001101001111101010101101011100001000000110110101011110000110010101110010110111100110;
#1 $display("%b", po);
# 1  pi=207'b001100011100100010111000100001010000111000111010110101011011111010010010011011100100111111010000011011001000001000101001111000101001100111100111001010000111111001011001100011110011011000100011100101011101001;
#1 $display("%b", po);
# 1  pi=207'b010111110011101101000011100101101000011110000100110011101111000110110101100001110001110001000010101001010110001000100010110111000000000110001101100101111101111001111101000111010101100110100111111011000000101;
#1 $display("%b", po);
# 1  pi=207'b111010011001011001001100010101011101000010011110110001110001000110001001010010101110100101110001001101010101100001011110101110101111011110011101001110010101111001111111110111111000011011011000101110111111010;
#1 $display("%b", po);
# 1  pi=207'b001001110111000101100010010011110110011110101110000100000100101111010010001010110111011101100010101001001111000101101011000110100001010011110010000010111010111001111010001111110110001110101011000010110111111;
#1 $display("%b", po);
# 1  pi=207'b001010111010010011001101110110010101001011000011101001100111110001101100101001001010110001000100011101110111110011010101000011101000100000110010101001110100010110101010000000001111110111000010100011101100001;
#1 $display("%b", po);
# 1  pi=207'b011001010010010110010110010100101001011110110111101111001100010011100000110000101010110111101011000000001000110011011011100001011101110011011111101101010000100001101111010100001001010111101100011101101001110;
#1 $display("%b", po);
# 1  pi=207'b101001011001000010011110110011011000011010111110000110011101111110001100100110110001010100001000101011010010101011000111110101010000100101011101101010111111101111100010110010011001110011100111111011100110010;
#1 $display("%b", po);
# 1  pi=207'b010000110011011010110110001000111100000011100111101100000010110101000100101010110011101111001010110011011101100000100000000111111000001100011011000010111111001000001010000010001111011101000110101011011110001;
#1 $display("%b", po);
# 1  pi=207'b101101101011101010110010101100000110101010011001011101110011010100011111101110000101011100011100010111001000111110010111000111111000000101100010111011011001011011000101000100001100100000001000000101111001110;
#1 $display("%b", po);
# 1  pi=207'b101100010111010111110101101110100001101110110001111010111110110011000011100110111000011100011101111110111101010010011000001110001101100010010101000110000010101111001000000111111100010010011101101000101110011;
#1 $display("%b", po);
# 1  pi=207'b101001000110101001011110000001000000011011000010000001100010111110111100001110000001001010000111110010010101101100010001011001110101010111101100100101111100011000010000000110000001001111101010000101011111000;
#1 $display("%b", po);
# 1  pi=207'b010000001111100100110001100100001010101110001111111000101110011010010000111001001100110011010000100011011110110101101010000101001111011111011000001010111001101111111010011000011000001010010010011011101010110;
#1 $display("%b", po);
# 1  pi=207'b100111001000100110010010001101101000110101100110111111010010101011101100100010010101001110100100011101010100101011110001001001100000001011101111010111011001110111101000101111100001000001010101101010111010011;
#1 $display("%b", po);
# 1  pi=207'b111110110100000011100010111101101111011001101111011110010011110000011101010101110110011100011010001100010100010111011111100111110111001100011000101110000000101100111100110100001101100010111110111001100100111;
#1 $display("%b", po);
# 1  pi=207'b110111100111111001000110110110001110100100011010000011001110101101111010011100100010000011111101011011011001100011000110010010110101000110001000010011110011011101101010010001110110011000011110001111100101011;
#1 $display("%b", po);
# 1  pi=207'b101011101010111100011010101011001110100011100100001001011011001101011100000001001001000001010110111000001010110111000100010001000000111011010000001011000111010000101011110100001010001001111010000001001111111;
#1 $display("%b", po);
# 1  pi=207'b100010111001001111000011001101011101000110110001101110001101000101101010000000110000111100011111010110010000101110000110110110100111001001100011111001111011000110010000100011100110110100001001011010111001110;
#1 $display("%b", po);
# 1  pi=207'b100101111110100111101000011010010111100111110001001111011000100110101011010111100000101111010010100110000011001011100001101100000011000001100110011001110010000110111001010111000101001010000000010111111110000;
#1 $display("%b", po);
# 1  pi=207'b001110101111011010000000000110011001000010110001000001010011001010000001111101111100111001110101010000011111110000000110001000110111100100101101101110011110001101100110101011011011010101000110011011101011011;
#1 $display("%b", po);
# 1  pi=207'b011101111000010000000101111111100010011111111000101011011010011010111000110111100101110100101101011010111011100101101101111001100000111110010011000011010110010111010111110000011001011001001011101001100011101;
#1 $display("%b", po);
# 1  pi=207'b000110101010111001001000010100001110001000001101011001110001001001000110100111101110111110010110011010110110011010001000110010111000100101010011001101011000001000100101100110010000011100110100110010101011110;
#1 $display("%b", po);
# 1  pi=207'b010101001001001010011001100101001100111010111100101010011111001000100011010000010000100001110110110011011111100101011110010100110001100100110000101110000011000001011000101011100101110110001100011110110100110;
#1 $display("%b", po);
# 1  pi=207'b111111110100111101100000100100100100000101101000110111101110000011010000001000000101101111101001000100001001011001111001111001110101001111001011011000011101111101101101101111000111111011000100011011111101001;
#1 $display("%b", po);
# 1  pi=207'b100100001010001010110101100100010101101111100100101011010101010000100001010100001011110100001111010110100001011010001101111010011101111110010101001010010000010011101111000001001001011000110110111111010000100;
#1 $display("%b", po);
# 1  pi=207'b101010111100110000010101101101000110101111110011000101101111000110001010101111001011100010111101111001111010000001001100001001010000011011101101101000111000100000110001111011010001110101000000010111101011100;
#1 $display("%b", po);
# 1  pi=207'b110000000011001011010110100011111110110011101101010100000010010011000010001010101111111010011001100111010110110111101101110010101111101100010001100100111100101000100101001110110110111101110010101000001011010;
#1 $display("%b", po);
# 1  pi=207'b010100010010011010001011010100110101101111010100001001111010101011100001110000101011001111100111101000010111110001001000000111110101110011101110101000100000111111010110101000100111111001010100110001110010000;
#1 $display("%b", po);
# 1  pi=207'b110010000001101000011000101101110001000000010110010000000000001101100000011011011110011010100001011001101000110000101001100111100100110110010110100100111101111011100101010000001010110101100000111101011011011;
#1 $display("%b", po);
# 1  pi=207'b111100110101110010110001010010010100010010010101100000111101110110111001001000010010110101100111001010101101101101011010110111101111010100010111110010010011011101111001001110001010010001101010010001000100111;
#1 $display("%b", po);
# 1  pi=207'b011010001010100101000000011001010100011001011010001110101011000101000010011001011101011101111100000000110101110100011000110101110010111101110001111010001110010111001011011010000001001011101100101011100101101;
#1 $display("%b", po);
# 1  pi=207'b101010111010011111101111101010001001111101010100101010011101111001101111000000101001110010001010010101101011000001001000111010100011000100111111000100110011111010001011100000011001111001001011110101110101000;
#1 $display("%b", po);
# 1  pi=207'b111010010000111110000101010001101001101111110100001111001101010011010110111110110001110111010000011110101000001011100011010111110001000001011100011000011111110000010100001110100001011010110000011010110101011;
#1 $display("%b", po);
# 1  pi=207'b000011110000010101001100010110101110100001001100111000111110101100000010010010111110100111101101011000101110010011001000110111001010100010011110100111110100011001101110100101111110101001110010101001010110100;
#1 $display("%b", po);
# 1  pi=207'b001011111000011100110111010000001001000010101100110001111101100111101001111101011001110000101110101001011100100010001000010111011101111000110000100011010010100011010101101101010101100000110111011010110011100;
#1 $display("%b", po);
# 1  pi=207'b010000011010000100101011000111110110011010111001100101111011001010111011010101100010001010100001111111000000000000110000110100010010111011100010111001010011001000010111111110100100100001111010001001101011001;
#1 $display("%b", po);
# 1  pi=207'b101001011011000010001000011001010101001100011001001111000111000000101101100011110111111101100101010111110110101000001011100111110001110101000011100101110110111111111010111001100100101110111110010001011111011;
#1 $display("%b", po);
# 1  pi=207'b000001101010000001011111011011110101001101101110101001100111100000110011011011110111000000011100110011101110001100100011100000000110001010101111000001010001010000011101101111111011000111001110100101100100100;
#1 $display("%b", po);
# 1  pi=207'b100111101001111001011100001100100100010110110011110100000000101111100000101100011011000001001100110001110100101001101000101100100110000001111011000110111101010010001100100100010111110011110001001001000111111;
#1 $display("%b", po);
# 1  pi=207'b010011011100100100001110110110111011100011001000100100100001001110111001010010111011010111110000000000100110101001101011111000101000111100001001001101111111011111111100100100011000001110011110110001000100001;
#1 $display("%b", po);
# 1  pi=207'b100000010000110001010010101111110000010110001001110100101100010001011101110100111000001011110100011001100010110000010010101011000101000010001110100110000000011111001001110101000100011101011100010010100111110;
#1 $display("%b", po);
# 1  pi=207'b000000110110111011001010111011111001010111010000000001010111010100000110111111000101011010011011010010110110011110011100111010111101110010011011110011111110011110010100101101010111100010011011111110001011001;
#1 $display("%b", po);
# 1  pi=207'b000100110011111010101010011000000011010011100001001110011111101101100000011010111100000110010010001011000101110000110011101101001001010010010101110011010110010011110111001011011111001101011010101101001111110;
#1 $display("%b", po);
# 1  pi=207'b000001100000011111000000010001101010100010000011100001010110001000111100110011100101010101100000010000111100111011001111101111001111111101011101101011010110111100100100001001000110110101000000011011110011100;
#1 $display("%b", po);
# 1  pi=207'b101101101101110101101101011110000001110100010100011000010001010001011101001010111011011101111001101001010101010011000011110010111001110111100101001010100110001001111101101110010010110100000110110010011000101;
#1 $display("%b", po);
# 1  pi=207'b111011010111101001001001010000000101000010101111000011111110010101000101100010111110111000111001001100101000000011001101110110011111101111010000000100010100001101010110000110000111000000010011100111011001111;
#1 $display("%b", po);
# 1  pi=207'b000101011100010011110000100011010100110100001011000100001101001000100000011110100110010010001011010001000111001010001101011001101001011100110010101001010110001001110010110010001010111010100101111100101011010;
#1 $display("%b", po);
# 1  pi=207'b011111111101100111111101011010000100010111000011111001010001111101110110001000100011110110000001111101100000011010101100110100011000100000001001111010100110010001001010011100010111111110100100010110011010011;
#1 $display("%b", po);
# 1  pi=207'b100100110011000110100000110011111001011000111101101101111111111101011111010101001011100100010111001111110011111111000011110111110000101000110001110011100101010110100101111100101110111001100110000101100111011;
#1 $display("%b", po);
# 1  pi=207'b010111100010110100101101010101101111000010001101100000100111011100110101001000011101000100100110101000011111001000000001111000010011110101110110001110111000110101011000011010010010001100000111011010001000001;
#1 $display("%b", po);
# 1  pi=207'b101010110111001000010101100100000000101110100100111100100110110100000010001101011000000011110111010000101010000101101110011111000011011011110010011000111110110010111110010111000011101011110101111011010000010;
#1 $display("%b", po);
# 1  pi=207'b110011011100111011011011010100011001000001101011100000110100000110001111100010011111001000100001011000011011000010111110001111011110101100100010101111011001011001101101011111111111110111100011001000010110001;
#1 $display("%b", po);
# 1  pi=207'b111100110000010010100010001001111111110110001100101101001111010000110000001001100000100000010001110111000011001000101110010001011111110100000100110011000110000010100101111011111111011010101110011101000100001;
#1 $display("%b", po);
# 1  pi=207'b000100101000100110010000111011000100001111110100100110111111011010000101111001111001010110111000101000010110100110010101000111111110110111101100100110101110010011110111110100010110111110010000001111001101000;
#1 $display("%b", po);
# 1  pi=207'b011001000000001100111110101100111010111011101000010110011110100000010101010101011111000011100011110100101011000000001010010000101100010100001001111011000111011010100111110111111101000010100111110010101011100;
#1 $display("%b", po);
# 1  pi=207'b010111100011111110000011111111101001010011101001011111011111110110000011100100110010101000100111111011000111011000001111000101011010000011010001011101011111110110100010000001001101111111000001101001110010011;
#1 $display("%b", po);
# 1  pi=207'b111000000100011101111000111100110010011001011111110011001110101011101010111000000101101100110011000010000010100100001001111000000110010010011000100001001011111100110000111111101000110101101110010010100001111;
#1 $display("%b", po);
# 1  pi=207'b101000100011100101001100000101111101100001001011100011110101000110111101111011111011100001001000011110101101101100100100111111111001000100001011010111010010111101111110111011000110111110100001110101100001001;
#1 $display("%b", po);
# 1  pi=207'b000011100001011111111001110011011010111011111000111111100001110000110000111101011111100000110101111001011101101100110010101011010110110100011100010101110011000101010001010011010111000111000110011111101101001;
#1 $display("%b", po);
# 1  pi=207'b101100001111001110011000101100011011001011010100011101010101000101000010011110011100011010010010000100111011101000110111000101100100011111101110000010110011100000101001000110011010011100100111110101110001111;
#1 $display("%b", po);
# 1  pi=207'b111101110000100010110000101000111110101110000111011010101101100000110000011001011100010110110010111000000011001010000100001100111001010010001111101010010010101110101001101000010100110010011100011011100101010;
#1 $display("%b", po);
# 1  pi=207'b100010000010111110101001000100000101011000011100001010000110001011101001000010001101100010110011001001100110101111111110100110001010110011011011001010010010011010111000011111000111010101101100011010111010100;
#1 $display("%b", po);
# 1  pi=207'b011011100110111000111111101111010101101001000000101001000011001111000010101000111010011010000000110010110000111100011100000010111011110111010101101111000111101100010010111111101011110010100110101001001111001;
#1 $display("%b", po);
# 1  pi=207'b101010110001001010011110110101011110111010001001011110010101010101101000010000111000000001011001011111011101110001001111110111111111000000001110000000001110011011000000110111011000001001101110010100111100111;
#1 $display("%b", po);
# 1  pi=207'b100110110001111100100110110101010100000101100110011001100011001110001101011001101011100101011010011110101110011100100101111010010111011111001110010100111110111101100010011000111101000000110010111010110111010;
#1 $display("%b", po);
# 1  pi=207'b011110110101111001001000111101100111110111110010000011101110011010000010100100110100001101111100100000001110111011011011111001010111110100110101110100100100101111110001101100010110110101011011101000010010001;
#1 $display("%b", po);
# 1  pi=207'b010010111001011001010011110110000111010011111101000100100111011000101100101000100101011001001010011111100010101011111011111110100000001001011111101000000011111010000101111110010100110111100110110101100100000;
#1 $display("%b", po);
# 1  pi=207'b011011100111001101101100100101011010000000010010111110010011000111110101110001100011010011010011001101100101010011110111011110110111111111010110101011011110011010100000000110111011111001000111011001011001101;
#1 $display("%b", po);
# 1  pi=207'b011000111010110111000111111011001111010100101101011100011110011001001100000010000000110101101101011001010101000110001100010110000110111001001100110001001001111100011101111001010111110001011010101010101000110;
#1 $display("%b", po);
# 1  pi=207'b011010110101110010011100011010001001110000110101100010101001111110101001001100100001111110110001010010110000100101001100100000000101110110000100110000110011110101100011110011011011111011100000110010111111110;
#1 $display("%b", po);
# 1  pi=207'b101000011000100110001111011110001111100001001111100101010100010000111111000111110101011110011110100010110101110100011101100011010110011010010101011100001100001000010110011111101011100111000001010111000110111;
#1 $display("%b", po);
# 1  pi=207'b100101110000001110000100110100110010110010100000010101110010101011010110111100011010011001000010110010001100000110010100111000001000000110111110100001101111001010110001110111111000110010111101001000110110001;
#1 $display("%b", po);
# 1  pi=207'b001010000011000100001101000100110011010111101011101101100001111111010001100000110110111101011001011110110101100011001101011010111000101001011111111010000100000100101010101111011110001100101001010111111010001;
#1 $display("%b", po);
# 1  pi=207'b101100100110111011010111011110111111111000101111111000001110001010001011011001011001001101001101110110110000101010000110110100111110100011100011100110111010101101111111011010000110010010101101100010110101011;
#1 $display("%b", po);
# 1  pi=207'b111110110111110100001111111000001001011101010111101101101100010100110101110010001111010000101011001001000001101001011010001101101110010101111101111101000111010100111100110111010001101001011001110110100101010;
#1 $display("%b", po);
# 1  pi=207'b100011000101001010001011111011001101001010111000001110000010011011001011100000011011110111011100110100011110101111111011101001000111110011001110110010101001111111011011001011000101100000011011101110001110101;
#1 $display("%b", po);
# 1  pi=207'b100010001101101001110011101000001000000010000101011010110101110011011111000110000101011111001110100101111001010110111101110001110001100011111111001110010111010010011111101100101100010000101001011011100011110;
#1 $display("%b", po);
# 1  pi=207'b100011001011111101010000101000110011000111010111001111110011110101101100010111011000101000100011001100100000100001000101010100010011011111000010010011011000111001011110100011110100010001010010100111001001111;
#1 $display("%b", po);
# 1  pi=207'b110101110001100010111111101000011010100110100111111011110001001000001011011111011101000010101000111000111111000001100101111011000111000001011100100101010100111011101101110001010010101010110110001001010101011;
#1 $display("%b", po);
# 1  pi=207'b101111000100100110010101010101111110010101000111000111110001000111101111110100110100001111000111101101111001001011100010101000111001111100100100011010111001011011010101011110001111110001101111111110000001011;
#1 $display("%b", po);
# 1  pi=207'b001000111011111110011001010100111010111101000000111111101000001111011101101100110001110101011000011101011001000110001110111110001101101111000111111011111001010110110110101001000000110011010110100101101100101;
#1 $display("%b", po);
# 1  pi=207'b110100000001010110100101111111010111111111111110010110111111011110101110010000100111011111100110111100010010001110000010000000101011011110011001001001101101100111101010001011111000101010110101111011010100001;
#1 $display("%b", po);
# 1  pi=207'b100100011101110000000110001000111110001010000111000110110001001000110100110010000001000010000011100001110001110100101110111110001010111001101011000100110101001110000000111011101011011000110110000100000100100;
#1 $display("%b", po);
# 1  pi=207'b111100010111101011001110110101011010001100011101111111100111001110001011101011100000010110100001010110110111111111110101000100011010000000110000011001100100010000011010101111011011010111001100101100101000110;
#1 $display("%b", po);
# 1  pi=207'b010110001100011110110110011000000111100100001100100011000001110101011111111001100001010010001110001101010011111010101100010111001100001011001010110111111101000111000100000100001000000000001110010011000110100;
#1 $display("%b", po);
# 1  pi=207'b100100000000011001101111010111010111001011010111111010001011001010110000110001000111100000100101100101100100000010000000001100000011001010011100100110000000111001110100011111100000111000011001110100101101100;
#1 $display("%b", po);
# 1  pi=207'b111111100000100011100111001100110100011000011100001001100000000010100000101000100000001011100100010010101001011101010011001011101011011111111101011111011101001001100001000001001110100011101010101000101111111;
#1 $display("%b", po);
# 1  pi=207'b101001011011011010111000011011001000001111101100110100001010100110111000110100101011001001101011000110010000000100101011110010101110110011010101011111101011110101100011110001111100100001000111001111111010000;
#1 $display("%b", po);
# 1  pi=207'b001010011101000010100010011001011101100010010110101100000001000110110111110101001101111001000011110001010001011100010110000000001000111001111111000100001100110101101001000101100110111001100010110001001001101;
#1 $display("%b", po);
# 1  pi=207'b000000101100100000111011100011111011010001110100011011110000111101011111100000000001111110100100001010110000010011111100010000000001111011110010111101111010111011111101010001110010000101101111011111010001001;
#1 $display("%b", po);
# 1  pi=207'b000111100011001010101010011111011110001000111111001011100101010000000110111101101110100000111010011001110100000001000001110110000101001111100111000101001110100110010100010011001100100001000011100110000001000;
#1 $display("%b", po);
# 1  pi=207'b010101010010100110011111100010000011110000110101110101010110000110011010000101011101000110011001011111110010000100010010111000110001010000111101100011110000011001101110100111110001010111101001011111101011011;
#1 $display("%b", po);
# 1  pi=207'b100001001110110011110110101010011111011000010010110001011000001100101011110100000000001101010011101000101111110110111000001101110010110101001001011110000001000000001100010010011110011100001001001010111110011;
#1 $display("%b", po);
# 1  pi=207'b111101110101001000001111010001011111101100101011011010110000001111101110100010111111011111001010000001110100111011111011101001010100100110000101001001110100000110100010110111001011010110100001101010110001000;
#1 $display("%b", po);
# 1  pi=207'b101111010001111000011011001100011101000100000111100010011001001011010000010001000111110001000000010110111010101010000000110001111000000011000001010101011101110110000001011011000111111000110011001100111111000;
#1 $display("%b", po);
# 1  pi=207'b101001001110111111010000110100100001100011100001001101010001111001001000011111001000100100000101110110010110111110000111011111010111000011001110111111101001001111110000000011011110110100011010001011100101110;
#1 $display("%b", po);
# 1  pi=207'b100100010110110001001010011100001110001100000011000010110000001001111111000100000110000101001000101000010000101011111100111001001001000010001110001110000100010000111110001010101000001010011101110000100001110;
#1 $display("%b", po);
# 1  pi=207'b111001110101001101011111001001101110100010110111000110011001100110011010101100001111000111111011100110110000000111010001100000100101011010101000101011010110110001001000111011010110001010110000000000011010000;
#1 $display("%b", po);
# 1  pi=207'b100101100001000000100101011000100111000110110110101001111000001010000101010011010100011101111011010000000110011101011101011100100001101001100000001000011100000011010111110001001010001100101100010010101001111;
#1 $display("%b", po);
# 1  pi=207'b100000011000101100001110010100010100111111101010011100010101111001000100110101100010110101001010000100100001000010011111000100000100111000000101101010101101001110011101111010100000101110110101100000011100110;
#1 $display("%b", po);
# 1  pi=207'b111111011001101000100101111111110100110000011101000101110010010111000010000011101111000001100010000010101110101101010001011100101110110010000001001010100000010101101000001110011010010110001110101000000000101;
#1 $display("%b", po);
# 1  pi=207'b000000010100011010111110101001100110110011101101011010011011111101110100011100100111101011110001010000100010101011100001110001101011000011100011100000111111111010101011000100110110111000000000110011111110000;
#1 $display("%b", po);
# 1  pi=207'b111011110000110011101001100111011111010001111100101111110010011010111001011110101011010000111011001100100011011100000011000110000000110111110101100111111011010101111101101100100110011101001110010100100111101;
#1 $display("%b", po);
# 1  pi=207'b000110001100000011111101111110100001101110011000100111001011100000100101000000101100110000000010001000011010010001111101000110100111001001110101100000010110110100011010111100000011011000001000111111011010101;
#1 $display("%b", po);
# 1  pi=207'b101011110110001100110111111011011111001111100101101101011111110011010011011000101111101111000010110111110010110111001000001101100001010110001101010010000010001110000001101001011011011111101100101101101011101;
#1 $display("%b", po);
# 1  pi=207'b100111100110110011101010010011000010101010101010010001111011110010000100110101010101010000000000100011000110010101100010011100101111011010001000101011010011100000001110011010000001000011110110110011111010110;
#1 $display("%b", po);
# 1  pi=207'b011110110101010101011111000010100111111010000100001101001011100110000010000110110001010101011100101011001001010011010100100110000010110000000111001100110111010111110010011100011101111100111111110100000000101;
#1 $display("%b", po);
# 1  pi=207'b111111010100101000110110110011100101010001010001110110001000010011100101110101001111110111001010000101101110100010100101001110100101110010101101010100001101111110000110100000000110101111100000001111111111101;
#1 $display("%b", po);
# 1  pi=207'b100011010000110010001101001101011010000011100101110111100001011110101100010111100011111011111111101000110011011100010111010110010011011110100010001011100100001111010010010000000100001010010101100110001000110;
#1 $display("%b", po);
# 1  pi=207'b111000110001010010111000111100000000101011011110001000000010011111001001110011010110010110011010101111010010100111110100000111011011011010001000010101100011011001110011100001000000000101110111010111110001101;
#1 $display("%b", po);
# 1  pi=207'b110001010010101010110011010110011111010011101101001001001101111100011101101101010010011101011110001110110100110111111010100010001100100101111011110100010100000100101101110111000101001000001111001101001110001;
#1 $display("%b", po);
# 1  pi=207'b001001010011110111110011001110011101111000000110110001011001011111010000010000001101100010011001110011011001100110110011010110101010110010001101110110010000011111110111111100100011010001101100100101010010001;
#1 $display("%b", po);
# 1  pi=207'b011101101011010010011011000000000100110010111000001001101011000111111110001010100101010000001000010110111100011010001111000010101100000100001110001000101100011110001001111011011100010110000101011010011001101;
#1 $display("%b", po);
# 1  pi=207'b010100110111110001110110011011010110011001111101010101110101111001111001001101010101110011111011110110011011001010110000110011100100111000000101111101100011001111111000010010110110101111011110100100111000111;
#1 $display("%b", po);
# 1  pi=207'b000010101110001101111001110101010000111000111000100011010001000001010000101101100111011110011100111000110000111010101110011000110110010001000000010011111100011000010000001000000100101010011011011000101101001;
#1 $display("%b", po);
# 1  pi=207'b110001000000011111010110110110100001010110111010010111000000010111100000100011000011011001101000010111011000110100011011101110001010001101110011111110000111011001001000100011010101010110101111110101111101011;
#1 $display("%b", po);
# 1  pi=207'b111100001000111001000100000000001011010100011011010110011110011111101000101001000100000110000111011010001101111111101000001010011111000111111101110001011010110011001010001001000000001101000000111100011100100;
#1 $display("%b", po);
# 1  pi=207'b100001001111000101000110011100101011010110001001111011000010000010000110100011111001010101001001011011000010001011110000110011011110100111010011101001100001101001001110110000000101011000001111011011111001100;
#1 $display("%b", po);
# 1  pi=207'b000011111000010100100110011111110110101010110100001100011000111110011100111010010101000101001111111001010100010101100101001101100010011000010101011101110001010011001111001101010111001000011101011011001010111;
#1 $display("%b", po);
# 1  pi=207'b110001111001110111000100110110110110001000000011001101000000101101100001101111101111111101100001011010100000011110111001110101111010101111000000001101100110001100110011100010010101100000001101110111110111010;
#1 $display("%b", po);
# 1  pi=207'b011110110001011101000010101101011101011101111010010001000000001010100110000011110111101110010101100101111001100110001111101011100101100010101010001001110111000010010111011110010011001101110111110001100100100;
#1 $display("%b", po);
# 1  pi=207'b000101011110100000000011110101100110110110000100110010110111000010000100001011101110111010000111100110100111111010001011001000010010010001101001010101110010101101001110110110011011000001101000010001111010010;
#1 $display("%b", po);
# 1  pi=207'b101110110110011000001101001111000111001011110000000001001001000100000100010001000110110000010001000011001010110101011110100101010111101101011010001010111100011101101110100010010000100000011110110110101010001;
#1 $display("%b", po);
# 1  pi=207'b000111101010011110000010011011110110001010100101101001000000001011010011100111101110111100011000110011110100100000001111010001001110001100001001110011011000111001011101110101000101001000110000011110110110110;
#1 $display("%b", po);
# 1  pi=207'b001000101111110011010110110101110111100110010110010101001111000110010011011001011101101010000000111101000011000011101001110100010111010100111011000111001100010001000011001100101011110101110011010001100111011;
#1 $display("%b", po);
# 1  pi=207'b001111000100101110100011111101111001110000010101100000100111000011000101101101111001000000010110111100111111010000111101011101001010100001101101110111110101000011010111101101001101111111001101101010001101010;
#1 $display("%b", po);
# 1  pi=207'b100000010000010100010011110001111000001111000101111000011011011001010000000100011011011101000111100100101100010011111110001111011001111001110110110000100111001100010010001110001110100000010111000001000110001;
#1 $display("%b", po);
# 1  pi=207'b000010101100100111101010111001111110101001001101110001101011011011010101011011011100110010111000101111101100101101001000010110010001110101110000110111111110010101001100111101101100100010101010001111010010011;
#1 $display("%b", po);
# 1  pi=207'b111001100110100101010111010100100011000100111111101000110101000001010010110101110100100110011010100100110001100110001110001101111110110001011111100010001000001110010100000111000100010110010000110111011001110;
#1 $display("%b", po);
# 1  pi=207'b001000110011010100110100010111110111011101100001010100001111011001001101111101011111100000111100110010101111011100101000110010100101100011111010101100111001110000000010111100101110100100101001111111010001111;
#1 $display("%b", po);
# 1  pi=207'b101000001011011100100011101010001010010001001000011111010111010001110001101000110000001011100010101110100011100011000001110111100010001111100100001100110011111110100111000101110001011111110101010011101100110;
#1 $display("%b", po);
# 1  pi=207'b100111111011111011001011101100110001110011001111000110010010001000011011100010001101001010000110111101101001011000001100001000101101000101000100011000110010100001010100110011101001101110100011000111000100010;
#1 $display("%b", po);
# 1  pi=207'b001101110111000100101110111011000111011110000111001011110000111101111100100111010110011110100001101101010010011101001110100011110111011001010101110010010011011010010100110001100010001011100110000101001010101;
#1 $display("%b", po);
# 1  pi=207'b000010001010000110100001111111011100111101110001100000101100100101001001110100110000101001000011011001010011011000111111011010110110111111000011101110001110101000001011101110101010010101001000001101011010110;
#1 $display("%b", po);
# 1  pi=207'b110110011111111111010100011110000101001011110001001010111100001011011111100011101101110100100011100101010010100010000001110100101110011110000000000001111001101011100100010000000100100011010010100100100100100;
#1 $display("%b", po);
# 1  pi=207'b100000101110110010011001101100101010101011011101001100101001100010110001010100110100110010010110000100010111100101011000011001010101001110010101100000101111000101101010101100010001110011011101100011100010001;
#1 $display("%b", po);
# 1  pi=207'b111110011001101001110111111110110010010010111010110010110000011000110011100011001001100000100001101011001011011010100011101000010011011011110000100010001110000010000000011011000100111001100001111001010000000;
#1 $display("%b", po);
# 1  pi=207'b000010110010010101001001100001001111100101101000101100011101101010111100111001111000001100110001011111010101011011001001010101101000010011000011101000011101100110001111000001001000011010101000011000010101001;
#1 $display("%b", po);
# 1  pi=207'b101010010000111101100010011001010011010110001001101110100011110001101100101111000110101111110010111010011001111000101010101001010000010011100101101010011110001110001010001110111001001001000111010111010011100;
#1 $display("%b", po);
# 1  pi=207'b011101001110000101100110110100011010110100010101100101000010000000010100001100010001000011111001101001100110011110110010011100001001110000100100111110101011001101001111000001001000101011111100010100011000111;
#1 $display("%b", po);
# 1  pi=207'b000101010011111111100011100111011100010010111101001110000011000010010111000101101111110000111010101010101100010010111101010101001101010010100111101010001100001011100110001111111001110101001101000010100100000;
#1 $display("%b", po);
# 1  pi=207'b100101010101100111100111010100001010000001010011010000110000100110010110010000111011001001000010000111110110010000101101111010010011100100101011111001011010001100101000111011001000111000110011010101000011110;
#1 $display("%b", po);
# 1  pi=207'b000011101101001100011000011111000111010110001001010110010001111011001001101010110111010011001000101110001010100000101110110010100010101111101110001011110100011100101100000001100101000100101110010101111000001;
#1 $display("%b", po);
# 1  pi=207'b000111010011000110110010110000011011000101111100100010100010111100011010010100001011101100100111001111010001001010101100110010111100100100110010011000111010011100000101111110011110000110001111001110100101100;
#1 $display("%b", po);
# 1  pi=207'b000000010100000001101101000110110111011001011010001010001110010011000001000000010101100100110101001011010000001101110001111011000101111010001101101111001011111101001110000110010101010000000011101010100011101;
#1 $display("%b", po);
# 1  pi=207'b110111101101000011011011000001110111110110001001010011101010110101001001000010011101101011010001100011010111000110000110010100010001100000011011011011011101010101101101110110110010011101111001110011001011011;
#1 $display("%b", po);
# 1  pi=207'b001011011111000000100110010011011111101000001011101001001001001010000111111101001101000111110101000011010011100100010000001010011100101001100111110011101111000110111111000000000000100011100111010001011001000;
#1 $display("%b", po);
# 1  pi=207'b011100101011111101001111110110110100111100100110111011101001001111110100000100100101000100100100111101100010001011001001100100100000010110101000100111000011000101010001010000110110011010011111000010110111010;
#1 $display("%b", po);
# 1  pi=207'b011010100101101111110101110110010111100001110110110001001010110111001011001111011100011111010100010000011100001010111100001110010001011010111001000111101110011111010101011011000111111110101101001011000000000;
#1 $display("%b", po);
# 1  pi=207'b011100010001111011111111111000110100000010111001001001000111000110010001100100010101100000100110011000101001011011010110011011011000011000000110111011001001110001110101010111011000111100110010100100101001110;
#1 $display("%b", po);
# 1  pi=207'b000011010101011110001000001100101011001101101100000111001100011000101010011010011111001001110100110110111011000010011011100101010101101110111000100010111110100111011011111110111101001011011101011010110010011;
#1 $display("%b", po);
# 1  pi=207'b111110010000110100011001001111001011000110000001001110000000011000100001100110001100010001100111101111111000111000000110000001000000010110101100101100110110001011110100111101011111000110011001110100000110100;
#1 $display("%b", po);
# 1  pi=207'b001010111111101110110010111111000000101110100001010011001010110011101101110110101100000101110110110000000101011011111101110101100110000010110011100011111001100010100001110000100110001010100010110111010100011;
#1 $display("%b", po);
# 1  pi=207'b100011111010110110110110000011101110001111001001110001011100110001010101110101000111000010000110111010010001011110011100001110100011011011111100001000101011000100101110011100001000010010001110110100011011011;
#1 $display("%b", po);
# 1  pi=207'b010110101010111110000100110110010101110100000011101101010010010010101010111111000011110111110111110001001110111110110000111011101010111001111111111110001000100101110000100010110010011100010011111100001000111;
#1 $display("%b", po);
# 1  pi=207'b110000001111011111001000011001110100001101001011000101011111100110010111010011001001111110111011001100011101011001010000110000000100110101111011100010010010101100111101000110011011000111010111100001011010100;
#1 $display("%b", po);
# 1  pi=207'b110101011110000111100110101110001110010100110100111110011100100000111111011110100101000111010101101101111101111001000101001111100111010100000001100100100111000001100000011111011000001000111011100101110100101;
#1 $display("%b", po);
# 1  pi=207'b100100010011110000110000101011100010101010101000111101010010000101110010001111011000010110111111010000011100111101110000011000000111110111001111011100001010101111101110110001000000010000000010001111010101011;
#1 $display("%b", po);
# 1  pi=207'b011111000000011111100101111001010010010000110010001111110110110101011000100111001111000000101100000000000111110010011000101110011011100001001111011011011000000100100001111111000011110101101000001000101011000;
#1 $display("%b", po);
# 1  pi=207'b100101000101100010101101011001011110011101110100111001111110011100100011110001010011011000001000100010011001101100011000011101100110000110000100000011101111010011110110100011011101111001011001010001010000101;
#1 $display("%b", po);
# 1  pi=207'b111001000000111001010000111111000001101000001111000100010100011000010011100101001101000100100100001110011111001110111000011110010010011011000100010100110010110100011101011000011101011111100011010110111111100;
#1 $display("%b", po);
# 1  pi=207'b100000000111110011110110000010111110001110001011010111011101001101010100101000101000111110010011100110011111000110101000100111001000100010111000000001100011000001101100000010111111101111001000111110111001110;
#1 $display("%b", po);
# 1  pi=207'b110010000101111010010001100110100000100011101111111101001101111010100101000001110000111100000001001110001110001010111010100110001110011111110001000010001100010011110011001000000100011111010000000100100111001;
#1 $display("%b", po);
# 1  pi=207'b000111101000111010001000101111010011010001111110001011011001011000111010110000111010110110000010001011111111111111010001010100101010011110101111100011011011101010010010100011000011010010011110101010111111000;
#1 $display("%b", po);
# 1  pi=207'b011001101001101100100111111011110111011111101011100110001001101110010110001100011101001001111011110010100101011010111101111111000000110011100010110000001011001001110110000110110110110011010110010000011110100;
#1 $display("%b", po);
# 1  pi=207'b110100111001111000010100111010001110111010010110011100111010111100100100110011100001011100110010101000001001100100111111111000010110111010100000010100111100101000011001001001001001111011000110000101101101001;
#1 $display("%b", po);
# 1  pi=207'b111100000100101101000011101010000110111101100011110111101100001101110000010111101011111100100101101101110101011110111111100001011100011011000100100110000011101111011111000011011101000011111010110100010001111;
#1 $display("%b", po);
# 1  pi=207'b001110000111010000111100100101110101001101010110110011010101011101000000110011000011000111110111110001101110110010111001011001101001111011101101100000010111100010000101101001011010101111000010111011110110001;
#1 $display("%b", po);
# 1  pi=207'b110110100010111011111000100001110011010001001001001010001111000101000010010001011000100111001011110000100001110100001110110100101011110001101100100000111100001111001010111100111111011101010100111111110111010;
#1 $display("%b", po);
# 1  pi=207'b001010111010000100000001001110000000100001101001000011000001011000010001011011011001101101101110111111111000101111100000101110111100000101100010101101011000111111000000010010110111101111010110001000111101010;
#1 $display("%b", po);
# 1  pi=207'b001101111111101000010101001111011110111101000000101110111000101110110101110111101010101010101110000011011110011011011010111001111010000100100110001000100110111101101000101010010010001110100111011111100011100;
#1 $display("%b", po);
# 1  pi=207'b111101100011011001110111011001111000011101110000101111001011100111010101101110011011100111100011111000101001101010101010111000100010010010100011000000001011001001101101000000000010000110101101110001010110011;
#1 $display("%b", po);
# 1  pi=207'b011101010011000010110011110011110010101000111111000000010111101000001011011000111011100101111001110100101001111111011110100101000111011101000111101100110101000001010000011000110111000000100111001010001010111;
#1 $display("%b", po);
# 1  pi=207'b001111101100010100111010100011011011010000010100011001001001000000101000110000010011000101000011011110001011110110010001001010110100001000010100111010111011001100010111011101100111101001110010100001011101111;
#1 $display("%b", po);
# 1  pi=207'b111011110000101110111010100110000111010010110010001010011100111001001000101101110100010100101010011000101110001100111111010111110100000011101111101110111101101000010011010010111111001100110100100111000111101;
#1 $display("%b", po);
# 1  pi=207'b100011101101010000001101100100110100001001110110000100100111101110110111110110001101010000010010001111010110011010010110101010111011110011100000110110101110101101101011010011100001110010011011110010001000111;
#1 $display("%b", po);
# 1  pi=207'b010101111011000011001001001001110111011010110000001111100111111110000000110101011011101101001000110001110010111001010011001001110011110100000111100100100111100010111011011110110011011000001001100110010001111;
#1 $display("%b", po);
# 1  pi=207'b110110010101000001010101000011111110011000100011100010001001110010010001111100101100110011101011001010011110101111101110011110011110011001101010101110001000000101111100111001010010000001100101110110011010010;
#1 $display("%b", po);
# 1  pi=207'b110111101110000001110000001011111111000101011100001000011100100100010111011101111101001000011100011010100011001011011110010000010111000100111101010010101011111001000101010101110100011011100011001000001000011;
#1 $display("%b", po);
# 1  pi=207'b101101000000110110111010001000010011001011111011000000011000100011010001011000100101001101111111101000101100001100011101010101011000001000101110011111010111110000010001111001110010010000010011110110010010101;
#1 $display("%b", po);
# 1  pi=207'b001110000100101010100110000110101111011111110110011011100011011110101000011000011100011110100001110011100100011001001010100100000100001010110101000110001000001000110101010011000111000111111010110001101010000;
#1 $display("%b", po);
# 1  pi=207'b111110110010010011010111111111100110110100001001010000101100011001011000101000000010111111110111000001110001001101101110010001101001100110101100110101001010000111011101111010000110011110111011100110110101001;
#1 $display("%b", po);
# 1  pi=207'b000101100111111011010101110000010000101100101001011011101011000000110001000010001011000100110111010000100000110000001000110110110001000111001001001001100110011010001100000100010100011110010001001001111111110;
#1 $display("%b", po);
# 1  pi=207'b010011101110001010001001000100000011010111001111100001100100111011110100111100011100100001001001000111010101101000111010010111111101110110111100010101111110110101101010100111000101010011101111111010011110100;
#1 $display("%b", po);
# 1  pi=207'b001000011100001011011000010101100100110101010101100111000101110110110110000101000000101001110000010001000110110000100011011011011111101000100011010000100101011110010101100100000100001011010111110101111111100;
#1 $display("%b", po);
# 1  pi=207'b110111100101101011000110010001100100011100100110111001110001101010011000101100100100111011110010001001101101000001101000101111011110011101011011010111101011111110001000011000000010011101111001101010101011001;
#1 $display("%b", po);
# 1  pi=207'b111110101111010001110101010011010011101111000110001011001111110111001101010000001010011101001010011000010101101000110010011101010001110101100001111000100001011011010000010010011001010101010101110000110101010;
#1 $display("%b", po);
# 1  pi=207'b110000000011100010110101001100100001110010110000100010000010100010100101110110110010010101001101011100111001111011110110000000101101001001111000010100111110110000100010101100001000101100110011010000111100100;
#1 $display("%b", po);
# 1  pi=207'b111100010010100000101010110000100111100000010110101110010110100111011101001001110100010101010000011001001101011111111001100100101101000010110010100100010010101011001110110111101000011100101111011001010101011;
#1 $display("%b", po);
# 1  pi=207'b011111010111011100010111000010011111010000011001011100010010100111100000110110110000100100000100010101000101000001100111001010011001110000101000000101110010001100100011010110101111010000100000101111000011000;
#1 $display("%b", po);
# 1  pi=207'b011101101001011110011011100011010000010001000111100011001000100000101110111001000100111011111110111110011111010110011010111000011011010001010000011000001110101000101110111101010000100001110001011001000110011;
#1 $display("%b", po);
# 1  pi=207'b010110111000001101001000111001010101011110001001110110111100110100010010011111100100111111111110101010100101110000001000011000100010111000100010011101011001101101010000010001010101111000000010101001111101101;
#1 $display("%b", po);
# 1  pi=207'b011111100111100111010100010111110000110001001100100000111100001001110101000101010000101110100101111101111101101011111010100101011101011110000110011010100101100101001011101110110011100010101010001110010110001;
#1 $display("%b", po);
# 1  pi=207'b000101110101011111100001101101111110010111100100000111100111110011100100000101001101101101111100011110101001111000100010001000000001110000000001101001000000011011010010101011110000100000111111101111101100110;
#1 $display("%b", po);
# 1  pi=207'b000011111110110001011100111100101101011100101001100111100010110111001100110001011000100001010111010111110101000010000101011010111001001101100110000111110101010101111111011110000001101111101001100010111110100;
#1 $display("%b", po);
# 1  pi=207'b011101001000011011111111010110101100110101111011001001111111001111100101011010000100010110000000010001011000001111100010010111101111101001110111010001010110111110110000111111111101010001001000110001100000111;
#1 $display("%b", po);
# 1  pi=207'b001000000011111010011100000101000011011100011001100100110100110000010000101000010111101001010000010000011000101010011111101010011001000111011001010011101010100110110011111011110110000011100111001111011110000;
#1 $display("%b", po);
# 1  pi=207'b011001110010010100110100011110100110000111001110100010001101100010101011101101111001000101111101110111101001110001011110111010110111110101011101101111001110101001011111110010000000100101010000001011100101001;
#1 $display("%b", po);
# 1  pi=207'b111010101101111000110101101011110011000000001000001101101111101100010111011001110100001111000001110100101010111111101111100101000001111111011110000001101011001100000011100000001101001100111011111000111111110;
#1 $display("%b", po);
# 1  pi=207'b110100001000010000100101000000100000000000110110111100000101110011110011100111000001011101101110010011000001110001011000011101011101110111111110111101011111111011001000111011110100111001001010101001000011011;
#1 $display("%b", po);
# 1  pi=207'b001010000010010101000101110111111001101101011001011001001111000010010101010010001101011011100000001111010011111010000000001100000100111001111010100100011101000111011010111110101101010010001011110001100100100;
#1 $display("%b", po);
# 1  pi=207'b000100111001111000001011101110010010111000111000011000100101000111110010111001011000111001010001011011010000001011100001100000001001111110010011110000110101101110100111011100010001100101011100100101000011000;
#1 $display("%b", po);
# 1  pi=207'b010101011011010001011001100101011001000000111011011110100011101010010101010010110000001011010010111001101111101000100110110001100100011010001110011110010111000101000000011001000000100001111111101100101010000;
#1 $display("%b", po);
# 1  pi=207'b101101100010000110001010111000110101110010110110000001010110011000111010001001000010100010010000010111011000100000011110010000111010110100110011000001001010110110001100101010101101001010011111010110010110111;
#1 $display("%b", po);
# 1  pi=207'b100010001001001100000110100111110001010000100010101111111011001001011000100011111011001110101101110011111110010110100110110001111100101001011011011101011001011010100010100011010111101101110010100001110110000;
#1 $display("%b", po);
# 1  pi=207'b101110011100000000011001100010001001001011110000100111101111101111111001000101001000011011100010100101001011110000010000100111010010010100110010010101010000101101011110010111110110101100010111001101001110011;
#1 $display("%b", po);
# 1  pi=207'b001001011101000011011110010111011110011001101110001100000101001000111001100001011111111101101100001001000111000110000010110111111101000111101010001111101011110101111000010101101010010100000110100000111000100;
#1 $display("%b", po);
# 1  pi=207'b100110010010011110100000100001101010000111011100010101100010010001111001110110011000111011011000010111001110101110000110001001001110110000011111001001100011010110010101010111001110000000111011111100000101101;
#1 $display("%b", po);
# 1  pi=207'b001000001011101001100100100001110101010100111110110101101000101110001111100110111100011011001010000100110011111010010101000100101010110101111111111111011011010011110101001001010001111100100110111101111101001;
#1 $display("%b", po);
# 1  pi=207'b001000001011100110000111000010100110111110010100011111111101100011101101111001001111110000000001110000011011011000111011011100001111000110000001110111011010100110111001010000011111100110111100001110111101100;
#1 $display("%b", po);
# 1  pi=207'b100110000101000001101111101000110110000110101110001111010000000111100100001110101010101011100000100001010001101000011010010111000000010110110101000010001111000111101011010010010010010011101101111110011110000;
#1 $display("%b", po);
# 1  pi=207'b000011001000000111001000111110011111100100111001011111101000110111011111111010100101101101111111111001101001100001111010101110110111111111001001101000010001100010101000011101111001100111001110001100111010011;
#1 $display("%b", po);
# 1  pi=207'b111001110110000100100010001100001110111100100100100011111111000111001000001001100010001100001111101001011100110111111001100101010111110000101101001111001100110011111111000110010110000011010110110010010010010;
#1 $display("%b", po);
# 1  pi=207'b101010000101101001000100110111111011111011000110101110110011110011111010101111100011000001100100011001100000111000110011110001110010111111011110101011001110011010001010010111100101101100110001011000110011110;
#1 $display("%b", po);
# 1  pi=207'b010010010101011011101011011000110110100011110001110010001000110010010000111011010111011101001011011100000110010110111110010110100101011110011110010100100010100010100000110101111111101110000011010010111010101;
#1 $display("%b", po);
# 1  pi=207'b101010011000101010011010100001110011010110110011111000010010111110100011010010111101111001011101111001001010100000001011010010010000000111010011110111010100100010110001110100100100010011100001001000011011001;
#1 $display("%b", po);
# 1  pi=207'b011011101010110101011010000100011110100110001111111111010100111001001011000111011101101100010111100001001001100001011100111000010011001101100001001011000100111000101100000001001111000101011101110000111111011;
#1 $display("%b", po);
# 1  pi=207'b111010101110110011001101001011100100010111001110111111111000010010011001011110011010111101001100010010100100101101000100000011110111000010111001111001110110000100110000110011011110000100110010010000101001011;
#1 $display("%b", po);
# 1  pi=207'b010111011010101110101100111010111010111011001000000110001111101001011100001100010001100000011011010000010101100100011000010111001110001110110011011011000101011010110011111010000001110101011010000100101110001;
#1 $display("%b", po);
# 1  pi=207'b101110000100111011100100011011111111111000001001010011100101110011010011111110001100100011000110110111011111011010010100110011010100110001101011111011110010111011011101010011101010101011000000110010110011111;
#1 $display("%b", po);
# 1  pi=207'b101010110111100110110010011110101011010001100100011011110100110111110100111101101101010101011110011001101101101010010101101001011100101111110011100000111111010001000011111110110010010100101000101001100100110;
#1 $display("%b", po);
# 1  pi=207'b110001100001101010110011110000100100010010110110011100111000011010010010110000100111010101110011000000001001110001100110100010100111100001011111101000110111100010101010111000001100100111101001111000011001000;
#1 $display("%b", po);
# 1  pi=207'b101011011001111101110001110111101011110111001011111110010110111110111111010110100110011000111011001010101011000111010011101101100010000101110000001100000000011101110101011101010111111100111100110001101010111;
#1 $display("%b", po);
# 1  pi=207'b001000110000111011111010110101011100110000010100010100101000100111110000110000101010011100010100011001010000101100111110010101000011010111101011111001101000000111010111101101010101011100011100100100010101111;
#1 $display("%b", po);
# 1  pi=207'b100110101000001110001110111011001001010011000000001110111100010000100001000011110001011111101011101100010011001111010100010010101010101111000110111110110110111011011111000001001101111100000011010001101101010;
#1 $display("%b", po);
# 1  pi=207'b101010001101110000100101110001000001110100111000001011000010110000001000010110010101110010001001110001111001000001100000100101100111111001101000101000000000001110011101111011010100110010011100111110100001100;
#1 $display("%b", po);
# 1  pi=207'b110111010000100111010100001000011001001001111101111000000101001100001010010010100001010011111001111101011100110001101010111101010010100001110010100110100110101010110011001010011001101110010100111000001110110;
#1 $display("%b", po);
# 1  pi=207'b010011000000101111111101010001101000101100100011011110011011111001001111100000100000010000100001101000001000010100101001011101101100001001111001001011010110110101110010001010100011111100001100001010000100100;
#1 $display("%b", po);
# 1  pi=207'b001110111100100110010000111010010011100000000001001101000010011011000001100101100110100011010110110010011101101000110011110100101011011000001001100001011011100010010011010100111110101100001110100110101011001;
#1 $display("%b", po);
# 1  pi=207'b101110100111110000111011101110110101101100010111000111110110010011001001101001010111111010010000101001010010111001100100101110000101001010010100101010001010011110101001010110000010001101100010011000001100011;
#1 $display("%b", po);
# 1  pi=207'b110011010000001111110111101011101101010011100010110101101001110011100110001111010011001111001110011111110000101100001111111001111001100111111101110001000000100111001100001011010111100100110110011001110110011;
#1 $display("%b", po);
# 1  pi=207'b001111000000011000011110000001011111110111101000000011011011000111101100101000101100010001000100101000010011000000001000011100011001001011011001100000010111000100111010010111101100111010000000000001101010110;
#1 $display("%b", po);
# 1  pi=207'b110111011110111100100011110101000000100001011110010111100100010101110111101010001001101101011000110010010110000000110101010010100010010001010110110101111011100100101010011001010000100001111001001011100000010;
#1 $display("%b", po);
# 1  pi=207'b111011110011110001001000010000100101110011101100001011001010001000101100010100010011111101100111001001011011001100100101111110100100001100110010001011101000100010101001000110010010001010110010011011111111011;
#1 $display("%b", po);
# 1  pi=207'b100101110011010101001010000010100000000110000010000010101111111100011000111000001010111010101010010011111100101001011111111111000001010100101111100110010110111001111011001011100010001001010000101000010011100;
#1 $display("%b", po);
# 1  pi=207'b111111110001001111011100100100111010011001110011111010110010111111010010001011100001011000100100010101001001010111110110111101001000010001000101011001110010010101011001001000110111000111101110100001101010010;
#1 $display("%b", po);
# 1  pi=207'b100011000000100010010011100111000111101111001100000010101100001011000011101101111001101111100010010010010100001000000100111100100111101101110100111111101000000101101101000110001101010101000100100010111101101;
#1 $display("%b", po);
# 1  pi=207'b111110010010110101000101001100100001010101011010110000101100011000001110001010011000110010101111010010010101000100101010100010001011110110111100100110001111111000111011001111110000110001011011110000100011010;
#1 $display("%b", po);
# 1  pi=207'b000001111000101010101111000001101001110000011010101010111111111010011110000001010011110110111000010010110100001000111011110000001000001110000111101000100001110110101111110100001101011011111010110001100000000;
#1 $display("%b", po);
# 1  pi=207'b001010011111000001000010110000010000110110111000001100000010010001001101100101011011010001001101101000011101000010011001001100001000000100111110100001011000011110000111110000111011101010011011000100110111001;
#1 $display("%b", po);
# 1  pi=207'b110000111110000000000111011010110110010101111001100000001010010111011110000101101001110000011101011011111011110110100111011011011111001011000101110111001000011110101001110110011011111001000001111100010101000;
#1 $display("%b", po);
# 1  pi=207'b000000110100111111010011010010110110101110000001101111111010101001100001110000001000111101110110110100101000100110100101000100111001001111011101111100110101001100011011110010000111010011110100110001000100000;
#1 $display("%b", po);
# 1  pi=207'b011101011010010000101111010110100111000111001001111111010111000011001101110111001111010010111010010001100011000000001010111101101000110100110001110000101011101101101111000011101011000010011011001110010100010;
#1 $display("%b", po);
# 1  pi=207'b101000001010111000111010111110011101001101000000000000111101000111001110000101111000111111100101010110101101101010110111101000010100011001011000111010001101101000101100100000110100110010110001101110000110010;
#1 $display("%b", po);
# 1  pi=207'b111110101101011100001000101111001000000011011010001101100010110011001011101111010011001110111111000010111001011001100010010010111010011000001110111010011111111001110000011001101010000001011111101110010010101;
#1 $display("%b", po);
# 1  pi=207'b011010101001011100100101001011001100001100000101001001101011001001100111011101101001010111001010110110101011001100111111000110000011011111110110000100010110010110100000111011111111010111110011010111001011111;
#1 $display("%b", po);
# 1  pi=207'b001110001100110010101000100111110010000001110001010010001100011100010011111001110101111111000000010000001101110111101000001111110110101111001001110101001001000010011111111100111100100001110110011010101100111;
#1 $display("%b", po);
# 1  pi=207'b001001000111100001000000111011000000101111000101100111101011010101010011011001101000111100110101110100011010010100100111001010011110110100011000011010101000111000111001101110010011111111001001101101010001100;
#1 $display("%b", po);
# 1  pi=207'b010000010000111111100100010011001011111101010110011000101111011000001111110101101110110000000001111000011011010110111111101010110101111100100101101010110011111110000000101101100011010111011000110101111010000;
#1 $display("%b", po);
# 1  pi=207'b111011110011100101000111111101111011101111101111111101011100111000101111110110011001100001110001100111111111010100010100001001001010110000110110110101101111100110111100111000110111011010001111011011011001010;
#1 $display("%b", po);
# 1  pi=207'b000110111001111111011100111000011110011101010110100000100000111110001001100111111011110110100100001001110100000111001110111010111111111100101110000100011000100110001001110010000111000011110001000000111001000;
#1 $display("%b", po);
# 1  pi=207'b010001011110100010011000000011011011010100110001001001000101011001111010100101010110110110011101001011111101110011110010001111110100011110110101000010000001110001101100011001111110110001000010111110110110011;
#1 $display("%b", po);
# 1  pi=207'b100000001010001011111111111111001110100000110111111000110100001101111101001110101101001000011100000011011111001011101101100101110100000101001001111000011110111100110010110011100010110011011001110110101011001;
#1 $display("%b", po);
# 1  pi=207'b110100010110100110101101000001101110000001100010101100110100001001011000100001010100110010101011100110000010111010100010111011010011111010101100000011111110010001110101100000010011011000000110000101000110111;
#1 $display("%b", po);
# 1  pi=207'b101000110011011101110010110010111111000111101110110010011110000111011010000001111110110010011100101001010100010001011011011001110011100011100110100101011110001010010000000001110000101000010111111111101011101;
#1 $display("%b", po);
# 1  pi=207'b110011101001101100110101100001000110101111110101101100101011000111001011101110010101101000110100110101011111000111011111010111010011100111000011011000101010101010000101011000100011010011010010110111111011101;
#1 $display("%b", po);
# 1  pi=207'b001111011101011000000001100100110001110101110001000111011100110111000101110110111001110101101110110001011110000001110011001111101010110110111011011100111010111000110000110111110101100100011110010100101111001;
#1 $display("%b", po);
# 1  pi=207'b110011000101000100011100011110011010011110110101000111011111110110010101110000011100110110001111100111001011101110010011010010100110001110101011100111101011101111101010111111011000101010001110101100000001101;
#1 $display("%b", po);
# 1  pi=207'b111011111101101001101011100100001010101111011100010111001101001001100100001111001010101011011101000010010100101001011101001000001101011100101110100000101110110101000000000010000111100100000111101010100101011;
#1 $display("%b", po);
# 1  pi=207'b000001011000110000011001110010101100000110000111011011011110100001111100010100110000011110011111101000101010110111011011001001111110011011100100100100100001110011100100001110111111011001011100100111010001110;
#1 $display("%b", po);
# 1  pi=207'b111001011000000100001010101100100111101101011000001101000111010110110111100001101111100110001101000111000011111001110110100100001000011110100001100011010011100101101110101010100000110101111001111111110000000;
#1 $display("%b", po);
# 1  pi=207'b010010010101000011000000000011010100111101011011001101110110010001111110111011110110010110111110110110101010101101101100110101100000101101001001001100101000110110011001000011001101010100111010001000011111100;
#1 $display("%b", po);
# 1  pi=207'b110100001110010111100111000100110100100010101100100111011100000111011010001100110100011111110110011010000101110110000001001101101010001100111110111100100110101001110010010011001011001000110010101010101111111;
#1 $display("%b", po);
# 1  pi=207'b001001111100111100011111100000001010110011001100111011101100010000001000000111001101001101001001000011101110101000110001101011010001101100101110100101001010111010010000100010011111101100001110010000111101000;
#1 $display("%b", po);
# 1  pi=207'b110110111010111010101111101111101110000110110111001100001110011111110100100011001101101101001001110011001110010101010000111111100100010010010000111110010110010101110111101011111011100010111110111000001111111;
#1 $display("%b", po);
# 1  pi=207'b100011101101000100000101011001101110100011101100110010101100010110010011010100110100111000110001001100011101001010110111100011110011001001110101101110101000110111101011111010111010110000010001000011010100101;
#1 $display("%b", po);
# 1  pi=207'b100101100110110001011100001000010111010101100111101000011000010011011010000110111100001011110000100010101000001001011100001110011100111101101101111111010110000110010001011001101110011100000110110100101110111;
#1 $display("%b", po);
# 1  pi=207'b010001010000101101011111101000011011101001110110101100001011010111000000111100101101101100100010101000001001011111011100111100111000101110011010110100100111010110011110010101010101000111000110000010100101000;
#1 $display("%b", po);
# 1  pi=207'b011010010111000011100011000001101000000111100111010010011010100011001011000001111000110100110011111010010110111111000111001101000000111010001000111001111100100100000101010011110100000010011010010000001001100;
#1 $display("%b", po);
# 1  pi=207'b110000011000101011011011001101101010001100010110100110101000011111010110110100000000101010001100011111011011101100111111101111101000100000100001011011100010011100001111001110110100111010011000001111111111010;
#1 $display("%b", po);
# 1  pi=207'b000100111000010100001011110000010110100101100010111000100011101101110111001010011110110001010110101100010100101010110001101001110100000000101001101000100000110100111111000101100000010001111001110001101001001;
#1 $display("%b", po);
# 1  pi=207'b000111111100011110100101100011000000000011001000011110111110101001000001010110011110011110111101111001111010100111111110110100001000010110100101110101101110100011111010010000101011111111001001011100001011100;
#1 $display("%b", po);
# 1  pi=207'b100110000100101010101111010001110010110011111011101010011110100011001000101101010100100001010100011010010100001100100110111101001011011010100001100110000011010111101100010001111011111111101110010000110001100;
#1 $display("%b", po);
# 1  pi=207'b111011110110111101001100010101000001110110001101000011010001001110110010000100111011000110001001001111100010000010001101000001011010111110100000101011111010100000010010000100100110011100010101101111010000000;
#1 $display("%b", po);
# 1  pi=207'b001000110100011110000011111111010110011111001111000010011010010001111111110000000101010000101100001101001011100000101110000111100011001110101011101010011101010100110000101001111011100000101010010000011100101;
#1 $display("%b", po);
# 1  pi=207'b001110100110111000010101101001100110110101110000111011001010010110100001001000000110101001010101100100010111010110101100110101111111111110100011101011000000110011010101100001111100110110001101011110000010010;
#1 $display("%b", po);
# 1  pi=207'b100111101111000011111011011011011000010010111011001001111100111110010101011100001101100001011001110110010110101011011100011000001000100101101010111000111010100001101010100111001010100101101000010111101100111;
#1 $display("%b", po);
# 1  pi=207'b110110100001110101110100010000100000010000110111001101101011101011101000101100011111001110100110100000100100010110001000001100100110001010000110110101110110001100001101010100010011000001111000001100010101101;
#1 $display("%b", po);
# 1  pi=207'b001100101010101001100110110001101100001011010000111000100100101111101100011100101111110110100101100000010100111111001111101100000101100001101001010010010110000110110101111111111101110010111010111111010111000;
#1 $display("%b", po);
# 1  pi=207'b000111010001010000111011011110100011010100010100111101001110110110000111010000101101010111011010001011100111101000111101000011110000011011111100101011101011011001100110010000001001110110111011110100000000001;
#1 $display("%b", po);
# 1  pi=207'b000011100001111000101010101111000000011100001100101111000000010010110010001101010111110011110101110100001101001011010110101010000110111001011100111101000111110111011101000010011011010001001100100100100001011;
#1 $display("%b", po);
# 1  pi=207'b110000011101000111111110010010010001111100100010111001000010000111111001010111010010100100100110000110011111001011110100110111011001000010011010010011000011101000010101001010111011010100001101100111110110100;
#1 $display("%b", po);
# 1  pi=207'b101001111010101101110000110110101111111010100000111000000110101011101111110111110100001110001011000001110011000101111011111111110111001101000011101110110001101000000101001001001111111110101010011101111011110;
#1 $display("%b", po);
# 1  pi=207'b111110000000111111110011110111111001011101010110010001011000111010110010000011011001101100101010000100110000101000011011010001100100101101000000000010001010100001011110011100011011101000000001000100011111001;
#1 $display("%b", po);
# 1  pi=207'b011111100100000100101101110011000111010111111110011001111001000110011001001100001100011010010000110100110110001011010000100011111101111000101110101000100000110011100000100011110010000110000011100111100100100;
#1 $display("%b", po);
# 1  pi=207'b111101011011110000110011001111100110000000001110011000101011101000100100111101000110000110110001110011101000000101010011001111101100001100010010111010111101100110110111111010110100010010111001101011000101001;
#1 $display("%b", po);
# 1  pi=207'b110101100100100111111001000010100110111101100011101100001000100100011110111001010001011010110001101110001100101011100010111111110010110011011101010101111101110101001111111110000101101010001111110111111010011;
#1 $display("%b", po);
# 1  pi=207'b100100011000000100111001000010111011001111100101011011011010010100000111000101000110011011111101111110011001000110111100100100101110000101000011011100100110111111000011110010111101110010101001000111111100110;
#1 $display("%b", po);
# 1  pi=207'b110000100111100100110110111110111111101111000000111010001010001001011001111101111110010110111000001011101000011000101110111010110101100110011001011110110110100111001010111011001110010010011100001011110001010;
#1 $display("%b", po);
# 1  pi=207'b111011001011111110100100010000111001000010011000111100011000110000101100000001000011001001001100111110001010010001100100011011111000010101001000111101101100011000100001101110011101100000001110110011011011100;
#1 $display("%b", po);
# 1  pi=207'b010011010001111110001001001110110001110010111100001000001000111110100110011001010000011100110110101111111101111010111100011101110011000101101010010110001111001001011111110010010011010000011001110101000010001;
#1 $display("%b", po);
# 1  pi=207'b000111010110011000101101110111101110110111101011010110011011010101111010001100100110100001000110011100100110000010000111101011010011000011010110011000011100000110011111111001010110010111111100000011000001010;
#1 $display("%b", po);
# 1  pi=207'b100101110100100010111001100001010110111111111100000111110110101001101110001001101010001010000111111101000110100110001110011100000000100001100010011000110010100100011000011010110001001111100101010110010001011;
#1 $display("%b", po);
# 1  pi=207'b111111111010101011001101011011010000001111010011110100010101010110001101100100110100000011001101101110110100001100111001010101111101100011010100101010000111000111111101010110010000110011101001101110001011101;
#1 $display("%b", po);
# 1  pi=207'b100000101011001000101001100111001001111111100110000111110110001111010101100100101001010001101111111011000010000101001111011001011000010111100011001010001001001101100100010001010010001110010011111011000011101;
#1 $display("%b", po);
# 1  pi=207'b001001011001111100000111100100011000100001011000110001110101100110011101011001001011100110111000011000001111010000111111011011000101010001101011010111001010001101000011010110000111011111010001001110111101101;
#1 $display("%b", po);
# 1  pi=207'b100100111101111000010010000111100000100101110100111101000011101011100001111000110010001001010101010111001100100111011011011101100101001000110111000101001011111010111010001010011111010110001110001111110110100;
#1 $display("%b", po);
# 1  pi=207'b011101110010110101100100101000011100000111110110000110011001011111110000000010000001000000111011010100010000000001110100001100101000001001011000100100000011001111110110010000011001101111101100111010010110100;
#1 $display("%b", po);
# 1  pi=207'b010010000011111100001000110010010101000111011011101010100111101101110111011011101001011101000001110001001110011000111010010000010000010101110111110111100111101110111101010110101010101001000110000011100010000;
#1 $display("%b", po);
# 1  pi=207'b111001011010011001011111101010001001001010000100101110110010111011111100001001000110110101100110100111100110010110010111001010101011011000000111101111101101001000101001001100011010100111100101010011001100101;
#1 $display("%b", po);
# 1  pi=207'b011100000010111010100101110011100110000111011001000000100001100000100011101111000011011111000110111001110000100111110000001101111011001010111010101001100110010100011010001011011000101100100101111101101010110;
#1 $display("%b", po);
# 1  pi=207'b101100011100001011011011111110101110001000110010001011010011110100111100101110111001011101010011111001101110100001011101010100010010110001000100011111110100000111001110011011111000100010111010111001001001101;
#1 $display("%b", po);
# 1  pi=207'b110000011010110000110100101101000110110101011010001011100110011010101101110011101111010010010001010000110110101101110010010100101000000111100110101110000100111001110011101100110111111111000110010000001100011;
#1 $display("%b", po);
# 1  pi=207'b110100101011111001110011000010110000110000010001100010000000111011100001000010001110001110011110010101010100000010011001101111101100100011000111111000111100001000101011001010011000001000101000111101111101101;
#1 $display("%b", po);
# 1  pi=207'b111001011011011011011110011101110111010010100001010010100000010000010101000110110000101001110000110110101001110111110111101011101100000001000011111101011000001110100001010110111000011111111101111101111000111;
#1 $display("%b", po);
# 1  pi=207'b111110101101001110101111011011110000011101001011111011111111011100011100000111011111111011100111111101110010101110011011111101000110000111010100010101011010100011000100110111011010100001101111000011111001011;
#1 $display("%b", po);
# 1  pi=207'b001001010101101110001100101100111110011110011011000010101001101111111110101001101111110001010011101000110110110100111011100001101000001010101111101110101100110001110110110000011101001001001000101001000001000;
#1 $display("%b", po);
# 1  pi=207'b101111111000101111001100111011001111110110000000001001100001111100011011011100101010100011111010110010000001101000010010001100010101110001000101010111100010111010000001010110000100111110100000011001000100010;
#1 $display("%b", po);
# 1  pi=207'b000010110101110011100111001101100100011011100110100000101010111110111010110100100010001010111001101101000000101011111000001110110011110110111100000010011100000111110111111001111010101000000111101001011001011;
#1 $display("%b", po);
# 1  pi=207'b100011010101011010001001011101011001100010101001110101100010000100111000000010110011100010101101100010000111100010100011011010011100010111010001100000001010010110111011000101110111001111000000110111000111111;
#1 $display("%b", po);
# 1  pi=207'b011110000000010001110100011000100001100100000011111000110001011110101011100101100011111110100101001100111010110000111010000000111001001111011110011110000101010101101010100100010110001010001101001010101001000;
#1 $display("%b", po);
# 1  pi=207'b111001011100010100101101001101011100001101001101111000010001100100000110100011100010110000101000000100000101111011110011111111000101100111100111101011100011010011111111011110010100011011100010100011110001011;
#1 $display("%b", po);
# 1  pi=207'b101011110010101110110000111101101000001011011110010110000111011101111000111100001101111001000111001010100110101001000011001100000110111000001111001010000011000101110101110110001010101111010011011011011101111;
#1 $display("%b", po);
# 1  pi=207'b110011110011000011000000011001000100110010100011011100000100011000101000001000011011010001100010110001011000001011001011011010100001101100011110001110100100000000011000110111110101000101010101001111011111100;
#1 $display("%b", po);
# 1  pi=207'b010010101101001011110011100101011101101111000010000001010001110000100110000011111000111111010000001000010001011100000010011001011100110001100010001101000110010001100111011101110010010110001101100110010011101;
#1 $display("%b", po);
# 1  pi=207'b110100000010011010011000101011101011001100001011101100110011000110001011011000000000110010001011000110001100010001100010011111001000010011100110100111011010000001111000010110001000111110001110000001111100000;
#1 $display("%b", po);
# 1  pi=207'b110110001000101111100011001000100101010000010000101100010110111111111110011010011111010101111111001100001001111110111001111001100011111010010100100010101101110101110010011010100110001001110100001001011100110;
#1 $display("%b", po);
# 1  pi=207'b101010111101100101111101010011011110110010111100110001011100000001000110010111001000000100111001010000010000110000110000011000101111011100001101111100011010011000000101001100100110110000011001111111110111011;
#1 $display("%b", po);
# 1  pi=207'b100100000010010001111110111011111001111001111111101100011111010111011000100010111100111110111101110010111101011001100011010001010011101111001001111011001000010110101111001001011001111101010110111001110011000;
#1 $display("%b", po);
# 1  pi=207'b100101011100111110110000011000110110100111100001101010111001111011010011000010000111111101110000111110000101010110110101111001001110010110011111111101100000010111000110110111110010010100001010011000011001101;
#1 $display("%b", po);
# 1  pi=207'b101111110010101111010011100110110100111111011010010011110000000101010000101101001001100011000011001100100100101111010110011001100011000001001000000011100001110001110011111000110001001111111000100101001001101;
#1 $display("%b", po);
# 1  pi=207'b000110010011000111111111010100110101010111011000101110111110110000001100100000011001101111101011011001100110111110011110001110000011010010100011000000111001101001100101000101010001011100011010111010100010001;
#1 $display("%b", po);
# 1  pi=207'b101110100000111101001011111000001011110011001110011000110110101100111001110101111111101001000110110110100101010101000001001010000111110011111010110000111101010110111001000110011001110111110000010111100011000;
#1 $display("%b", po);
# 1  pi=207'b001010011010100000010100010001110011000001011100111001101001101110000110010111001001101100001111111010011000010010101111110110110110111000001111001001101001000101110100110000011101000111010001011101101001011;
#1 $display("%b", po);
# 1  pi=207'b011000001000100100111011000010100010110011011001101111101011101101101011010101111100100101011100000000000101101110101010010110100110100101111111100100110100010100101110100101111101001000011100101110001010000;
#1 $display("%b", po);
# 1  pi=207'b110110000111011011111101001101010101011111001110100101000011010001110111100100111011100101010011000000101010001000000101101010010010101001100000000000101010100011110100001000011000111110011001100010010100101;
#1 $display("%b", po);
# 1  pi=207'b110101111111111101010000001000101101000001001010101000101010110111100101101101001101011110111100010100110011111001100100111011110011101011110100011010001010100011010100110000000101000001111111000011011111111;
#1 $display("%b", po);
# 1  pi=207'b011011101000010011001011011011011000000011001101100111111011010011011001101110110100111111001010000101100110100000000010001010110000110000101000101010100101111111000111011011101000010100011101001010110111100;
#1 $display("%b", po);
# 1  pi=207'b111011111101001011111101000000100011111010110001001101110100101101100111100100100110000000011110011111111100111011000010011001000000100000100100000000100001011100011100111010110111000001010110010001010001000;
#1 $display("%b", po);
# 1  pi=207'b100111101001101001010101010110111011101101100110111010111010100100111100001010001000001011110111000111001101110101100110111111101000011001110010100011000011001100000101111000001100101110001001001010000001010;
#1 $display("%b", po);
# 1  pi=207'b010011001001000000101100101111101110100000111010100001101001011000000001111111100110100000001110000101100010101011111010101001101110101011100110011111101001101001101100101010010010001110001011000100001100110;
#1 $display("%b", po);
# 1  pi=207'b111101101111111010001001011110001110001001111001011100100001000000101011111110001101110111100010101010110000111000010111010011001010110100100000101001101101101011101111101000000100100000011111010100001111011;
#1 $display("%b", po);
# 1  pi=207'b011110010110111000001000101111110011000001011010101111100010110001110011000001101000110000100110100010011001011110001110010110001101101000000111000100100001001110110101011001010100111001011100110101101110010;
#1 $display("%b", po);
# 1  pi=207'b010111001001000101001011111100011011110001010011110110110000111110000010000100010010000110011110001000101001001011001110011000111110110100010010011110110110010101110100101000000001011010000111101111010111010;
#1 $display("%b", po);
# 1  pi=207'b110001010001000110100100111100110101100001001010011101110101000000011000001011100010000001010100000001001100111110100011101000000001001101100110110100100101011110000000000000101011000011100011110101111010010;
#1 $display("%b", po);
# 1  pi=207'b010110101001110111111111001011000001010011000101001001101011100001000001010000000100011100001011011010101010101000111101000011111101001001101110001010110001111000110110101001110101111101111111001101110110100;
#1 $display("%b", po);
# 1  pi=207'b111011011110111110011000010111111100000000101011001001111000111111110111111001110000011111101110010110000011110111100001010011010100011101101100110110001100000111000001100011001110001110011101100111011111101;
#1 $display("%b", po);
# 1  pi=207'b000101010110101011100101101011010100111101010110000001010010100110000010010011001100010010100000110110010001010100101100101101111010101010101000010100011010110011110001110010001100010001011101010100110101110;
#1 $display("%b", po);
# 1  pi=207'b101111101000000001010011010010110001100101011010000100100011011111101100110111111110101001111110110101101111101110000000101011011000111001000100001100100110010110111111111011011011101011110010011101001011110;
#1 $display("%b", po);
# 1  pi=207'b100100001100010010100111111111010100100100110101000100111111000111111100110110111110000010111101111010110001110010110100010110000010010001011000100010010110100110111111111010011110010000100100001000111010000;
#1 $display("%b", po);
# 1  pi=207'b000101001001010110000010010111011100001100101001101011010101010000100100110110101111000010101010011010100101000101011001011000101011100010101011011111110001010000010000010100000000101010010111000001101111011;
#1 $display("%b", po);
# 1  pi=207'b010010011001110000111101101011110110111111010101011111011001111111010011110101010110100000010011011000000011010010100101111100011101001010011010010110100000100000111000110111100110001101001011011010110110011;
#1 $display("%b", po);
# 1  pi=207'b011001100001011010100001000101110100000111001010001010111000000011001100010111000001000111011101011011000100000011110100010010111100010000111010011101100010010001101111111110000110011110010000010101001011010;
#1 $display("%b", po);
# 1  pi=207'b111000011101010111100010100001010000111001100010111111010110111110011000101000111010101010101101101001011111011100111000000011101010101111010110100011100101111011000011100000011010101111001110111100000101110;
#1 $display("%b", po);
# 1  pi=207'b011001111110111001100000010101001011000111000001001010000100001111000110111100011000100100010110111100001000000001010101101010001000110101000100100111011010111010110000110100101100101011010001101000111011011;
#1 $display("%b", po);
# 1  pi=207'b100001110000001110001001111101000011100001001000100001101101101000001101111001110101011000111001001111111010101001100110010011001001100011000110000110101100110000001010010010111000110111011001111101110000111;
#1 $display("%b", po);
# 1  pi=207'b001011111000010101001011100010011110110111101100111111100111111110001101101110001011101011011010001111111101100100001111001100101011001010001110100000000100100010110000011010001111010011110111100111101010100;
#1 $display("%b", po);
# 1  pi=207'b100001100000010101100111001000011000010100101100010000100000110010000110011000100001011010000101010111011010010010101111111001101111001010111000100010010110101101010000110001101001011100001100001001010010110;
#1 $display("%b", po);
# 1  pi=207'b001101101001000101011001010101000101010011010110001111110100001000000000101010010101110001111011000111110111001101000000110100110110111100101010000110001111000110010111010011010000011010011000101001101111111;
#1 $display("%b", po);
# 1  pi=207'b011000010110010011000010100110111001101010000101010011010000001110101000000101011011110010011001000000110100111011011010000101011101001100011010011011000110011001000100110101100010001110011110010110001000000;
#1 $display("%b", po);
# 1  pi=207'b010101001011101110011101010110101101000010001110010100010000101010110101010011000101110000001010101000010101100100100010100000110011001111000110110110001001100101100101110100101100100011010001010101011001001;
#1 $display("%b", po);
# 1  pi=207'b010100101000000000110000001010010001100001000101010011011110100010111010011100011111110110000111010110100001101011010001101011011101001110100001100001111011110011011001001010110110000010100111110001011100101;
#1 $display("%b", po);
# 1  pi=207'b011110001100111100000111100100100010111011110110000110000011001100110100001110000010100010100101101101101000111111010110110011010100010100101110101000000100001111111011001011111011000000110001111111100001101;
#1 $display("%b", po);
# 1  pi=207'b001111110101011101011011011000101010011111010110011010011111111110100110100010001110011001110001100110111011101000010011010001001101010000110110101100001100010010001000000100110001010000101100101010101010101;
#1 $display("%b", po);
# 1  pi=207'b100011011000110100100011111111101010101111111101001110011000100101100011010111010000110111110011110010110111000101100000100001000010010010110000101111111010011010001100100001011101111100011011011111010000101;
#1 $display("%b", po);
# 1  pi=207'b011101000001110110000001001111111100100010011011011101000110000010101111011110100111000001101011001011010100011011100111010110111100000011111011011111101011100001111010001001110010011111111011101100100111101;
#1 $display("%b", po);
# 1  pi=207'b110011001110000011001010111100110111100000010011100001010001010110101111110101110010100100011000011100010100111000010010000000011100111111101011100010001010000001011100011010101010111101010110011101010001000;
#1 $display("%b", po);
# 1  pi=207'b001110001100110101111101111101001110011110101110001010100100010110101111000111101101010000010101011001100110110000101110001011000011011010011000111000001111111001011111111000001111001011000000111111001110101;
#1 $display("%b", po);
# 1  pi=207'b110000111000001001110101001001110100010000010110100001001111110010111101111101110011010001000110100001101100001100110000100100100001001000000101101011001100100001111111011001011111111010111010011011100001000;
#1 $display("%b", po);
# 1  pi=207'b001000111110011001010110101011000110101101010011101001010100010101001110101000100111000000010101110000101101011100111110011000101101000100001010000000100001000010110110110110111000001000000010111111100111010;
#1 $display("%b", po);
# 1  pi=207'b001010000100000010110001111011100011011001101001110010101000100101001110011001001111100110110101111101110100010011010011100010111111000110000100011000000101010101000011001100001101011111110100101101011110110;
#1 $display("%b", po);
# 1  pi=207'b111111010110011001101010010110101011000110111110100100111000010000011101010100000000111110011000010100100101011001010010110000110011001000110100000110010111110010000110010000110110010100000001101011011111001;
#1 $display("%b", po);
# 1  pi=207'b000111011100111000001011100011110000111101110000111001110101101010001101110000001000011011001011011001000110001110101100001100100001100100000000000011000010110011110110001001110110000000100110010100010100110;
#1 $display("%b", po);
# 1  pi=207'b001101010011111011000110011100000010100011011110100101101101011011100010101111100011100000101010010100111110011011100000001111001101100011111011000101000001001101101010011010010111001010101111110011010110001;
#1 $display("%b", po);
# 1  pi=207'b111111100110100101101111010101101000001100100010000001111001100101010111110011100110000011010111111101001110011001000111011000100110011110010011111100010100110111101010000000010111001010011110100001110111110;
#1 $display("%b", po);
# 1  pi=207'b100111111101011010001010010010111111111011100011000000010011100101100011100101011000110101110011000000011001101000100011111010101101000110111001000101101100011111010111001010101110111001000110100000101011000;
#1 $display("%b", po);
# 1  pi=207'b011011001001011001011100001111111110011001100101110111010111000000110000100000101001101010110000011101011001111001010001001100010011111001000101001101111111001101111011111000010110101100011010000001111011100;
#1 $display("%b", po);
# 1  pi=207'b011000111101110001000111100010001000101001100000010001010000110101001011100001001111011100111111111010010000100000000001110010001011010101111111011110110100011111000001000011000001100111100111011011011101010;
#1 $display("%b", po);
# 1  pi=207'b010000001001110011001010000110010100100001011100101011100110011110001110101101010111011110010010111111110011110111000000011110000001011111101001110000011110010001011001101111010100110100100010011100010010010;
#1 $display("%b", po);
# 1  pi=207'b111000010011100101010111111010001000011010011101101001010100100000000011111001110100001110110100000111111110110100100110111001101100010101101001111100010100101101110111101000111000010100000100010000010111111;
#1 $display("%b", po);
# 1  pi=207'b111010110101010010101101001001101100111011000110110000010011100111011001101101011101010001000001111011101110001111000111101001010110110100100111111101001111000000111101100101010000110010100101011111010010111;
#1 $display("%b", po);
# 1  pi=207'b011001001011110010000101011010000110100000000101110111101011001100111110010011110110001000100101011000100011011010010010011010101101100110010100001110111110111100111111110111101101001110101001010000001101110;
#1 $display("%b", po);
# 1  pi=207'b100011111100101100100100101110100101001111110110000110010011000010100010001001110100110000101111010110100111110011111111100100011110100011010000100011010101100101101010101101011101000010100000100111011101001;
#1 $display("%b", po);
# 1  pi=207'b101001010110100010001101000000011110011110001011100011010101111101010000010000100100000000000011100101011101000001010001000100011010111111110111010000010011111001000111111010111111001101101100001101101010000;
#1 $display("%b", po);
# 1  pi=207'b011100001101010100001010111001001000011110100101011100111110111100001000110001010011000110001000101001001101011001110111111011100000001010011111101010111001000000111110101100000001110100101011000011100010101;
#1 $display("%b", po);
# 1  pi=207'b001001110100101001100010111000000000101110100101111100000011011010101101110100100011000000000010001000110010100011111000010111000101011110010010110000011010111100001011100011101000001000110101000000100110110;
#1 $display("%b", po);
# 1  pi=207'b010101101000001011111100101011100110100101001101001010011100011110010001011011111000101000001010101111000100011101000101111011001000000101001011000001001001000111010010110101000101111010000001010010001100010;
#1 $display("%b", po);
# 1  pi=207'b010001101100101110100001010011000111000110111100111111010001010111101100111011101101100011110011110011000010000000100110001000001101100010110010001110111010100100110100011011111000010011101011100110011100001;
#1 $display("%b", po);
# 1  pi=207'b010111010100100101001101101010010110101011101111101100010000101111010111011101110101101100001000100001101011101100111111111001100111000011000001011011001001010101100111101011110000011011100011101001010111010;
#1 $display("%b", po);
# 1  pi=207'b100000010100000110010100010011001011000110001011001110011101010110100001110010001010011110001101100010000111011001010101111011110000001100011111100001100101111011100001110011000001100110111010011010010110000;
#1 $display("%b", po);
# 1  pi=207'b101110101010001111000001010011100010100010011010001111111001101111001001110010010111010110011111001110010011111100001010101001011000111101101101100100000010010010111101100010111101000000100111011000100010001;
#1 $display("%b", po);
# 1  pi=207'b110100000011110001101010001101001001100101000110100000110001110010000111011111001110101110010000001010100001100111001000011111011011000011101011100000110100100101010011111000001100100111110101001000100010011;
#1 $display("%b", po);
# 1  pi=207'b010111110011100010011110110011110000000101100101110001110111000001111111100110011011001111100010011100101001100101100001000110001111110100110000001100000111100100110010010100011001010000111001001111010010101;
#1 $display("%b", po);
# 1  pi=207'b010111000000010110001100110100001000110011010011101110100010001110011100111111110001010100101101101111100000101110111010111000101101011100101011001100000010110110011110101010100110011001110001100010001100111;
#1 $display("%b", po);
# 1  pi=207'b001100010110111011101101111110110001001010010011111011011101110010110001101010100100010000010001101111001000000000010101001001101000010011011011101110000011111110011111110010100101010100011101001011100101111;
#1 $display("%b", po);
# 1  pi=207'b010110000111101110011101011000000010000000011001011000100000110101001101010110000111000111000110011101110101111111011100011100101010001000001111111000001011001101001110100100011011010110101110010000001001101;
#1 $display("%b", po);
# 1  pi=207'b100001011110010011100000001011110110000101100100010011101110010011010101111101011110000001110010001111100010111101100100101001000001100011100000001111100110000000101011001000111001100100000010000001000110010;
#1 $display("%b", po);
# 1  pi=207'b010001110111010101011111110001101011000001011111101000101000011111010100000100001100100101001101101110100111101010100001010101110011011101010110000010100110101110100111001001111110100110100101110001010001001;
#1 $display("%b", po);
# 1  pi=207'b010111111000110001101000010000010001010010001010000100000011010101101010010001101001001000111111100011010010010110001000101000100100001000011111110001111101101101101001001010001110101000010000011010100010100;
#1 $display("%b", po);
# 1  pi=207'b101011110001100000100100100111101111110011010100001111010011101000000010001000100110110111100010001110000110010110010001110101011011000000011101010101010101000110001101011011001101001010100101010110111000100;
#1 $display("%b", po);
# 1  pi=207'b110111011001010111011110101010110110001110010110001011110111101111100010001000101110110010001110011000111111101011101111100101010110110111010000101010000111101110101001110101111001111111110110000001101100000;
#1 $display("%b", po);
# 1  pi=207'b000100110110111010100000101100010110010000101101000001111001000101011101110111000001111111111100010001010101111010010101001000110011010000000000001010111111101110111000010101011011111011111010111100110000000;
#1 $display("%b", po);
# 1  pi=207'b011100000111111111000101110010111111100111000111000011000000000100011011100101110111111011001100001100100111111001001110110111111100110000110000010000110011001101101101100101000101010110010011101111101110111;
#1 $display("%b", po);
# 1  pi=207'b011111010011101101100000100111011010001111011001110001101011000111010010001101010100011001100001010111111101001010101110001000000101000101000110000110111001000101110001011011000001111011001011100001001101011;
#1 $display("%b", po);
# 1  pi=207'b110101110001111110110010100110111011011010100100101101010110011011001011101000011000000111101010001110000011100101000001110001110110011100000111101111011111100110000101111000111010001100010101100001110100010;
#1 $display("%b", po);
# 1  pi=207'b110001101101100011011110111001010101111100101100001111001001001000111101100010000101011001100110001000011100111100011111010110001110000101001011000111010110100001010110001110001010010011100000001011001100000;
#1 $display("%b", po);
# 1  pi=207'b111101000101010000010011011010010010110110110101001110110100000001001011001101110111000010100010001001111000011010001011001100100001011100001110000111101001111000000001001110110100000101001100010100001000010;
#1 $display("%b", po);
# 1  pi=207'b100101110101001001011010110011001010010000100001001000111011011010100011111000010011001011100011010111010111010111010010111111110110000001101000111111010111001111000101100100100100000100000010101111111111110;
#1 $display("%b", po);
# 1  pi=207'b110110101001101110110111011101010110001110100010100111111011110101001000001100111011000001001001011111010000000001110001101000001110111111100100011000011110001011010001000011111100101001110001001101111001111;
#1 $display("%b", po);
# 1  pi=207'b110001110000011001100000111111001010110010000001000110010110011101100010110011000011010010101111011110111111001001111110101010110000011100010011100010010011011111111110001011101001110100010100010101011111111;
#1 $display("%b", po);
# 1  pi=207'b001111001001110101001001010111011010010011001001011010111111011100001010001110101000110101100110011011111101010100110101000011001011010101110101000010111111100010111010000010010001111010010001010000010010111;
#1 $display("%b", po);
# 1  pi=207'b010101100000000001100110010000000011101010011010101101100001000011110001111100001000010000010010011111110101000001010001011000000111101111000010111000110100001001001001001011100001010101001100100011111110111;
#1 $display("%b", po);
# 1  pi=207'b100111111111000010101111001000100011110100000010010010010011101110100000111111101001101110010100011000000000101100001110011011111101110100101000001010111101111010000111110110001110101001000110011001100010000;
#1 $display("%b", po);
# 1  pi=207'b001111111011111000110000000000111011001100011001001111100100010011111110111110100011100011000101000111010101111100100110100110010000101001011000101111101101110110000110101100101010101001001100110101111001011;
#1 $display("%b", po);
# 1  pi=207'b110010101000111101111111101100010011111101101010011000100100100010000010100101000111100100101100011110101111100111110111011111000010110011010010001010001111111011001000011011110001111001000010001111110101001;
#1 $display("%b", po);
# 1  pi=207'b110010100000000101000111101001011001000111111101111001011100110010101100011110101010100000101001001100010010011110111000010101000000000111110100111000000111010001110110010011001110100110011111000110001001000;
#1 $display("%b", po);
# 1  pi=207'b011000011010110010110011010010011101011101110111101111000110101011001011001110011001001100010001001000101110110101110111110001100100101000100011101011100111111110011010011111011011100100100101110100000100010;
#1 $display("%b", po);
# 1  pi=207'b011101101110101000010111001001111010100000001000011100111110000000101001011101010010111110101100110001101010101101000110111000010011110100000001100001000011101111010101011011011101001001100011000001000001111;
#1 $display("%b", po);
# 1  pi=207'b000011110100010011111011011111111110110000110010011011000100011101000001001001101001011101100110100100000111110111111000010011010011000100100011101011000111001101001111011011000010010100111011101100100100110;
#1 $display("%b", po);
# 1  pi=207'b011011110101000101100011000110000110001000011100111110000111011011100110001110010001000010110010110100100111000000010011111111100000110001011010010101101010000110110001000010110001111011001001110101111011101;
#1 $display("%b", po);
# 1  pi=207'b111111110001010010110101110001110010111110001111110111011010101100011010110111000000101111001100101111100111100000010101011000000001010001110010111111111011110100101011001011101101000111111001010010111011101;
#1 $display("%b", po);
# 1  pi=207'b001100101100001010100101010110000100011000001001111110000101110110101100011110110111001100000111000011111010110101111100100011000101111001011011001001111110100110010011011001010100111111001010111011101000010;
#1 $display("%b", po);
# 1  pi=207'b111001011010011000111111000000110111101111101010001100101100011101110000100100000100001110111111101110100101100001100011010001101110100111011001000010111110100101110001101011101100111000111011010011101101110;
#1 $display("%b", po);
# 1  pi=207'b111101111100101110101101110001100011000100010101001110100110000011011000000000010000111110111110011110010001100001110111100000101110010111110011001001100011001010101110010111010101001000000111001000110000110;
#1 $display("%b", po);
# 1  pi=207'b010001010010011011000101100111100011110010101010011100101000110001010111000110111001000000001011111010100010101010111100011110101010011010110110110011000010000010111000110011010011101111011000010000011000100;
#1 $display("%b", po);
# 1  pi=207'b000110011111101000100011100000101001111110101010111000110010100100001010001011101111100010001010110011011100000010100011100111101001110010100001110001100111001011111011100011111110110000111001001110100111000;
#1 $display("%b", po);
# 1  pi=207'b101100000001100111100000010111101000101001010100110100101001111111010100100110110100111101110000000100100100110001100001001010000010001000110100001100100110010110110000011101010001100111110110100111110001011;
#1 $display("%b", po);
# 1  pi=207'b101111001111010111011001010100000011111010000100111000110000000101010110000010001011100011001011010000110010111110000010001001110001110111101101100010111011000000100001011111001101010010000101101010101010000;
#1 $display("%b", po);
# 1  pi=207'b100001100000010011100001101100000101011010101011110101101010101010110011011010010000010110111000011101101101010110010110011001000101001000010001011001000011001111101101001100001110001100101101110110110110111;
#1 $display("%b", po);
# 1  pi=207'b101101011001100101000010010110010101011100011101100010100100000010001011110010100001001010100001010000110011100100000000101101100100100100000000010000101111010011111100100001001011101011011000010101111111101;
#1 $display("%b", po);
# 1  pi=207'b100100100000111010100111100100100101001010010101001111100001011010000100111110010011110000001010000111100100011110010101011000111100001100110110100001110101110110101101100011010111101010001100101100001011110;
#1 $display("%b", po);
# 1  pi=207'b010100110001000100100000100000001000001010111110011100101010011011000101011101011000100010010011101010001001001001101110001011010011010000101010010111001010111110001001001001011110110011011111100000111010111;
#1 $display("%b", po);
# 1  pi=207'b110011000101010010001010001101110010001011110001110110001010101110101110000011001010000111110010001101101100000011000110111000111011001110000000101111001101110111111001010011110100011100100011000111111111001;
#1 $display("%b", po);
# 1  pi=207'b111010010011011000100001000101110011001100011001000001001110101010000110110010000010010110111010000101010011000111100101110001111000111001100000111011010111000011001010010001000100010110010010101111010111010;
#1 $display("%b", po);
# 1  pi=207'b100000111010111101000001001101111111110001011110101001010001010001000110011011100011001101111011011100100010001101001110100011011000110001110010110011000100001110101000001010011101101100000100100101001001101;
#1 $display("%b", po);
# 1  pi=207'b100100101000110111010111110001010010110010110101111001011001110101000011010000010001110010100111010011111011100011000100101100000100000110111100100100110010101000001011010001111110000011001100100110101011011;
#1 $display("%b", po);
# 1  pi=207'b101100101001100000100010010100011001100000011001101100100001101100011001000111011111010001101100110100001100110000000110001100110001001100000011000000001011011010001000011010011111010000011011010111101010110;
#1 $display("%b", po);
# 1  pi=207'b011110101010000110001110000111010100100111111011110100110001111100011111100010100101110101001100111101100101101111100001000010110001001011101000110101000100000100010101000101110101001011110010000100001000111;
#1 $display("%b", po);
# 1  pi=207'b000101111101000110111101010010001111100111100101010111001111001001010101001100100010011010001100110100101110111101111000011000011101011110101101000101101100111110011110111110100110011101111000101101101011001;
#1 $display("%b", po);
# 1  pi=207'b111010001010111010110011100101000100001111110100111100111001001000101100110001111001010100011000011001011000001101011000101001001010100111111010111001100111110011010010001011101001011111111111100011000100000;
#1 $display("%b", po);
# 1  pi=207'b100010110011111010111100101110011101100010100111101010010010001111110110010010110111001111010100001001011110000111110011101000101110111000110111110110011101100100011001111100100111011101101110001000100101110;
#1 $display("%b", po);
# 1  pi=207'b101111011010101101011011001111000010010101000000000100101011100101101110011111001000010000100010110010110001111101111111110100110101000010000101010000111111001010001011110111001000100111110101110001110010000;
#1 $display("%b", po);
# 1  pi=207'b101100100011101111011110111110110100011100101011101111000011101011000001011100001010110011011110101110110101001000111010101111011011100001001101001001001101100000111010110111011101110011100111111110110001101;
#1 $display("%b", po);
# 1  pi=207'b110110111100111110101000101011011011110000000001001000010011000000111001000101101010110111010110101100110000001000010010011110001000010110110111000010011100011110101001100000110110100010111100111001111110111;
#1 $display("%b", po);
# 1  pi=207'b101111110001010101001100000100100010101011101110011100100100111000110100011101101011001011100000110110010011111010110100010101110110010000111001111011101110110111100011110101010100000110111110110101101100100;
#1 $display("%b", po);
# 1  pi=207'b000001010010000111000000111100010010001000010000010111011111011001010110011001001010110111100111100000101010000010101010010010011100011101011011011100110001001111110101111010000100110011110111110100001110100;
#1 $display("%b", po);
# 1  pi=207'b011110010110101010001000010010001011110111110111101110000111001110100100101100010010101001001000001111011010001010001100100110101010110100001000100100010010000001101110001010011110101011101101011111110101101;
#1 $display("%b", po);
# 1  pi=207'b100100110111010000001110101001110110111010100111000101110011111011111100010110001100110100000010001010001011100110011100011001111101101111001100011011111010000011111011011110100111101100110110101000111111010;
#1 $display("%b", po);
# 1  pi=207'b110011100101011100101011100001001111001101001100010111100100000110001000000010101100101111111001110011101010110001001011010111011010001101110111100101100100011101011011001100010111010010000111000110110011111;
#1 $display("%b", po);
# 1  pi=207'b101011110110000011101101111001111000001011111010110010010101011110100011100101000001011111000000101111000011000001000010110101110110010011101101110100111100001010000000010100001110100010011010110101101011101;
#1 $display("%b", po);
# 1  pi=207'b100111100010111101101011011111010101111000010110010111010001001010011011101000101010110100010001011111110000110111101000010101011111100001011011110011011001011101000100101101011000111010010001001111101001010;
#1 $display("%b", po);
# 1  pi=207'b001101111011000000010010101000010100001110111011000110111010101101100100101111010011101101000111100111001101001101100101000111101010110011100001100001101101001100101100110100100111001110101011010011001111000;
#1 $display("%b", po);
# 1  pi=207'b010101001010011001000100110000001101111010001000011001110010000110101001011110001101000010001100001001010000000010101110110100001011010000000001011011010111110110001001101011011101100100000010010011011011111;
#1 $display("%b", po);
# 1  pi=207'b101100000000011111001011000110010110111100001100111111001101000110011100100000100101111000001010010001000100110110101101011011010111000010011111010101001001001000011000010010110100110010000011000100100010110;
#1 $display("%b", po);
# 1  pi=207'b011010000101000001000000010111100010000101111011000000001101011001011000101011001011001100010101100110010011000111011111001111101001111101110011110001110001110100001101010000100101111101110101000000010000110;
#1 $display("%b", po);
# 1  pi=207'b100000000101001111000000000001001110011100001111101110010010110000101001100001101100011111101111100101111100011010000001100011101111110110010010101001010011111010011101011001000110101101000000110111001111011;
#1 $display("%b", po);
# 1  pi=207'b110000111001111101101000000111111011010010110011001100001010011111100000101010100000001000011000000100000100100101101011111100111100100110010010110000100100000000100000111101011011001001111001010011101111101;
#1 $display("%b", po);
# 1  pi=207'b100101100111000110010111111100100100010001001000011100011000101001100011100010100010000110000110010111001011011111100111101110000010100000001001111111111010010101100100001000011111011011101000111110111000110;
#1 $display("%b", po);
# 1  pi=207'b001101001011011110101100101010010000110011100011010110110000010101100000101110111111010001100111110001011101000110000011011000010001010110111100101111000010011010011010000010101011000000110010110010100011110;
#1 $display("%b", po);
# 1  pi=207'b001001110111011101011111010100110000010001000100111110010100101000011010101001110111010000100101100100000000001000001000110111111000110001011011110000001100101100101011010110011101101000001000011101101010010;
#1 $display("%b", po);
# 1  pi=207'b100001011110001011000011000011001111011000010010100111000010010110011001100011101110001010100101001011011101111111010100010011101001101001010110100001100001101010110111010001110111010110111000011000001101111;
#1 $display("%b", po);
# 1  pi=207'b000101110111010010100010111010011001111110111011001010000110100100000001011011011000011011010110010101000101000001110011111010101110101010110101011111000010001101000111111010010001111011011111111010101010110;
#1 $display("%b", po);
# 1  pi=207'b001110010100111001001100101110001100011000100111111111111011001101110100101000011000111111100001011111001110110011100000100000001101010100010010000101110000011101001000011010011001000101100111001101101111101;
#1 $display("%b", po);
# 1  pi=207'b100101000110101001001000111100000110001011000000110110111100100100100110011100011110110000101111000101101001111100110111110010000010111100011111111110101011100011001010111001100001001001100100101101101100101;
#1 $display("%b", po);
# 1  pi=207'b100000001101001111101000110001011010000100001000111110100111101101000001111001011000011000001111010000010011100001011101001000010011101001001111010100111001110110010100000101111100110000000111110000010111011;
#1 $display("%b", po);
# 1  pi=207'b001011011101010001100101100001100011110100110111111100001110000110101101100001110000101111011010111111010010100011000111100101010111001110010100001001010100000011100100111000011101110001001011101110101110101;
#1 $display("%b", po);
# 1  pi=207'b011010101011111011110110011110001011001111010101001010010010110011101011000111100010010111000010100110011101111000010011101010111101000110011100010001111000110001111001111111111010000100111100001000101100001;
#1 $display("%b", po);
# 1  pi=207'b010011110101001010000001100001010000100000011100001111111100101010101111111010110101011110111000011111010011101110000001110110001011101001111011101110110111011010000101011111000010000110011001111100100011100;
#1 $display("%b", po);
# 1  pi=207'b111110101111101111010101101010110001100110101101111101011000001110100011011010000010011011000011001011111010111110010000100010000100101100010111001100011000100000001010101011011010101111111101011011100111000;
#1 $display("%b", po);
# 1  pi=207'b100101011100100100110010111111011010011111011001010111110001001001111111110101010110011000000100101001110000110010110010101111100000101111100110011101010100000111110100011111100011100011110110111001000011001;
#1 $display("%b", po);
# 1  pi=207'b000000111011111111001100010111110010111000101000110111010010101001011100011111101010101010010000011010110010001011011101011011100110111111000001100100101010110101000101011100110101010000111110000010000100110;
#1 $display("%b", po);
# 1  pi=207'b101011100010100101111001000100010111101001001010001111011011101001100011101010101101110110010001100111111001010110000000111001000010000101101110110101101011011100001000001110010010111101000101010100100001011;
#1 $display("%b", po);
# 1  pi=207'b111101001101011011001011000001011010011010011010100011000110011001001011110100101111010111000111001101010101011001011010110101101101111011101100100001001110000101001010000100000111101000000001101000001111011;
#1 $display("%b", po);
# 1  pi=207'b010110110111010110100101101111100111101000011101101010010010001111110111000001100011110110001111011000111001110001101011010111010010010111011110110010100010101101110001100100011101111100111101001111000000011;
#1 $display("%b", po);
# 1  pi=207'b110101001000100011001110000110110010000000010111011101110100100111100111010101000110000101111101111100101000110110010101111011110100011110000001011010001100111011101111001100100101000100100000011000001110111;
#1 $display("%b", po);
# 1  pi=207'b011011010110101010110001111011010111100011000010110100001001000000101011011101101011010111001100111100011101011001111111111010010010011110000001000110100111010111111011110100010110110010001001101010000101011;
#1 $display("%b", po);
# 1  pi=207'b101111001011110101111011110100110101001111000101010010111011001100100011110000101111001000110001010101110101100100101101010110100110011101101000011100100110001000000100111110001101010110000111100101110000010;
#1 $display("%b", po);
# 1  pi=207'b010010000101001001001110000110011111011101011010100101001001101101000010101111001100110111001111100110010011111110110100010100011111000100110000011111110000011001011100010100101000001010000100001011111001111;
#1 $display("%b", po);
# 1  pi=207'b011011111010110100001111100110011001000011001111111111111001011100101000110100001010111100011001110001110010111110010110100110010100001100011000011001101101111110001011111011101011101110001100111110100110010;
#1 $display("%b", po);
# 1  pi=207'b011110010111100010010111101001111001010000001011100011011111001001010101000011010110011111000111010011110110110010000000010101101100101111001110111100111000101110011000111100110111110100011000100001011010010;
#1 $display("%b", po);
# 1  pi=207'b110110110101110000101101101101100011111110000010011100000000111010110010111100101011111101011101110010101101110101010000011000000111010110100100010100010111111001000001010101100101010010011100001110100101110;
#1 $display("%b", po);
# 1  pi=207'b110011111111101110010101000101000111100111111011010001110000000001011110101010001110011100101100101110111001001001110010011011101110100111000101000101111011011000010111110011110010011110011110011011101110100;
#1 $display("%b", po);
# 1  pi=207'b100010001111001010000100001100101001001111001111001001001101011000011110011010001110101011000111101110110111110000100101111101000101100110000100101100000010110010100110111010000111110110001100010000011000000;
#1 $display("%b", po);
# 1  pi=207'b010110010101010011111000001001110111110101101001111011111010100011111010000011010111111001101100000010000010101000001001010110011011011111101011101001110110110011101100000011001111001010000110110111011001110;
#1 $display("%b", po);
# 1  pi=207'b101111110010010110111010100010000010101110110100010000110000000111011001100010100001100110010011100010101010010101111010100101011011000000011100101011000100111001010100001001101101111101100010001111001010000;
#1 $display("%b", po);
# 1  pi=207'b101011111101101101011000011001100101010000110001001110011110101100000110011101110101000101001010000010101111000110101111110000111111000000010110110100101100100100010101000111010100111110111100111011000100100;
#1 $display("%b", po);
# 1  pi=207'b000110101101100000101100001111011110110101001111001011010011110000111111111010111100011111101011011000001011000011011111101110001010110001110010011100100001111101101011111001000001101000100001000100100000011;
#1 $display("%b", po);
# 1  pi=207'b001110101010001110101100010111011111010000111001101011101111110001111011000111111101111101110001111011000101011010100111101111111010110001101001000010001101011000110000110000001100110101101000011100100100011;
#1 $display("%b", po);
# 1  pi=207'b111000011110110110100110001000111000000100010011110111000111011000111010010100001011010011011000101001000001010001100011010001101010101011001001110100111111111010100110111010101011111111010101001110100111001;
#1 $display("%b", po);
# 1  pi=207'b001001101111110011001100111001100111010000100011010111011010001101000110001100100100010001101101111000011010101111101000011111011010011001111110101101001000011101011011000111101011001011100010100011011011100;
#1 $display("%b", po);
# 1  pi=207'b010011100001100110101001000010010001000111011001001011110101110001000111111100010001000000101011101110100110110011010010101010011101111100001110100111001111001001110010111110001101101100000010100101101011011;
#1 $display("%b", po);
# 1  pi=207'b111100000011001010011011110111101111101100011111110101010011010101100000111000111000000011101001001011110000000000110111110011010100111101000110000000101110011001100000100110011111000100011100000111101110101;
#1 $display("%b", po);
# 1  pi=207'b110101010111011010111010100101010111100100111101010110000001000111110110011100100001010010110100000110011010100010010010111001001001110101001110010111111101000001111010111111001101011000110011101010010011000;
#1 $display("%b", po);
# 1  pi=207'b100010011001000001001000101110110101100110011111110111000010011101100100111011010101111100000111110111000000011100111000110111110101101100000101010001111000100001011000110100010011011010000111000111001110001;
#1 $display("%b", po);
# 1  pi=207'b001001110110010101110111111110101000100010110100000001010010111010111101001100010001100010010100010111010111110011010010101111000100100101100111100100101011100111001111101111101011001100000101010111111000110;
#1 $display("%b", po);
# 1  pi=207'b110110100010101001111001111010100110010011001101110111111011101011110001001100110001101110110010101001100110110110111001000100001000101001000001101010000010010010000010100111111110100001010001100011111111000;
#1 $display("%b", po);
# 1  pi=207'b000001010111110010011001000100110010010100010101001000010100100101011001101010101111101100110101011011110001011000001000110000011001000001111000000010011010000101111111000111001010110101110010110000011101110;
#1 $display("%b", po);
# 1  pi=207'b110110000001010010110101100110101011101100101011011001111110011101010011001000001000010010010000001111000100100001101010111100001101001110010011100110000111000010100001111110011001011101000001001010001000100;
#1 $display("%b", po);
# 1  pi=207'b010001100001100000101100010010101010111010110000001010001101000011101100000000110101011010110011001010010101011001010000011111011111100110110011000001110111111110001101100001000011011110110100110001100111010;
#1 $display("%b", po);
# 1  pi=207'b100010001011100111001001111000111001101011100100000000110100011001000000011111111010010110000010011011110001011000001000000111110000101010011011001110001111011110101100001110000000100111010100010001011110101;
#1 $display("%b", po);
# 1  pi=207'b011010010111101101011101100001111001100011001110101111010010000000110101101010111100101111110111000001000010001011110111001100110001001001110111011100000001110001100101010001001111111100001110110000100010011;
#1 $display("%b", po);
# 1  pi=207'b010000011011100000000001111111011101100010110011100001111011100101000110001100101100010101111010010100110001100110000001011001001011000110101010001110101101000110011101010001100011100111000101100101101111101;
#1 $display("%b", po);
# 1  pi=207'b101101110001110111000101100000001111011100011010111010011101110101110111011001011011011101100011111111110001001110111101110101111001110100010110011001100000001010101010000110010011010110110100011110100000111;
#1 $display("%b", po);
# 1  pi=207'b101011100100001001011000100100111001011111111100000100100111011001001101000011110101001000000110011010010100010011100110110001000000010011101101001101001000101100010001101000010111111011000111100001010010001;
#1 $display("%b", po);
# 1  pi=207'b011111100111101110110100100101011100111110001100100011100001111011011101111100100111111101001111111000100011111000100010000011111001111001011101000101010101110010000101011110111111101001100100100111000001011;
#1 $display("%b", po);
# 1  pi=207'b000001011110010010110111001111011111110101010110001000001101111111010100100001011110001100010101000111000011110010111110000010110010101100011100110011001100101010101100011101000111011101100010011110000101100;
#1 $display("%b", po);
# 1  pi=207'b101010001101110000001000010101000100111011110001011100100110011001110001101000101100100010001110001111101011001110100001110011101101000110011001100111010010010100011000110111100111011111100000010001011001001;
#1 $display("%b", po);
# 1  pi=207'b101001110111010001100000110111111101011111001000110010000011100111010010010101001101100111110000101010001010000101111101011111000001011001001100100110011010001101101101011001111011000111010000011111011110101;
#1 $display("%b", po);
# 1  pi=207'b111100001110000101010100100111101110000000011011100011011110000001101001011000001011011001010101001110010111000011001110111111110111110110101001111011001001010011001101110100101110110000101110111111000111000;
#1 $display("%b", po);
# 1  pi=207'b001001111110100011101000000111011100100100100111001111011000001101001110110001111110001101000110101011101011110001011011000111110111010001101010011111011110110010000101100001001010010100110111110101001110011;
#1 $display("%b", po);
# 1  pi=207'b100101011111000011101100101001101100001110100111001100010010100111001101101010111011101101011101011010101110110010100101000110100000100101101011001111110111011111101111100010011010111110011000100011000100001;
#1 $display("%b", po);
# 1  pi=207'b100010101010100110110100001000111001001111110011110111001010001001100100100000110000111011111010010110101001100011011111010100011100101110111000010100100000011110100001001110011100000100011010001111000101110;
#1 $display("%b", po);
# 1  pi=207'b110101000101110101101110010000110101101010101001111110010001100100101101011000001110110110111101101101000001101011001010110110101100001011011000100111100101001000000010110101111010100100001000010010110010001;
#1 $display("%b", po);
# 1  pi=207'b101111101101101010110110110010010000100111110101001101001000010000000111001011000101110011011111110100000010001010110110110011100101001111100101100111010000011001011100011001111010000011111000011110110101111;
#1 $display("%b", po);
# 1  pi=207'b010011010111011011100000111100100011011110111011100100101000110101100000011101100011011010101100001010001001001001101000001011100110111000111000111010100110000100101001001110011111101001010001101001110110111;
#1 $display("%b", po);
# 1  pi=207'b000111110011011111001011110011011010001110001000000100111000111001001000000101100111100100001001010001000110001011100011001010101011100100001110001010101100110101011111101100001011100110001001101010011111101;
#1 $display("%b", po);
# 1  pi=207'b100110011000010111011110010011011010101101010010101100010000000000001001011101100100101100010100001001011000110001001101100110001000000111000000110110000111100100010110111101110101010000111011110101111010111;
#1 $display("%b", po);
# 1  pi=207'b011110110111010111011011001111101110100110000110101110111111000001110100101011010010111010011011010010100100110101001011110001010101010110100100001110011010101111000010011010000001000010001010001010011001101;
#1 $display("%b", po);
# 1  pi=207'b111010110101100010101101111101001000110101001010000011101000100011110111100110001110100011110111010001101100000110101110011000011010000111111001101101001101101011100010010000110101001111010011111111101011100;
#1 $display("%b", po);
# 1  pi=207'b000000000111100000110111000000001001100010000000111100001000110001111110111100101010001110101111000010001111100000000111010110110101111010001110000000011100101001111011010000100100101001010000110110010100010;
#1 $display("%b", po);
# 1  pi=207'b110001001010101100100000010011000001001001011110010000010001111110101110000110110111111010100110110000001100110111110110100110111101000111000011111001111001111111110110011110101010110110100001100000101011010;
#1 $display("%b", po);
# 1  pi=207'b110101110000000101101110111111000110000111110111001011110101010000101111100100010111001001001101000111001111001010011001011101111101010110101111111111010101000010111010110100010100011101100010101111110110110;
#1 $display("%b", po);
# 1  pi=207'b100111010000001001010000111110010100110000010101000000111100001000111001011101110100111101001100000110011000011111000011111100111011010011011101000110011110111101111111010100010001010110010011100100111000000;
#1 $display("%b", po);
# 1  pi=207'b111000100100110010010001011101011010011100111100010101100110000111000101101100100111100101111101111001101101100101110010000010101000101010010111000100111001111110011010100101010111100101110011011010010000001;
#1 $display("%b", po);
# 1  pi=207'b100101110001111111111000001100000110001110010101101101111110001010000101011011011011100000101001110001101010001001011101011100110101101001000011100100010000111111010101100010100111100000100100111100101000001;
#1 $display("%b", po);
# 1  pi=207'b110010100111011011011011101101010111110011000111111100001001100011010101111011100000100010101101110111000011000101110010110110001001000010111101110100101010010001101001100110110010101101100100010010001011001;
#1 $display("%b", po);
# 1  pi=207'b110011100110011100011000100000011101100100101011100101110111100101101100001010100100011001101110110001010111000110001010111111011011010010010011000101111011010111100010111111110100010000100000110000110001001;
#1 $display("%b", po);
# 1  pi=207'b010111001000011010011000010110010101101000111001000101111000001000110110100100011101010110010101101010011011010011101011011000100000010110100001011101101010101101111111000011110010101010010110010110010101111;
#1 $display("%b", po);
# 1  pi=207'b011001001100011111000101010100110100101110000101110110101101001010110100010100010010111110101000001101001101100110101011000010000101010001001110010000010101001010111110001001010011110000011111011100110001100;
#1 $display("%b", po);
# 1  pi=207'b101111010000011001111010111011010011001001000101001100101110101101011110010111100010011010111000100100100010011100001000100010000100011000011101010010010001000100110001010110011011100111001101110100110101011;
#1 $display("%b", po);
# 1  pi=207'b001001010101011011101001110100000111111110110100100111100010001010100000010001010111001001101100001001001111110001011101111001111000010011101010111001000001100100100010111101101011011000110110000010111111011;
#1 $display("%b", po);
# 1  pi=207'b001001110110000101011001111001101011111110011010111000110110110111100110100111110000001101010110011010010001111101100111001001111001110011100100100000100111101000110010110101110111100000111000010010001010101;
#1 $display("%b", po);
# 1  pi=207'b100010110010001100001101010101010001100111111001100111000101011111101101000011111001001001000110111010011011000011001111101001001011100101110101011001000001100111001100110011011100111100011111110000010010101;
#1 $display("%b", po);
# 1  pi=207'b101110001101010011001000111110000010010100011100111110101010110011001111100110011100110110001000001001000010010110111110110111111011010011011110100011011100011001001100011101010100100101001001010011010101111;
#1 $display("%b", po);
# 1  pi=207'b100011000011010011001000111001100100011111100010100101111101111100011010010101101001110010111110011001101000010001001111101001000001000110000001110100101000000101111111010010001111101100110010000000011100111;
#1 $display("%b", po);
# 1  pi=207'b001111111001001110110001100011110010110111010000100101000010111000001000100010010110111100001110000110100010111101001001111110101100110111110011001000110111010100101001010001111101111110100110111100100101111;
#1 $display("%b", po);
# 1  pi=207'b111100111101101011010100011111100111010110101101111011111001011110010111100001011111111011100000111010111010010010101101010111110010010000110010111111100101001100000110100110101010100111010110111111010100100;
#1 $display("%b", po);
# 1  pi=207'b101000100010011011111010001001100010001100001111001010100111100110110010010101001110000001101000100110111010011100110100001111010001100100010011100111100011111100001100001111100011101111010000110011101111001;
#1 $display("%b", po);
# 1  pi=207'b000000011011001110011100101111001011110000001001010101100000010101101100111101010101101011011010100101110001011100001010110110100001000100001101000111010110001011000100011111011111010001001101010001000000100;
#1 $display("%b", po);
# 1  pi=207'b001100100111100000001111001001101000111110010111101000100000011111111000011000001111110101011110101100010110111100000011101101111101100111100010100011001011110000100001010101001000101000111000110011010101010;
#1 $display("%b", po);
# 1  pi=207'b100001110011101011100001001110101011100111010111110100000111000001110110110011111000110110110001011010011111111110100001011011101010000111100110010100101011100110000111001010101101100110101101101111111111010;
#1 $display("%b", po);
# 1  pi=207'b100101100011010111010100100101010110110010110000011100000010101011110111000000001101011010010100101110100100000111111001010010011010101100101000100111111010110100011111011011001000011100010110110011010100101;
#1 $display("%b", po);
# 1  pi=207'b110100010110000010000001110110111010111101000010101000010011001010000000111011111011110110011111101101000010111011010001001011110100100101111001111101000101111101100011111001111101000110001010000001000000101;
#1 $display("%b", po);
# 1  pi=207'b101001001000010111001110010001011100111011010111111010000111111101011110101010111000110110000011101011101101110111001111001001110001010100110111011011110010101000010100100100010101101101100000010111011111010;
#1 $display("%b", po);
# 1  pi=207'b000001010111011011011101100100101111101010110011001111100010101110100101110000000101000111101110110111111110100110000000010010010111001100110110000001010010110100000100110111001100111000110101101110111100100;
#1 $display("%b", po);
# 1  pi=207'b110011100110011010100000110011011000001100110000101100011100010010010000001001011100000110010001001001111101001010110000100001101100110110111000010101110110101111101110111000101000101110010111000101110111100;
#1 $display("%b", po);
# 1  pi=207'b110111110010010011011010001011100001100010110111000010100010001101001101011100001111101010011110000010101110110101000010010001100110101010111111101101010000001110101001110011011101100101011110011000100010111;
#1 $display("%b", po);
# 1  pi=207'b110010100100101011011110101000111110100011111001001010011110111100100010101110111110000101010001110101101110001101111100110001011000010001001001101100011111100011001100110110011111101010110001000111111011010;
#1 $display("%b", po);
# 1  pi=207'b110001001101110101010000101001011110000101110111001110110000011011010111110101111010000100001111010001011110011011100000000010100100100010000101111010011111001100111011011000001100101101111010011000000010111;
#1 $display("%b", po);
# 1  pi=207'b001100100110010010011100000100101011010110011111111100100011111011111110100010010111010011001110100011011110110011100101100111110001100000111111101010000000111101000111001010101100010011001100100001111110111;
#1 $display("%b", po);
# 1  pi=207'b100100110011011010011010100110011010000001101101010000010111011011100110010111100000101111010100101110001111111111101010100110100011001010100100011101000000101011011000101100000010010111000110101011011110011;
#1 $display("%b", po);
# 1  pi=207'b101011000101110011100101000011001100111100011100111000100101111000111011101011111100011101001010101110100100010001011100011100001110010001000110110010100000010110010101110000101101111100101011001010010101001;
#1 $display("%b", po);
# 1  pi=207'b111110001000101100110001011000011010100010110100011100011101100110101110100000110000110111111110101111101001101011100111011001101000010100010111101001101111101100010100111000010110011011000110101101101000000;
#1 $display("%b", po);
# 1  pi=207'b000110101011100101111010110010110110000100100110001100011001101111010010010010110111110010110110110011110001100101001011101111001100111111000111011001110011100101010010001010001010101001111101100101010011101;
#1 $display("%b", po);
# 1  pi=207'b011101000011010011011011001011011000110110001010000001011010110010011101110110001110101111100010110101110001110000000001101100101000010000000101001100010111010010111001001111011111110010010100110011011010110;
#1 $display("%b", po);
# 1  pi=207'b111011001110111110001111111110101111100000100110001100001011111110011101011010011010000010111111010111001000111010111010111110111111010110010111011111111010010110000111111100101000110000101001011001011110101;
#1 $display("%b", po);
# 1  pi=207'b111010011011000000011100111111011010001111100101001100010101101101010111000011101101111100011101101000011110100000110001011010100101111101001011110111010010100010101011001101000000110100010011110010010010110;
#1 $display("%b", po);
# 1  pi=207'b111011001000010110000110010010100000110011000100010001000001010011100000110100101110000110101101000111000100011011110010100001011111111101101000100001000110110001011111100101111101110111011010110110100001000;
#1 $display("%b", po);
# 1  pi=207'b011010011000100010100110111111101001101010010001110100111000100111111100010001110111111110011010000001001100101101110101111101000001000011110110110100010000100110010000101111000111011011100110101011010110111;
#1 $display("%b", po);
# 1  pi=207'b111110111001100111010101101110101010010011110111000001111111011001010101100101100101001011110101100010101010110100100100001001110011110010011010100101010011000111101101111110010110111111111111001001001001001;
#1 $display("%b", po);
# 1  pi=207'b010010100011000001101010100010101010010111101010100010101000010010001010001001100001011101010100011001000111000110011011111000101011110010111111010001101000011110101011111011100111101111011010101000111011011;
#1 $display("%b", po);
# 1  pi=207'b000001001110000011101111111111011011001111111110101110010000101111011110100101100001011000101111111000111101101110101001000110111110110111001111011101111011110010011110011000111100111010100111010000000111000;
#1 $display("%b", po);
# 1  pi=207'b110010011101100100000011110011001101101000000010111110111011100100010101111100111111101110011001110111100101001000001111110111000011100000111010011111001000010011010001011101110100001011101101000001001111010;
#1 $display("%b", po);
# 1  pi=207'b010110111110101000001100001001001110001100101110100100100000101100100100001000111111001011100001101100100000101101010100101001011110101001010011110110000111010001001010010111011001011000110010100100011101111;
#1 $display("%b", po);
# 1  pi=207'b111110111110001001000100100111000011100000101011011010001010111100001110100000011010010010010000001011011101011101101000000101100011100100001110111010111011111011010000100111111000110110110011010101100000101;
#1 $display("%b", po);
# 1  pi=207'b011010110111011110100111110101100110000001011001111000011100001111110100010110110100011110101000000010010101010111000100111110101111111100010100101100000111001011000000010100011001111100100000100011110010011;
#1 $display("%b", po);
# 1  pi=207'b000100101100001110101101110011111111110000001101111111010110010001100000111101101110010001101100101100101011100110000001001000101010101000111000110111111101110100000100100111000110010011110110011100000110010;
#1 $display("%b", po);
# 1  pi=207'b111010011100011101101111010001000001011010100010100010000010100010101001101101110110001101010111001111111110010010100010000111110001000010001111011000110111001110010011001101101000110000010101111000110001101;
#1 $display("%b", po);
# 1  pi=207'b000001011111100100111100011010110111011001001001000001001001110000111100101111101010000100110001000100011010001010100111001111100001110101010111110000011011111110000110111110100010111100101111101100111001001;
#1 $display("%b", po);
# 1  pi=207'b110100001011010111000110011101001110100101001001110111101111010110100011110110100011010110110011011011000100111011111100100110001011111110110110000010000010111111001000101000010100101100001001010010011110111;
#1 $display("%b", po);
# 1  pi=207'b111111101000011001001110001001001110101001000011110001101011001011110011000110101110011000110111010000101111011010000011110010001110011111111101101110000101001011011110001000111001010101111011001111001001011;
#1 $display("%b", po);
# 1  pi=207'b101111000010011010101110110011100011001100000101101101001100010000100100110110001110101000000110101000101100100101010100101100001001011010111000010011110110001011100010000111100011110110000101110111111001011;
#1 $display("%b", po);
# 1  pi=207'b010110111111010100101001000101111100111001110101111111100101000001111011000011010001101100100111111010001100010101001101001110011101010101001010010010100111100111100011000010010011001010101000011111010101010;
#1 $display("%b", po);
# 1  pi=207'b110111100100001001011100001111110110111110110010000110011010111101010101011100110111000000111001110010000111100100000000000011000000000111111110111110001101011011111001010101011111010110010001110111000111101;
#1 $display("%b", po);
# 1  pi=207'b000110011010111010100010101101011011101111000100000010000111001010101111010000111111111110111000111001001000101011001111000011000000011100110100011011111101010011001101111110011001101101010110101111000010011;
#1 $display("%b", po);
# 1  pi=207'b001101101101011100000001101100000000101110100011000001000000101111100101010101110000110011111110001110011100000110010011000000101100101010101101101100000001110011001101100010001000000001111001001010110011110;
#1 $display("%b", po);
# 1  pi=207'b111000101000000110111110000100011101101011100011010001110110111111101010010010100111111000100110110001000100110100101110111011110000110111110011111010010011010010101101101111011110101101110010100111111010100;
#1 $display("%b", po);
# 1  pi=207'b100011011101110101111000011100110100000011111101111001110111111001110101001110000111100000101000011010111110010000000001011101101001101111010111000000110011110001010011101001010111001100110011001101000010000;
#1 $display("%b", po);
# 1  pi=207'b000101001010011011111011110010000101010000111001101000101101111001100101011110111011011101000011000101111111101100111001101111010010101000010000100111101001011100011000010100010000101000101111010111001110111;
#1 $display("%b", po);
# 1  pi=207'b011101010101000100001011001101100001110010110111001011111111010010000011101010100000000011001010111001100110100001001100100011101000000111100110100011000010011110000000111001000011111011000010110111000111101;
#1 $display("%b", po);
# 1  pi=207'b011001101110100110100111100100000000111010011000010110000010011001111111111010000000010010110000001111001001000100111011111110100110000000101110001011101010001011010101010111000010110000100110010111101001111;
#1 $display("%b", po);
# 1  pi=207'b001010000101111100101011111001010010010101010100101110101001001010110111111101001000101110010011111010011100101001001011111110001000111010011101111101101000010111110011111000010101010010110000000101011011011;
#1 $display("%b", po);
# 1  pi=207'b110000110110110000001011010100110001100001000011000101110100101111011100011100010100101101101100111010110100011000101001011010101001011110011000011000100100111111100100101111001010000010011110100101011100101;
#1 $display("%b", po);
# 1  pi=207'b100000010110100001010110011101101111001111111100001101010010001011111101100011011101010010010101110100000110101101110100010110001111110100101000011100111111101001001110011111010001011111010111101111111011000;
#1 $display("%b", po);
# 1  pi=207'b110110100101111100100001111001110010011101101111111001011100100001001101101110000101010101101010010101110111101111001111100101001011000000111010110101010011001110111110110100011000011111001011011011001011111;
#1 $display("%b", po);
# 1  pi=207'b011110011110000010001011001001001110000010100010111110111101101001010010101101100100000100010110101010010010011000100110110101001000110001000010101111110110000010001110010101010001110000000011111010001010011;
#1 $display("%b", po);
# 1  pi=207'b100110010101110001101010100010011100010010101101011100010011110010010100101100010101111111100011011010001001000110010011001100110010010110001010000000000110110001100100011111110111111110000011000010000101011;
#1 $display("%b", po);
# 1  pi=207'b100110000110100011011001001010001000111111101100010101110001001010011100000101001001000101000111010101100101011011100100000111010001000111000101010111101011010100100000101110100010000001001110110011010011010;
#1 $display("%b", po);
# 1  pi=207'b100110101101010100101110100001010100000101100111010100100111100001101000010011100110110110000111111110010001011100000101110010001000101111011011111000101010010001000100001011010100110001010111010101001100111;
#1 $display("%b", po);
# 1  pi=207'b110111110000011011101110111000001011010100001000010101000011111000010001001101101010100100010110100101000000001011010010111111000010101111101100110010101100111000011010101000011001100110100101010110010011011;
#1 $display("%b", po);
# 1  pi=207'b011001111110111100110010000110111000001100011100110010001011101101110000101101111000101101101110010110100000001010010110101101100000111001110010001000101101110110010001000010011110001000100001110011001010111;
#1 $display("%b", po);
# 1  pi=207'b111111101010100100000100000101010011111110001011000001100101101100010101110100100101110000010100101000011000100000001100111100101010100011010011111111111000110011111000110010001010110010101110111101101111000;
#1 $display("%b", po);
# 1  pi=207'b000010111001000000110111010011101111110010101110100101101010101000011100011101101011101010000100101110010110110010000000100011001011101111001111110101100011110010101101000011111010110010110011011101001110111;
#1 $display("%b", po);
# 1  pi=207'b001110111111000101101111100101001100010111110010011110101111100010100010000010000110111000011010111111011100001111010111000101100100010000100111001010100101101101110100001111011000110100000001100010111000000;
#1 $display("%b", po);
# 1  pi=207'b001011010100001111001100000001110010001010100001011000111101111101110111001101010001001001110100100010110011101110011110101111100110000111011111101001001011110100111111111001010000101011010110000010011011111;
#1 $display("%b", po);
# 1  pi=207'b010100101000111111100101100111011011110111101101101101111111001101010001011010011111001011111010101111001111000111011000100101100000100011001010010101110110111010100100100000101110010000010110100100000000110;
#1 $display("%b", po);
# 1  pi=207'b011111001111010101000110111101001001010110100111111100110101000100000000111001000010110010000010101101100111011110010000100001101110100000100001000011011011101100010100110010101000111010001110010010010101011;
#1 $display("%b", po);
# 1  pi=207'b111101000101011011101100000110001111111110100111010100000101000101000000111101001011100101110101011100011101000000011111111011010000100110100011101110011001010001100110100000011101101010101001011010100000111;
#1 $display("%b", po);
# 1  pi=207'b110110111110000100100101110111011001001110101010111100101001001011010011010110011010101101010111110111011100011100110001011000010111100011001101110111001111101010011111111001111001000101010101010011001011000;
#1 $display("%b", po);
# 1  pi=207'b100010110010111101000110110001101101110000011010111000011100001011010111011100110101010101111010001010011011000000000101111101010010100010101101111101101101100001001011100011100001101010111011010110110100011;
#1 $display("%b", po);
# 1  pi=207'b011101111010000000100111001111011011001011111001001111011011000001101110110001100001101110110010111101001011110111001011100000011110110100110101010011101111011111100010100110100111000101011110100010001110111;
#1 $display("%b", po);
# 1  pi=207'b101111010101010110101101110110001101011010000110011111011110101010010010001101110101100011011100111111111111110101111110000011110111001000000111011010110001001111000100010111010101000101010101111000100111001;
#1 $display("%b", po);
# 1  pi=207'b011001110101000000010100000111010000111000111100000110111001110001110000111100101010111011100011101000001000011101100101001000011100010011111001011101111011100011110110010000000110001010010110011001000111010;
#1 $display("%b", po);
# 1  pi=207'b111110011001001100100000001100101000110010110001001101010011100101010001001100100001000000101111011011001010001001110000101100001011001001000011111000000000001010110001000011110101001001010110000011011000000;
#1 $display("%b", po);
# 1  pi=207'b011000000010011100110101010010100100110111111011101111100101101101000000111010011110110001000101110001100110011010101101111000101000000100001101000110100110111011010011011110010010100110111011001101010111001;
#1 $display("%b", po);
# 1  pi=207'b011100100010000010001110000110110000011100110100010110100011010000111110001110110111010110111010011001101111101010010000011011101010100100011100111001001110100001111000101000001110000110010001100010011010111;
#1 $display("%b", po);
# 1  pi=207'b010100111111000100111101011001010110110001110011011011111001100100001100001100011111000101101100000110011111001110110010000111101101101110110101011010101000001100110011100101111100001101010110110110001101001;
#1 $display("%b", po);
# 1  pi=207'b111000111000110110011111001111000011000100111100011010111100011110101011111110111000110010011111110100001001100100010100100001011101111001001001010000001000001111001010000011000101010111101111000011110111110;
#1 $display("%b", po);
# 1  pi=207'b111001010110111110010010010000010111110011110101011011101100111000010110010010011010001110001111101000001000000011001101111100001110001011110010100111111001110010100000100111101100100101011010111011110101101;
#1 $display("%b", po);
# 1  pi=207'b011110111010010010101001111001001001100000000010001100111011010011110011110110111100101111101100110000101011100101111110100001101011110111100000010000100000100110001001010111010010001001011111110010010010000;
#1 $display("%b", po);
# 1  pi=207'b110001010110111010000100111100100101101100111010011001011111100010001011001010100100011000011110000000110010010101110011111000110010001110000100101011011111010011100010001001111000110001001010100110011010011;
#1 $display("%b", po);
# 1  pi=207'b010111100000111101110111101100111010100100110110001010101101001010110010110100000010110101000011001101101111001001010010000011000111100010101100010110111110001101001110011111100110111100111101100111011101010;
#1 $display("%b", po);
# 1  pi=207'b011111110011011000101111010001001101001010100010111010101110010100000000000000000101010111000101010001100011001000010010001000111010001100010011011001010111100110010110111111111101101111111000100101001101110;
#1 $display("%b", po);
# 1  pi=207'b101011010101101100000010010000000001011001001000101011100011001001010000100011111010101011101010000001110100101110110101110000011111010110011001110101001100110100110000011111110010100111100100111010110101001;
#1 $display("%b", po);
# 1  pi=207'b000101000110000011111110111000010010011000101110001011010101010000100010000110111011110110001101111101101011110000000110101111101011010110011010110111011100001010000110101010110101100111101100110010001111110;
#1 $display("%b", po);
# 1  pi=207'b100101010011111111000010110100011100100110010001001001001001001001100100001100010000010000010101110111111001000000000010001111111010111000001001101000111001110100001000011000110100100001100010011110001011111;
#1 $display("%b", po);
# 1  pi=207'b011011101100000001101010110110100011100000110111110111100100110010000011101111001000011001011111100110100101111101000101000110111001100000001101000111110101000000110100100011010111110000111100010011011011011;
#1 $display("%b", po);
# 1  pi=207'b000010111001111011110110000111111111101100110101111111010101101000111111000101000001110100111110001101100101010011010110111000011000010111000011100011010101111110101100011111111110001100111110011010011100001;
#1 $display("%b", po);
# 1  pi=207'b101101010101010110000101001100000100000001001011100000010110010001010110010000100001110010101110010010111010111111010010000011111001100011100111111000010011100011100111011101010111101010101110010000001101010;
#1 $display("%b", po);
# 1  pi=207'b011110110010001111101111100010101110100010101001011011011000011100001101011101011110111111100011101101010000111000011111100000010000010110101010001010111011001100011111001000111110111010011101000100101111100;
#1 $display("%b", po);
# 1  pi=207'b100010110001010111111000101110101001011100110000101100111001111100100011001111100010100011101011001110111101100100101001011010001011001010111010100011010010001100110101000110010101001001011100110011100110001;
#1 $display("%b", po);
# 1  pi=207'b010111011001010000001101110111010010011011111001000000000111101110000101101110101011110100101010101110100100001100000001111001110010001101011111100100011001100001011010010111000111001101010011010000101001011;
#1 $display("%b", po);
# 1  pi=207'b001101001011100111000101010011111101000101100110111110110010101011111010001100000100010011111000100011001101100000110111001010111110010111001010101101111010000001010011010011001110001000001000100011110011010;
#1 $display("%b", po);
# 1  pi=207'b100101110010001101000001100101010110011111110011010010001101111010000100000010010110100000100011010001010001010111111011111001010000010111111100001111110100110100110011111100001111110010010100000111110100110;
#1 $display("%b", po);
# 1  pi=207'b011101111010010011111110000110010111000011001011000000110010111001010011011011101100010100000110100100010100011000000110101010100000100110011101101000111010111010100111010010001001010111001100001110110010000;
#1 $display("%b", po);
# 1  pi=207'b110010110100110001010011010011110010001100010101010011001110010101101000001110011001000101011110100101110111010001010001000010011110101110101010100011010110001001000111010100011001101010110001000111000000111;
#1 $display("%b", po);
# 1  pi=207'b011010110100111101001000111100001101111110100001011011101001010010010001000001010011101010000001110001001111010101010000111011010111001010110000101010101101000000100010110100100010101010111111010100011010010;
#1 $display("%b", po);
# 1  pi=207'b111010101010111011010111000100110110100000011011111010111110011000010001000000111111110010000001011110101001110101000000100010010001101110110110101000100001111001101111100010111111101011000000100111110110010;
#1 $display("%b", po);
# 1  pi=207'b000000101111001100011001001001110010001010000000100011011000010001100101100111001100110101100100001101110010010100010011100001011100001111011101000110011100111101010011111011100111011100110110100110111110111;
#1 $display("%b", po);
# 1  pi=207'b010001010111011001011001100111010011101111110100111011010000110100000000010000100100101111110111001001011100010100110000111000010011111000110100100100000101001111111011111101111000010001110101010001100110101;
#1 $display("%b", po);
# 1  pi=207'b100100110011001110101010110101111000000010000110010110110010011011111011001111011110010100111110010010101100000101000111000001010111011000011111111100111010100010110001011010001000100101111100001011001100001;
#1 $display("%b", po);
# 1  pi=207'b001101101111001011001011001101011011000101110010001001001101100000011010111010101110101000000100101011000010010111111010110001111011110000001110001010111110101111011000000101001001011011110110111101000101000;
#1 $display("%b", po);
# 1  pi=207'b110001111101010110111000001001010000001100101111100101011001110001101011111100001101011110010111110000011001000100101100111000110001001111110111110110111111100000101010001011000111111111101010001110001000100;
#1 $display("%b", po);
# 1  pi=207'b010100100010101111000110101100110110110011100010010011010000001000110000010101100000011000111010110111011010010111001010001001100000000010100000101001111000010010111011100110001011001101111011111111001101011;
#1 $display("%b", po);
# 1  pi=207'b101001001000000111000111101010100110011111100110011100000011101101101010110010000111001000100110010101111111111110101111100100110001101011000010110010101100000011111000100000101100110000010000000001010001010;
#1 $display("%b", po);
# 1  pi=207'b111000100101101001001001011111101101110001100001000001011001111001101000001010011111010101110101010110111010010101101111010100001101111101010000111101011000101011111101111111010100010001101111101100000100100;
#1 $display("%b", po);
# 1  pi=207'b011001000011011101100000110011110110100011111111010000100011110001000110110100000111100010100111010111111001001011011101101100010110101100011010010001111111111110001001011111110011000101110010000110100100110;
#1 $display("%b", po);
# 1  pi=207'b010110101000101100111010011100111001110011110110000111111111101110110100011011000101100111001010101111110001001001011110101000001001010000000110011110001110111000011010111110001111000010100101110111010110110;
#1 $display("%b", po);
# 1  pi=207'b110111011011000000001111000000010001000100000010101101100001001000010000011110110111001111100000010100111101110110100101111000100001010011001000010011110001110110010001101110011010111111000101100100010101100;
#1 $display("%b", po);
# 1  pi=207'b100100111111100011100011000010111100011111010100000001010000111101111011110011100101110000111110011000101111111001111000110011110010110010001000100111101110110011011001000010001110111000111101011100011000111;
#1 $display("%b", po);
# 1  pi=207'b101100010110001100100001001110010101111111001011001100010101000001010110110010010100001110111010100100101001111110011101110111010101100111001110111110110101101010100010000010111101101100001000011000110010000;
#1 $display("%b", po);
# 1  pi=207'b010101111001110010010001110100001011110111101011101110110010101110000110010001010001100011110101000000000011010010100001011011000101111010110111011101110000111001111001101100101011100111001101111011001111000;
#1 $display("%b", po);
# 1  pi=207'b010011111100111011101101011010101010000110110000011100000010100000110101110010111010000000111100101101101011010101001001111000000111011100010101000010011110101000101100010010011011110010001110101100000111101;
#1 $display("%b", po);
# 1  pi=207'b111000111110111101100101001001110100101010110010110010111010000001000011011100001111110101000001100011010000010010000110001110110011100001010101110000010011010101000111001110001110101011110100111000010010110;
#1 $display("%b", po);
# 1  pi=207'b101111100101010010111111000000010101100011000011010010101011100100010101100100001101011011100101011001110101110111010000011001100100100000101111001011101001011101000111111010011111000111110111001000101111001;
#1 $display("%b", po);
# 1  pi=207'b111110011000111011100101011110101000011100011100100110100011001001101100100101010011100000010000001001001000001100010100100111001111111010011100110011011110111111010111101001010101000100010000001110000001100;
#1 $display("%b", po);
# 1  pi=207'b000100011110011110010101001101111010100101100111110100100111101011010100100001011110001011011000001010110101111000000011101001000110010011011111101100100001110000110001100010101100110111101111011101000100111;
#1 $display("%b", po);
# 1  pi=207'b111000010101011000000100001110110110010011000000001101101000000101010101101011000011000100010101010111010101011000110011111100001010100111100011000100111011111101101010100001010010001110111011000111000000101;
#1 $display("%b", po);
# 1  pi=207'b001000100100010001010111111000100110011101000101001001001101000111010111100000101001011110101010010101001001111001101010000111010101110000111101111011110010010011000101001000111111110000111111011101111000011;
#1 $display("%b", po);
# 1  pi=207'b011000000011000101100111001011000001010010010000000001010001110001110001110100011110010111001111111100011011001001110101101000001110101000011000111110011100011100010110001110110010101111001100010000110111011;
#1 $display("%b", po);
# 1  pi=207'b000100110010111101101110110101101010111000010000011000010010101101011011101011111100000011010100110101011101111101010000001011011100110010000000100000010001010001011011101010100011010101000011001110000011010;
#1 $display("%b", po);
# 1  pi=207'b100100001111110101000001100011110101100111010111000001110010000011101010001010100011001011100011011001111110011110011000011000111111111101010110100111000001000000000101111101010010100000011101010011111110101;
#1 $display("%b", po);
# 1  pi=207'b001001010111010100111111101001100011010101111110010010111111011100000101111100100011111010000011111101011000001111110001110010011111101001110101110001100011100011110111110110010011011110000010010010010000010;
#1 $display("%b", po);
# 1  pi=207'b100100011100110100111010000000010101000110010000001000101111001111100001000110000110100101000111001001100001110100001010100001011110001010000010111100101001000100101111110010011001101011100100000110011000111;
#1 $display("%b", po);
# 1  pi=207'b001100111111010000011000010000000000101000000011100010000110011010110111011010101010001001010110011100010010000011011011111000110110100010000101000001101110111001100010000111010100010010010011011111101010110;
#1 $display("%b", po);
# 1  pi=207'b000011000101001110111100110010011011110000011001101100001110111101011011111010011110011101000101010001111111110011111110001011100011100011101011010011000011111001000010111010001100101111110011111100000110101;
#1 $display("%b", po);
# 1  pi=207'b101011100011101010100101100000111100000100101011011010111010001110101101100000100000110000011111010001001000111100010001000011101010110110110110011110100110111111100101001111101110100111111101001110100101101;
#1 $display("%b", po);
# 1  pi=207'b010110000101110101010001101110010100011010100010100000101000001111110101110100110010011011001000100111110111010011011000011110010010101100100101110101000111111010001001001110101100110010101111001011100110000;
#1 $display("%b", po);
# 1  pi=207'b110010110110000100100010110000001110011001110000101011111000111110101010011101110010101100000110001011011110001000010011011001111100110011101001001000100110111000011110110010101011111110001001001001101110010;
#1 $display("%b", po);
# 1  pi=207'b100010001110010101011000111001010011110101111110101000111100000000001110110100100011000111110001111000101100110100100111111100110011000111011101101001000111011001100010101110011000010010111010000101001100010;
#1 $display("%b", po);
# 1  pi=207'b111010001110101010100000100110110101111011111000000001110011110001001101001011111010100000111011111010001110100101111001111111101010101001001010011001100100111110110000100111110100101110011011010110100101110;
#1 $display("%b", po);
# 1  pi=207'b011000101111000000010001110110111101000110101001110010011000101010101111111011110111000010011111011010010101001111000000100010100011011110011000011000001101011001000011111110010011010111001010111101110100011;
#1 $display("%b", po);
# 1  pi=207'b000000010101100001001101110111111100111011110010001110101110111001110011010010110000111110001000111000000101010010011010101100110111111110110100101111111001010010010111000010110010101001111110011000010110000;
#1 $display("%b", po);
# 1  pi=207'b000011001101000011101111100100011110010010111001001101000010010111001100001000101100101100000010100000001100101100010001101011000000101000110011110010111010001111100110011001011100110100111000100001011000101;
#1 $display("%b", po);
# 1  pi=207'b101010010001001001010100011010010001000110011001001110011000010010000111000111111001110001100100101001101100001010110100000000000011011101010001010011001111001101001000100101001011101110010110010000000001100;
#1 $display("%b", po);
# 1  pi=207'b111010000011000110000100111011001111100000010011010110110000001010000101000101001001011000101011100010010111101100010100111100011101000101101010101110010101000010101011101011011011111011110111001010101011111;
#1 $display("%b", po);
# 1  pi=207'b110011100101110001000110100101110001010000111010110100000001001111101110101001110100101000110101111001111001001010110101111110001000000001001111010001010011110110000010101010000001010110011100100000010101001;
#1 $display("%b", po);
# 1  pi=207'b101010100101011110010000100100010010110101101101110101001010010100001101010011011010000010110001100000101110000111000010100010011101111001101000010110000001000000100111001010011011011110110100010011011001000;
#1 $display("%b", po);
# 1  pi=207'b010111100110100110001001010001111010101000001110001110000110110101111001010010111110110110110101011100110001111000110011110000111000001001010000101110010110001101011101110111011100100010111001001111000000001;
#1 $display("%b", po);
# 1  pi=207'b100100111001101111000111011001001101101111001001000110000101001100111111101000001010010000001001010110011101111111010100101010110110101100101011011011110001110000110010100110011010100110101100110110000001110;
#1 $display("%b", po);
# 1  pi=207'b000001001101100101111000000110001101010111011001100000000111000101000000110100111000111010010010101001000111010001110000110001100010010111011100110100010111010001011101010000000000101110010000111101000111011;
#1 $display("%b", po);
# 1  pi=207'b101111001100000000100000101111110100000101101001110011000111011110110100111101110010110001010011110100101001010111001111000111100110100101000111111110101000010101101001111110101100100100011111111000101101001;
#1 $display("%b", po);
# 1  pi=207'b100011100011010011010100110100011000111001010010101101111101010010010110010000110111011101011101111100111101001111000110001110011101011101110011001111110010010101101001010011111101101010111011010110010101110;
#1 $display("%b", po);
# 1  pi=207'b111011001011110100101000010111001001110010101011101001000100010111110110000100000011110111111101011110000101011100000111111100011011011000010000000000010111110111000110110110011101110111101011010111010000101;
#1 $display("%b", po);
# 1  pi=207'b001111101011101011001111011100010001000000101010011111000011101100101101010101010111011011111010010111000100111011101000010011111100110011110101110100110110001111000011100101011100010101000110101111111000001;
#1 $display("%b", po);
# 1  pi=207'b000011111110000101010000001000110011101000011100111011010001011101101011100001110000100111000111100000101101101000101110110010010110000111001010010000011000100011001101001110010010111100101110100100111111011;
#1 $display("%b", po);
# 1  pi=207'b001101110111100001101101111111100001010011110001000001010111001110111010011101001010101011011000101101000010111110110011100101011101110101001111011110110000111111000010101111100111101111011100010100001100001;
#1 $display("%b", po);
# 1  pi=207'b001001101011011011000110100110010111101011000010100110101011110101110001110000000111011110111011110101011101011101010110110100010110110011010101011001001010001111101111000010000011011011110110111001001111011;
#1 $display("%b", po);
# 1  pi=207'b101011101010000110101101001011111010010000010111110101010110100011110110101010000011100001100101111010000100111100100000010010100010000000100000001101101101000101001101100110101100001011101100000001100001000;
#1 $display("%b", po);
# 1  pi=207'b000111010011001101011111011001011000111001001010110000011110111100011011000001001111011100101100000110110011110101001101001101110010101111001100101100101101011000010110011101010010010010010000010100110010000;
#1 $display("%b", po);
# 1  pi=207'b011101000111100101001100100100110100111110010010011100110101110111100010111011001100000011100001110010001000110110101111000000111110101101000000011000111101011000101001110001111100010110111101101110010100110;
#1 $display("%b", po);
# 1  pi=207'b100000011001110011110101101100101100100000001110001001000010001110110101111111001111101000100100000001111000111101100100010101100000000111001001100010000000000110110101101110011101011001100110110110110010000;
#1 $display("%b", po);
# 1  pi=207'b110001011111010000011000010101100011111111010000101100110010000010001000100101011001110101010011010000110011110011100000001000101001010110101101100100000000010101000011101110011101011111010110011111011101101;
#1 $display("%b", po);
# 1  pi=207'b110101111110000110010110101011010000011010000101000100000110001011011100100001101100111100000010100101000001110111111110011001010011110010000101010000011100110110110011011100110111000101000010110111111001001;
#1 $display("%b", po);
# 1  pi=207'b110010001000101101110111101001010000010001101000000001100101110101011001001111001010001111111111100111001101110001111010011010000101011100001110011001010010000001011011101100111111000101001101101100010111011;
#1 $display("%b", po);
# 1  pi=207'b100000000100001001011010001001000111101000110101100110001100111100011011101111111001111001001101111001010000010001110111100001100000010110111010000100101100010111001100011001110001010010000101000100110110001;
#1 $display("%b", po);
# 1  pi=207'b101100010001011110101010001011110111111111011101111011010101011111011110011001100000000111011000000010000100001000011010111110000110111000111111000011010011010111011000000000001011111010110011010100100111110;
#1 $display("%b", po);
# 1  pi=207'b000000101100111111010111000011011000001111101111001001111001101001000000111000101110010001110110100100000111111101001110000011001110101010111001010011000011000100110010101000101111010010111010000010000101000;
#1 $display("%b", po);
# 1  pi=207'b111111111011110110100000000010111110100001110110110001000110001110010010010000100111010110000011001001001000010100111101001111000101011111011010010011101000001100010110110001100000101011000111110110111001001;
#1 $display("%b", po);
# 1  pi=207'b011000111000000001010101001010001010111010111111010010000011000110100101101110110110000101111101100011101011111100011101100100101110011000000110101011101011010101000011101100000111000000110001101011010011000;
#1 $display("%b", po);
# 1  pi=207'b010001010100111000011110010101011011010111010101010101111100110011000000111011101000101111010011000100110111111100111000000010000100001100100010111001000000001010101111110010001010100011001001000000000010110;
#1 $display("%b", po);
# 1  pi=207'b101101111111011001000011001110010111101100000001010101001110011100010011011111111011111001100010001011110100110100110010110000000100100000011111101100101100101101010100110100010000110001001010001000101101110;
#1 $display("%b", po);
# 1  pi=207'b000001010110001110011110011010001101000100010010100010010011100110000011011000111011110011011010010000111111110100110101000100111000110010110000000101011111110000101011010000011010101010000011010010111010110;
#1 $display("%b", po);
# 1  pi=207'b110111100101011000011010111000010100010101001011110110011010011011010100001111000010110011100101110000101001000001101100110101001000101100101101100111011100101010000000111011101000001001100110111011011010010;
#1 $display("%b", po);
# 1  pi=207'b011110001000001100110101111101101111001111111001001001100110011000100111001110111010110110001110100100001010101000010011101000110010011000111110101111010111101101111001101111000110001011101000011011111010111;
#1 $display("%b", po);
# 1  pi=207'b100111011111000000111011110011011010000100010011101100100111010010101001011111011001011001001111000111110010000111000010110001001110010110000100101111011000001110111000011010101100000100110001101100010110101;
#1 $display("%b", po);
# 1  pi=207'b101111111110110111100001111000111000011011011000000001110010101011110100101000101110101000100110001000110110111111111100011100111111000010010011111100101111100100100010101111101101110010110011101111010111000;
#1 $display("%b", po);
# 1  pi=207'b010111111000010000110111001111010011000100111110100100000101001110101001101100001110001110101101111000001011000011000000110001011100110100101100101100111101010011111100100000101111000010001110011110001011000;
#1 $display("%b", po);
# 1  pi=207'b011110001011101000111000111000001011010001001010001101100100111001101010111000011110011110101111111111110100100101111101110101101010100101010011001110001111001110000000001011110100100010000000100000101110111;
#1 $display("%b", po);
# 1  pi=207'b010011001010010111010001001110110010111000111000110001110100001011011001101110101110001110010010010011110010010000011000000101111110010110101101000110001100000101000010010101001100101100001001100100110111100;
#1 $display("%b", po);
# 1  pi=207'b101111100100101100001110011101010000000110001101100101100001000010111000001100010111010001111010100000100011001100100110010101111000011110000101011010010010001011100100111111100101101001001101101000110110000;
#1 $display("%b", po);
# 1  pi=207'b001110111101110001010001010000100111000101001111011011100010110010011101011011010111001111001110110100100000001011100101001100010010101110000100100100100101100101010010100000000100011010101101010100000011000;
#1 $display("%b", po);
# 1  pi=207'b011110010111011001110011100101101011011001000010101111011001111111100000110100010000110101010111000001001110110110011001011111000100111000001010000100111101100000111110110111010110111111111000010111111001010;
#1 $display("%b", po);
# 1  pi=207'b001000010111001100101101100000111100100000001010110010011110110111100110010111111001100100010111111110110111110000100110001100110001010111111111010100000101010000110101010001010101110001001100000111111111011;
#1 $display("%b", po);
# 1  pi=207'b100101111101101100100010000100110011001001111101000011011100000110000101101011000100001100001001111001101001111101000011101110011010111101110001111100100110111111001011110100111001010000111100100101010101110;
#1 $display("%b", po);
# 1  pi=207'b110110000110100010110111100001111101001000101100100010111000101010100011011001101011010011101110100100100101010100110110100101011111110000111101101110100100110001110011000110110100110001101010001000011011011;
#1 $display("%b", po);
# 1  pi=207'b111111101110001100101100110011111010101011110101011100010001100111011100101110010011101101001011011011101001000000000111111001000010101011100001110100010001100001000011001000111001011000011010101000100001001;
#1 $display("%b", po);
# 1  pi=207'b011111111101010011110010111100101000111110001001001100011110000001001101010110110010011100110110010010000110111001101110111101100110000110100010000100111111010100010011001101010000011110110000101100001111010;
#1 $display("%b", po);
# 1  pi=207'b010100000111001101011110001100111101010000011100101001010010011010001000000111110000100110011101001110001111101001100000001101011011111001010001001011001000111111101111010000110101001110000001111001101100111;
#1 $display("%b", po);
# 1  pi=207'b010101001111011001110101010000000111011101011010111110000000010111001111110011001010010011000001111100010000010111000101111111111011000011100111001000000011111000001010111010111000101111011001111101101101001;
#1 $display("%b", po);
# 1  pi=207'b100111111001100111001011011000100100110010111011110100010111110000011000000011001000100011100100001111100011010010000000010110101110000110001110101010001101111111000111101001010010110110100011001111011110101;
#1 $display("%b", po);
# 1  pi=207'b010010011101101101101000110101101010010110010011011001010000110011001000010111100100001100100010111101101000100000000101101000000010011100010101111110101100101000001010001001101001010000100001000111010100001;
#1 $display("%b", po);
# 1  pi=207'b100111001000100010000100000001000110111010110000100111011001001001000001100111001100010011110010100110011000011110110100011111100001111101010000011100111001111111111111110011000000001011110100010111010101000;
#1 $display("%b", po);
# 1  pi=207'b001010011110110110001100100010101001100011001011110100011011011000000111111000011010110111100010000101100010110111100011010011000011100011010010110100111000101101111000100000110010000011010011111100100110100;
#1 $display("%b", po);
# 1  pi=207'b011111110011111001011111001110101110100010010110111110100011101001110011010010011011111110111000011000001101011110100000101100110110111001100010111111110011110111100110011110011000101000111010011110001110110;
#1 $display("%b", po);
# 1  pi=207'b101101101100100111110000101001110111111010010111000011010111000101110011011101110111110110001111001010100000001101100110110011000001100000011100111100110111100010001101101101101000110100000000101101000111000;
#1 $display("%b", po);
# 1  pi=207'b011101010001001110000011110110000001000111001111101010101010100010101011001000111011100001100001001000010101000001001111110000011001000010111011001001000100001111110010001010100101000111011111001110001000100;
#1 $display("%b", po);
# 1  pi=207'b100111011101101100010001000001001100010111111000111101111101011101110110110101011000010110001010110011000011010000010001011000101001001001101001001001111000111101110000011110001000011010101111110111010110101;
#1 $display("%b", po);
# 1  pi=207'b110010000000001011001001111000110100101000011101111110001011001000110101110001010100011111111101111110011010110100110001110000010110001001000001110001011000000001011100011011000110000010101011101101100110010;
#1 $display("%b", po);
# 1  pi=207'b100011101011100011010101100011100010111011100010110011001111001010110011010000101100010010011011101100100010011000111100001111000000101000010100010001101111011011001010110111011111011000100101000010010000001;
#1 $display("%b", po);
# 1  pi=207'b011011110101101110011110100011010011001010111110001010100010110001110111010100101011110010011001110101101100100000011110010101111110000000110100100000100000000111110001010101011100100100001110001001100100100;
#1 $display("%b", po);
# 1  pi=207'b010100111100100100111111010011000111001000111111011000110101010010010110110101000000000101110101011010010100111000000100000001010000111101000011001101111101001100100101110101100000111111100110001111000010000;
#1 $display("%b", po);
# 1  pi=207'b110000000110101110111010010010101111111000111000100110001010000111100010001000010101000110110111101101001000100010111100100111100100010000000101000001110001010000111001000100000101100011101101101110100001011;
#1 $display("%b", po);
# 1  pi=207'b101001110011101001110010010001110000110101010111111011101000010100110000010010110011001010111000110011000010100100011110011010001110100000000111111110100010001010010011001111101011101100010001100000000111011;
#1 $display("%b", po);
# 1  pi=207'b000100100000010010111110111110101010100001101000010000001010100101111101010111111110001000010110011111010001010100010100010110000101010001010010100110111010011100011010000000011011110110100000110110101000001;
#1 $display("%b", po);
# 1  pi=207'b011101111111000011000101100011010110101000010101101101111000011110000111111111001111000110001010011011010001000011000010100110110011100100111100110101000000001000100110010011101101010100011001110111100000010;
#1 $display("%b", po);
# 1  pi=207'b110010000010011101101000101100011011100101001010101010111011001101001110011101000110010000011101110110001111001011101110100100000101100000000000001000110010110110110110001110100010000001011110001101100100001;
#1 $display("%b", po);
# 1  pi=207'b001100010100001111101101100011011101101110001010011110011010000001010000100011111101011011010011000011000001010111111001000100111010111000100100010001101001101010111011101111010001111000101110010010010100000;
#1 $display("%b", po);
# 1  pi=207'b001101100100110101010010001101101100110100110111011011101011010111010001001100101010010011001010100111010000010101000111010100100001110001110000101100111011011111010101011100100111111110100111111101001001100;
#1 $display("%b", po);
# 1  pi=207'b101110010010010111101110001000111101001111100110111110111101011100000101000101100100010100110010001100110110100000010010001010111111111001110010010011101011111011100010110011000101111011100001111000000011000;
#1 $display("%b", po);
# 1  pi=207'b111111001010001110100110000011100001100101010111101011110111001010111010000111001000001101011000011110011001111010111101010000011111110000010011110010100101000100111000110001111100111000111011101110010001001;
#1 $display("%b", po);
# 1  pi=207'b101111101111000111100110001001000011101010000011001100011011001111101010111010100010111011101011101110001011100100010111101111000000001010110011011111100101111011011000110000000110000110010100111101000101110;
#1 $display("%b", po);
# 1  pi=207'b011111000111101001110101001110100101101101010101001010000000111110111101011110110111111111000000011010111111000110011110101101010110100100100110101011100011101111010001100101010010101101111100101001011001110;
#1 $display("%b", po);
# 1  pi=207'b110100001110011010000001111111111110110110011111100111010000001010110011111100101010111011101111101000100100110011000000000110001010111011100010001010001111011101001101111010100001101001110011011111110111001;
#1 $display("%b", po);
# 1  pi=207'b100110111010001110011100111001110010110110100101100010110011111100101010010000111011011110110010011000000101100111101101000010101101111101011110011100001010101100100100001111000000101111000001110101101011001;
#1 $display("%b", po);
# 1  pi=207'b100001010101000010010001000001111010010100100110100001101110111010011100101101110100000001100111110011111100000001100110100011010110101110110100010011110110011100110101111000010010101011001001101111101000101;
#1 $display("%b", po);
# 1  pi=207'b100110000011010001010101111011111001001000000001010010101001001101001100111011000111011011010010100100100000011010110011001111001100101010010101110010000100000100110000010101001101000110100110010110101110111;
#1 $display("%b", po);
# 1  pi=207'b101100101110100011100000110001111011100110011110000100101001010111100001001000011110000011101100110101010000011111001100000110001111101110001010010000001000100010111001000010000111100000110001010011011000010;
#1 $display("%b", po);
# 1  pi=207'b010100010011001010000011111000010110110011110111101100000100101100101100000000100101110010111010101111100001000011000111000100001110101100010010000010001000110011111111010010100010101010101010000001010100101;
#1 $display("%b", po);
# 1  pi=207'b001001110111000011100010101110001010000001110011111110110001110010111100000010001101010001110000110100010001010011110000010100000100011100000011101001010011101010011000111111100110010010100100111100010000011;
#1 $display("%b", po);
# 1  pi=207'b001011101001100101001011101111001111000110101000100010001111001001100011110011010101010101001110100011000100101110010010110010101000110100010001011000000110110011010001111011001110000000011100100001110010011;
#1 $display("%b", po);
# 1  pi=207'b100110100010100110100110110100110110101110001111100011100110100110001101110011101011011011011011110001001100111010110011000101100100111100001110010111110100010010000011010110011110100100001100001000000010111;
#1 $display("%b", po);
# 1  pi=207'b100000111010010111010100011111101000100001011001100101000001000101010001001111100111010000101001111000110000110000100111110101001100011010100111110101000010000011011010011000011011011111101101011011111100101;
#1 $display("%b", po);
# 1  pi=207'b010000111000101110101011101010111011111111011111110011101001100001100010010100000011111001011101110010111000010000111110100010100100010000101111100011110000011011010000111100011111000101101011101000110001110;
#1 $display("%b", po);
# 1  pi=207'b111010101011100010011110000010011101011100010000101011010101110100001011111001001001111111010011101000100010110110100010011011111010100101110110011001110001011010100100001100110111011000101011001000001111110;
#1 $display("%b", po);
# 1  pi=207'b000011001110101110000010001010011010010010110101101110101110010000101110101010010001101100100000000000001100101011111101011010111110001010001000111001101010001101010100101111001100101101101010110111011000010;
#1 $display("%b", po);
# 1  pi=207'b011101011100110111010100010000100011010100100000000110010000001010011101111001111001100011000101100110111110110110010010011011010100010110101111000110101111101101000111000110010111001001000100001011010001101;
#1 $display("%b", po);
# 1  pi=207'b110001011110010100100101011110010100110010011101011111100001111111000010101101101001101100010111011100111010011000110001011000101110000111110110010001001010100100110000100111100101111000100010000011110001101;
#1 $display("%b", po);
# 1  pi=207'b110100010010110001001111010100111110101010111111100011101001001111111000111110011110010110110111111110111010100111110100000101010111110101111001101110001101110101101100100100001110001001001011010111101001100;
#1 $display("%b", po);
# 1  pi=207'b011000000100010100111110100001101100000001101011000110000011110000001010110010010010010100001000100001110100010110100011011111110100010100011110100001010110010111101001000010100010111111010010100010010010111;
#1 $display("%b", po);
# 1  pi=207'b101111111000000010011101101110011110111111111001101000000000101111101110010000100101000100010011010001100000111101110001000100001000101111001101011011000000010110011101001110010110100111101010110101001010110;
#1 $display("%b", po);
# 1  pi=207'b000010000010100101001100100110010000000111000100011100001110001110010100110001101000111010110100111010111110000111011111101101111001001110101001010001011000110010110110001010110000110100100010011011011110111;
#1 $display("%b", po);
# 1  pi=207'b010010011001010110111001011111000011010111101010110111011100000101101010001101100011110110100001111001101001101111011001110100101010111010010101110000110011110111110010111010100100110101010110001010000010101;
#1 $display("%b", po);
# 1  pi=207'b000111001100111011101000100111000001010011010010001011001001000010010001011010111100010101100011111111011110110011110100110000111000101000000000001011100111010000001010100101010000000110110011111110000001011;
#1 $display("%b", po);
# 1  pi=207'b011011110111000000100001111001100001011011000000011001111000110110010000011011111101100110001110110001010110001001110010101011010110011110101100001000001100000010000110010011110000100011000101101001111000010;
#1 $display("%b", po);
# 1  pi=207'b110000101111010100110100010100011001011111101111001001111110011101010110011111100101001000001000010100010010001000110000100001101011101111111010110010110110011111000000001110000110111110100000010011001010010;
#1 $display("%b", po);
# 1  pi=207'b000100010010101111111010110100011101010010010111011011010000110000100011010011000010011001000110011011001110000010100001000111100111111001000001011011101011000011001100100110110000100000101100010011000110011;
#1 $display("%b", po);
# 1  pi=207'b011111001100000001001001011101010010101010010001000001100100000101111100111101101101101000001100001110001011100010110011110111000111100010100011000110101000001110000111001100001101010110110010100010111111110;
#1 $display("%b", po);
# 1  pi=207'b110101101110010101110001111000000000010110011101100011100000011101111001000100010100101100110111110010001010010010101100001101000111100110000011010110011011011010110010001001100000101001101110101110101110101;
#1 $display("%b", po);
# 1  pi=207'b100010101101100111010010010010110011000000111001100011011110110110010001101000001011111000011011000100011110001000110010111011111000010011111110101011010100001001111111111010001010000110110001000101011000110;
#1 $display("%b", po);
# 1  pi=207'b010101110010001110001101001001111010011101101111001110000010110100111110111101011001010110011100001101100010001110001011101111100010111101101111100101001001100111111111110010110110011111111110110000001111000;
#1 $display("%b", po);
# 1  pi=207'b100000101110011100111010010100110111111100011111011001000001101010000110111010011110010110011011000110111110000011001100001100000101101101001011011001101010111010101011100100001011000011000000010110001111000;
#1 $display("%b", po);
# 1  pi=207'b001101010011110000010101011010101100000010110110011100001110000010010011001000110001100100011100111000000111001011001000110001000001001001000100000111110101100011100111001000111111101011001011011001111100101;
#1 $display("%b", po);
# 1  pi=207'b101001011101111101010011000000000110100001000010111111000110011100111100110101110000100111010000011100101000110101111111111100001110110111011111011111100011111111011001001101011111101011010001110110110000100;
#1 $display("%b", po);
# 1  pi=207'b000001111000011000000000101100100101000011100110010100011110111101011100011101000110001111110000100101010101011101010001101110101101011100100110001011000111001010100100111011000001011110100100100111001001101;
#1 $display("%b", po);
# 1  pi=207'b001000110010100111001110101011000001011000100000000000000111010001001100100111101110001011010101001010010110011000010000100010100000010101000100010011101000001010011001110011110100100001000100110000110010100;
#1 $display("%b", po);
# 1  pi=207'b010100101011111101110110110011101110101101001001111111100011100100000101001111001001101010101101110001111000111010010111010000010000010001110011111010101100110110010101010100100000001111111100110011110111111;
#1 $display("%b", po);
# 1  pi=207'b100010100101101000000000011000100111100111011101000001010111100000101000110000101101000101010000101110111000110101001010001011110010011100000110001010010110011100001111111001001010100101100011100100101000010;
#1 $display("%b", po);
# 1  pi=207'b001001001100001000010110100111000100111001101101110000100100101000101100100010000101101111111001101001000101100111011001001000111001000011101011110111101101101011010100101000101000010000010011100110100011110;
#1 $display("%b", po);
# 1  pi=207'b101100010100101101110101101100110011001011101000111101011000001011101011011010101111000010111000110011101101011100100000100001001001100110010011100100011001010100110101101110111001011001101010100010011110101;
#1 $display("%b", po);
# 1  pi=207'b011111111010101001011101010011011010110100010111000101110011101111110010000001010011110011000101111100111010000101101000100010000001000101001000101100010001011011101011000001000101010011011011100100110000111;
#1 $display("%b", po);
# 1  pi=207'b111100011110101111001011010100001100011011100010110111010011101110011111100100010100000001111011001000111110101010100111001100010010110011010000111111110111100010000101001010101001101110111111100101001111101;
#1 $display("%b", po);
# 1  pi=207'b010001000110011001100101111011110110100000110011001000100111110010101011111101110001010101000011001011000110101101110100011010100010111011011111111010100100101101010111011010101001100100101101110000101100101;
#1 $display("%b", po);
# 1  pi=207'b001101101111110100100110011001010111111010111011110111010100100101110110100011111111101111100100111111110001000110110100001101101100000100111111001011110110010101110011100000001000010000110010111111010010101;
#1 $display("%b", po);
# 1  pi=207'b111000011010110010000010001101111111100011011100101011011001000100010000011010101010011000001100101111111111101111100000010110101101000010000111101011001101110001101011111101011101010101010101010011100011111;
#1 $display("%b", po);
# 1  pi=207'b100001001101110000110010100110100000101111111010111000000110101000101110100001101110100111101101001010010100011101011001111010111010010100110011001011011000111001111010100110111101010111100010101100001100101;
#1 $display("%b", po);
# 1  pi=207'b101001101101011111101101100110011000010001100000011101000111000100111001000100101000101111001010010110100011100010101100101011111010010101111011111100011001001000111110100110101110100001011111000101110011100;
#1 $display("%b", po);
# 1  pi=207'b101100011101001110110111011101000110100101000000001101011011110110010110110010010001011111111011111010000100001001110111000000110111111001100011100010011011100101000110110011100010100010010111111011110001001;
#1 $display("%b", po);
# 1  pi=207'b111111111111100101000011010110101011101101101011111110111100110111101111011100110011110111001110000110111110001111001110000100111110011000100011101111111110001000011011000111001110011101000110100011110101000;
#1 $display("%b", po);
# 1  pi=207'b001010001110111010011101001000100000011111101011101111101000000110011000111111000011000001100110010010110111110010001101111000101000000011010100110111110011101010100110011011010011110010001010100110100101001;
#1 $display("%b", po);
# 1  pi=207'b001101101010010111111011101011101011001010111011110101001010100101010111100110011001110111110101111010011110000111010110100011001011111010001001011100111111101110010011110101011000111100010000001101101011110;
#1 $display("%b", po);
# 1  pi=207'b000001110011110010010001100110110100000001000000100011001010110000001010001111100001000111000100010110111110010010001110011110000001000101100011001010010000110100001000001000100010000111011110000111101010111;
#1 $display("%b", po);
# 1  pi=207'b110011011110010000000001000101000101111101010100000001101110100111010101001110000001001100111110111000010001011010001111100000001110111111101101000001100101001010110010101011110010010101100111011100111011110;
#1 $display("%b", po);
# 1  pi=207'b101011100101001111000001110110110011000111100000001011000010110101011000101011010110000011110010111011110010000010111011110111011101110100011001100110100010110100011000011001100100101010011010010110010100100;
#1 $display("%b", po);
# 1  pi=207'b010111100110101111000101100110101110100011000111001001011011110111110101100101011101011100110110111101001010001101000110110101111111111110110111000100000101111011000011101010100101111001001011110010001100101;
#1 $display("%b", po);
# 1  pi=207'b001000010111101001101000011111010111001011010011100011011010011101010001010000110101110101111000110010101011010000000010110000010000010101101111000111110000111000001001011110110100100111010111111111001010001;
#1 $display("%b", po);
# 1  pi=207'b011010000001010101010101111101100010010011010010100110111100010101101111110011001100100110001001110101000000011010100011110000000000110011111001011110001001010100000001111000011100100001001001010101000110111;
#1 $display("%b", po);
# 1  pi=207'b010001100100101110000011111000110010011110011001010000010001100111101100001010101011011101100111100100101101110100001101100011010110101101100011110101111111101111011100011011111000000101111010011000011110000;
#1 $display("%b", po);
# 1  pi=207'b111111011101011111110101001111001010001000011111101111000011111000111110001011011100111010001110111101110011111010011000110110100011001001010011110100111000101011010011100111000010100100110001000010010101001;
#1 $display("%b", po);
# 1  pi=207'b101001110100011011110100011001101101011000011110010001101000001110000010000000011111011111001101110110011110011011111100111010101110100100010010001010000110101010101010111010001111110000111001000110001111111;
#1 $display("%b", po);
# 1  pi=207'b001000111101100111101101111100100101010100100010100011101110000010001100100100101101001101100100111001111011011010100000000011001001011001001010101011110100011100100000100011010100101011110011010010010010001;
#1 $display("%b", po);
# 1  pi=207'b011100111110100100100011111110011101011011011000001111110110110100111001010101110110001010100100110010111010111100010101000001101001011111101001000000111101101000100001100000000110111000101100000010001011010;
#1 $display("%b", po);
# 1  pi=207'b111001011101000111001001001110000111001001001101111110001101010011111111100100110101001001110111001001001001110100000010101001001011001100111111011101000001011101101110101110000111010001000101111001010000110;
#1 $display("%b", po);
# 1  pi=207'b111000001100000010100111100001101001011100110000000110011111101101001001101110010110100101110001100111001110111000110010011100100110101011010000111001111101111100111100000011111111011110001000001110001010101;
#1 $display("%b", po);
# 1  pi=207'b111110011000111110011011100011011110010000001000111010101111111101100111110100001111001001000111110101010000111001101100110101101011101100011010000101110011101011011110111110000111011011010001001110110011111;
#1 $display("%b", po);
# 1  pi=207'b011000001011111100000001100010010001010101101001010101111011110010110000000010010110101110001000100101110011001010111100011110000101010010110111101000011011111100111000010001100101110110101101111001111111111;
#1 $display("%b", po);
# 1  pi=207'b000100010010011011110110111110011101100101100011011001000000101000100010100010000011001100100010010011100111011011100111110101000001111001010101101011100011111000100101110000010010110100111010000111110000001;
#1 $display("%b", po);
# 1  pi=207'b010110110100010000010100110111001001101001111010100010010110001000010111011100000011100011010010011111111001100110110010000111110100000010010111101010000011111011001010111101100011101000001101010110001001001;
#1 $display("%b", po);
# 1  pi=207'b011010110001000100101100101011100111000101100011000100010110000100111100100100011000010110111101000110110000111111000000101110111111111110101000001111010001000101101010110000011001101110000111010101001111100;
#1 $display("%b", po);
# 1  pi=207'b011000100101100011111001000111001111001010101100001111110101111111111011100101001001101001110101001100001100101100101011001110010011101111101001000011001010100101010100111101010010000000011001001101000010001;
#1 $display("%b", po);
# 1  pi=207'b010110001010000100010000110001111111010000010011101101010100110101110110011000110011010011001011001011010001110001110000010111100110000011010010111110011000011011110111110100000010101000001110100101111101011;
#1 $display("%b", po);
# 1  pi=207'b000111011001010000000110010010001010110101001110000101010001001001110100100101100011110000111001000011100100010110110001110101000011011001101111010111010010001101010100010111001111100101000100101010100110001;
#1 $display("%b", po);
# 1  pi=207'b001010100000100100110101100000100111101000010110011000101000100010110000000100000011000010011001101001001010111111010000000001000011111000100111111000111011110010011010100110110010010000110000011100110110110;
#1 $display("%b", po);
# 1  pi=207'b011010010011100010111000111011110110110011010100101010101110111011000000100000011100001011100101000000111100101101011101110111100000000110000100111100001001101101000010110001000110101111010110000101110000101;
#1 $display("%b", po);
# 1  pi=207'b000111010110111000000101111001001101000111001001001001111111011001001110000110000100111001111110110100110111111011000011001010111000111011111101011001000000001011100110110011001110101010111010111001010110010;
#1 $display("%b", po);
# 1  pi=207'b001111001110100010111010010111100111010110011001100110100011101001011001100000111011010011110011110110110100001110001011011000011101100000001110011101110100110100000011111001010111111000101000011101110000111;
#1 $display("%b", po);
# 1  pi=207'b001101101101000111101111011001010111100100000100111111111011110100001001111000100110110111011010000000011000110001000000001011101011100001011100011111000001010111001101011011101100111100100100001110011010000;
#1 $display("%b", po);
# 1  pi=207'b001011000011100001011101111100111000111000101000101001010000100111011101011001011000101110000111110100000101010101111000001110010000011010110110101011101101100001101000100110110101111010010101000110110110101;
#1 $display("%b", po);
# 1  pi=207'b111101010100101101110100111101110011011011001110101101011011011101101100111011100101000100110100001000000101001011110101010100001110000101111010110011000001010101000010100111001110001000000111001100110100001;
#1 $display("%b", po);
# 1  pi=207'b111001001010110110000101001100111101110110101000111101110111000111110100111110101101010111011110100010010011101010000011001101000101111111011011010111110011001000001010010010110011011011010001101101110101110;
#1 $display("%b", po);
# 1  pi=207'b111100010100001010001111100001101010010000110110001110110000100011101000000101000011001010100000000100111011101000100001111000011001011101000000110010010010101101110011111000001100101111110100110110110001101;
#1 $display("%b", po);
# 1  pi=207'b100110100001101101100111001110000001000110001101111110010100000001101001111100110111111111100111010100100110110011011000111101001001010101100101100000010110010100010111000101100010100111011001111011011101001;
#1 $display("%b", po);
# 1  pi=207'b010100100011110101000011000100110010011101010100100111111111101100111101011010111110110111101010000111111110000011101111111001110101011000010111100101011000011001100011011100010011001100011001111000000000110;
#1 $display("%b", po);
# 1  pi=207'b110000001001010010010101100000111100110110101101110101100001000001011000000001100111000011100010000100100100100110101110101110000010010110010110111101101111010000110110001100100111111001011011100100110110111;
#1 $display("%b", po);
# 1  pi=207'b001100001001011100011110110011100111110000010101001101000101000011101101011100010110001010100001101110101011000100001000000011100101001110100000001011100101110010011000101110110011010101000001011110001010101;
#1 $display("%b", po);
# 1  pi=207'b001110110011110000111000010001000000101110100101011100001011011011000010011010001111100100001010011110100000001101101101101010011011100010000101111110010110010101000001110100010011000011100110101000010001110;
#1 $display("%b", po);
# 1  pi=207'b010010111100100101100100010111001110001111101001110101111010100001100010011010100000110011110101011101101010110101011000101011111000110100100101111001001011101110111100001011000101001110101101011101101001011;
#1 $display("%b", po);
# 1  pi=207'b011010111101010111010111010110100100110011001101110000110100101000101010101001010010101001100011000111110100100000001110011010010011111000001101111001011000111001101000100100111110010110101110011000101001001;
#1 $display("%b", po);
# 1  pi=207'b011010011110001011000111001011010011010100000011010100110101110001001011000110111110011010010100111101111110111111001111000000110101110011000111001010011010010101110111111001111000110111010100001110100101001;
#1 $display("%b", po);
# 1  pi=207'b011011001101010001110000100011100100011010101111000111010110100001100111011101001011101101010100101100000010011100101001001101100010100010110000100010001010000010100011010100100010001100100001001101110011100;
#1 $display("%b", po);
# 1  pi=207'b011010100101101010001110001101111111100101010110101111001101111000010101101010100010110101101110111011110001110000110110011111111000001111100000010101110010011100100001101111100110111010001000110110001110111;
#1 $display("%b", po);
# 1  pi=207'b010101011110100101001100111011111100011110101010100110010011101111110000111111011100000000010101111011110111001110000100100011010000100011000101101011101111000110011001010001010001101010010011111110111000001;
#1 $display("%b", po);
# 1  pi=207'b100100001011101010001110010010001011011011111100100001110111110111111011110010111100111000010111010110100001110101001101001111101111101011101111111110101101110011100000101111110010000100111000100110111011101;
#1 $display("%b", po);
# 1  pi=207'b010001111100010111100001001010111000010101000111100010001011101010011100011101000111111000000001001110010001011101010000110000010110001101010001111011110101010010000001101111111010010010000000101100111011011;
#1 $display("%b", po);
# 1  pi=207'b110011000010100110100011011000101011101100010110110110101010101100111011101011000110011111111101100110001011011010100101100000010000110011110111011100000001101000011110000111110110000110111011101001111011011;
#1 $display("%b", po);
# 1  pi=207'b011001011111010010001110000011100101011110101100001000100101001011111101100110001001000110001010110011100000101110101011000001101101101111101010011001111000111010100101011111010010111011000000000111111001111;
#1 $display("%b", po);
# 1  pi=207'b000011100101100000101010010011000010000110001000000110001010110000101110011101000010001001010101110101010101010111011011000011111100101001001000010110110110001111001001100000000110011011111000110011100100111;
#1 $display("%b", po);
# 1  pi=207'b010000001111001110110101101100000001001010000010000111100001100011001011100110110101110010000000000001000000000000110010100010000010011000110111111101111100100101001010101000000000010110001110110100000110010;
#1 $display("%b", po);
# 1  pi=207'b011000000100001011001011110111110001010001011010010101111100010000110111111010011100100111010000001100001011001110011001011111111001100010110111111001110111011111010100100010000111011001001100001101011101011;
#1 $display("%b", po);
# 1  pi=207'b110100100001000100001011101010100000101101100111111001110010110100001011101101110100001110110000000101011111000001001000011111000110110111111110011101000010101111010000001110111010100010011110001111111000111;
#1 $display("%b", po);
# 1  pi=207'b010001000000111100001100100110100110110001100101110101101110010110100011011100101011110101111010001011111101111001010110001010011100110100001010101100000100101111001110111110010001100000000011010001011100010;
#1 $display("%b", po);
# 1  pi=207'b001110010000111010011011110110110100110011111101001101101111100010101101101101110101100110101101100000011111100011001000111100000110111010000110110001111000011000101010001010101000100001001000101101011100010;
#1 $display("%b", po);
# 1  pi=207'b010011110001110010000010011100001110101111110111111010110010101011001110110011010101010101001100001110010000010011001100010100110110010000000100111101110100001111011001011101000110110110010111100010111110100;
#1 $display("%b", po);
# 1  pi=207'b011010001111010010110111100010110110110110000010001100011111011111110100101000100001110111101101011111111110000111001011110001111100000010111110100101000000000111010010011010111001010101010100101100010111111;
#1 $display("%b", po);
# 1  pi=207'b011100100101101111011011011101101101011001011100101001101110001100001000001111010010110011100000111001011100100011101001111110010101110101110000100110000000110010000111000001100010011101101001001001110100011;
#1 $display("%b", po);
# 1  pi=207'b101011110111110011011111110110001010000001011011011001001111011000011011011101001011011100100001111111000011101110000011110101100001110111010000111001011111110111100110100111111001001000000111110100101110010;
#1 $display("%b", po);
# 1  pi=207'b110111110100011110010111110011101110011110101110100011000000100010010010010111001110001010100111101100100110011000011110110000010111010000010010001111100110011011001101100110000101001000001010100110101111010;
#1 $display("%b", po);
# 1  pi=207'b010001010001110111000101101011110001110000100010101101100101101110110010110010000100101111010111010110100000001001010011110111001110001110011101010110010110111111011001101111011010000001101001011100110000000;
#1 $display("%b", po);
# 1  pi=207'b000101111100110000011111001110100001110000001111111011110110111110000000000101010110100100001111011100000101000001000010110100000000111001100001110010010110100100111101011110010010101110000100110101010110111;
#1 $display("%b", po);
# 1  pi=207'b000001011101110011111010110111000000111000001110010110110000001001100111010111000001110110011100000010010000110001001001001101001101000001101011110001000010101100000011101001110001101110001101011111100101100;
#1 $display("%b", po);
# 1  pi=207'b010110010010100110000001011110001000011110011010011000001110111011001001000111100001111001100100101101100001011100111101000001111100000111010110010010010001000100110011000100111011000011110110000010010000000;
#1 $display("%b", po);
# 1  pi=207'b100111011110001110100100101011110010000001001011110010100011010101111100110011110100010110011011110000101111000111110001000100000000000111101101001011000110101100010101101110100010101100000100001101100110001;
#1 $display("%b", po);
# 1  pi=207'b010001101110101000101000101000001100001100100111010010110001001100010010001011000011011011001111111100111000001011011101011000101000100001110011111111011100001110011111111100000100100101110001111101010000011;
#1 $display("%b", po);
# 1  pi=207'b111101111101010100110011111010100001001100001111101000111001000101000111011011001001100010111101110111001100101111010001000100000011111001011101111000110100101110100101001101111100010110001001101111010010100;
#1 $display("%b", po);
# 1  pi=207'b111001101111010001100001110001000100111000110111100111011111001101111101011001001011011101101010011100100111011011110011111011011001110110101000110111100111010111100011001101111011010110000100110000110100110;
#1 $display("%b", po);
# 1  pi=207'b010110100101100001111000110001101110001100100001001111110011111111010001001110000010001101001011110110110111001010101110010101000111100110010001001001000011110000010000010010110111110000110101100010110111101;
#1 $display("%b", po);
# 1  pi=207'b010011001010101101110001001101101011000101111010010000110100110011001101101110011111111111101000010010011011011110011010100010101000110110110100000001110011001011100110110000001101100111001001111010101111010;
#1 $display("%b", po);
# 1  pi=207'b111001000110010010110001101001100000010000111001111100101000011110001011001010010100000111101011111010101001100101100110011111000000101011011001011001010111010110110000100110010100000110000101101011110000100;
#1 $display("%b", po);
# 1  pi=207'b010100101011011010011011111101011101011110001010111011111000010011111001010000011010010101101101100111111010100111011001110110001000011011101110100010100001100000000000000001100011001001000100000100011011001;
#1 $display("%b", po);
# 1  pi=207'b101010100111000101100110110001010100000001101100001111101000011010011011001011011111011011111010000110111011110100111001100100010111010101101100010110001111111010110111111011000001010000001001101101101110011;
#1 $display("%b", po);
# 1  pi=207'b101011011000111010101111010001100011000001100110100011110100100101011100011001110001010110110111100110010100011111101100110000100111111000110111110000000101111111110010100101011111110010111010011011010100101;
#1 $display("%b", po);
# 1  pi=207'b101001110011001001111100100100101011011011010011001100111110001111010100101100011011001111110011110000110001011101011010110011000100011000001011010111001010011000100001111100000110100010100000110011000101101;
#1 $display("%b", po);
# 1  pi=207'b111000110011100000000100111111100000111110110000000011000111001000010000100110101001101110001111100100110101000010100000000111000011011101101111000110100010011010101010101000100110110010010110011000000111111;
#1 $display("%b", po);
# 1  pi=207'b011110010000101101100000101010100111100000011111010001001101100001000001011010011101100011000011000110110000011010100111110101100010111100100010111010010111101110001101110011000110100001001011001001010010110;
#1 $display("%b", po);
# 1  pi=207'b000100001110010110010000010110000011110001111111011110011001111110101001011110001011111101001011011111001011100011011000011011001011100000011001111011110011011100100010011101010101010100110011110011101100000;
#1 $display("%b", po);
# 1  pi=207'b101101100000001111011010001010101101010000000101011010010011000101011001111110001010010111010111000001011111100101111111110011001010010010011001101101011011100010000011010101000010011001100100001011010010110;
#1 $display("%b", po);
# 1  pi=207'b110000010010011000111100100101100100001011001101001010111001000111101111001000011110000101110111100100011110001101101100101010110101111100000111110000000100110001111101010110000010111100110000111011000010000;
#1 $display("%b", po);
# 1  pi=207'b100110011111110110101010110111110011001100101100101010101010101010010010000001001101110101110010100100011101100011111010110001000111101011100111001101111011001000010001101001100001100000001110110101111101001;
#1 $display("%b", po);
# 1  pi=207'b110100100010001001001100001101011011011010100110111001110111000111110111111100010101001011100111000100000101010101011111100011000100100110111001001110000100100100111100100101110110011011010110100010101110101;
#1 $display("%b", po);
# 1  pi=207'b010101111010100100010101010110110110011011110100101111111101111111111101000101001000100111100100011110100100001101100000111000000100001000101100000100011100010011101000000011001010000110000111001111110001111;
#1 $display("%b", po);
# 1  pi=207'b110011001100011001010011101010101010101101000000010100010000100000100000001011011100100010011101100100001100111100010011110101001100010110000111010100010101101110100011101010100011010001000100001111011000101;
#1 $display("%b", po);
# 1  pi=207'b011101000100100010101010101011010111111011111110000010001111101011110101111001111001111001000010110111001100100001101110001010111011011110110101101011111000101011110011111001111010101011110001111100100000001;
#1 $display("%b", po);
# 1  pi=207'b110010001000011100111001000011111111101000010100100001110111000100111011100111001000011000010111010101001101000100011010101111011100010000111001100111101111100011011001110010111010000101011010101110101111101;
#1 $display("%b", po);
# 1  pi=207'b001011010111000001110010101110001010010111100001101110100101011101100011100110111010010001001100010110010110001111010000110110001000111100111110011010000101111000110111000111110111001010110111101110110000010;
#1 $display("%b", po);
# 1  pi=207'b010000111000001000000110110000100011101100000000100110111111100000001010100010101000101011110001111101110010100100011110001011110111101100010100111011110010011001011000000010111101100101101100001101011110100;
#1 $display("%b", po);
# 1  pi=207'b100110011000111110100011111011010100100100001101011001110001010001111001110000001001100100110110011111010011101010001010001001111011101111110110000111101101011011101100100011111101110010101011111010000101001;
#1 $display("%b", po);
# 1  pi=207'b000101001111011111011011011000000101010110010000010010001010110011000101100101110101010010011100000100101111110000110100100000101011110010000100000111011000000111001001101110100001100100110010010101110111010;
#1 $display("%b", po);
# 1  pi=207'b001011001101010000110101001111100000000010011001111100011111000010000001001110110011000000010101001111010101000100111111011000100101111110111000111110000000001101101101000011001000110010000011101001101001001;
#1 $display("%b", po);
# 1  pi=207'b110000111000000111001100101101000111100010110101011011001100011100111110100111010000000111001100011010100111111000001000101100010111110010010101101001010010010111101100000010011011011101111101100110101111110;
#1 $display("%b", po);
# 1  pi=207'b000110011101000011011001011101001011111111011001101101110010101110010100011010100111010001101011010101001001001011001000011110101000101001001000000001000010110111010010111001100111110010101001001100111101011;
#1 $display("%b", po);
# 1  pi=207'b011001011110000001110001101011111011010000101110000001011110011010010111010001111011100000110110110010001111100101111101101110110011100111101111100001100101100010111011101000101001110011101001001010100011110;
#1 $display("%b", po);
# 1  pi=207'b010101001010000010100110110110011111011001000100111100001100111000110001110001000100100110111110001101000010011100011000110000100110111000011100011101111110101111100010111111101111010001001110100111101011101;
#1 $display("%b", po);
# 1  pi=207'b101010010110111111100101111101100000011111001111101010101110100111001110010101011100110101110010010101111101000101000100100011000011110000101111010011011101111100101011111101000010000101111011111101100100011;
#1 $display("%b", po);
# 1  pi=207'b001010010001111010011100010111100111110010001010011011100110110101001101000101000100000011001010001101101000000011000110001000011000010000010111110101011111001111001001100000010001011110000011000001110001100;
#1 $display("%b", po);
# 1  pi=207'b100111110100000011000010110011011100010001111011011101010001100100110010111100101101110000000001111100110011010100011011110100011101101100001001011001000010100100100000011111010110111111010101101000110001010;
#1 $display("%b", po);
# 1  pi=207'b100111000101010101111111110011011001011010111001000101000001000010001000111001110111010001111101111011001101000110001101001011110000000111110100000100100100000110100000101101101101100011101101000010101010110;
#1 $display("%b", po);
# 1  pi=207'b000001001111000011000110110011011000000110101000111011001000010100011101111110101011100011010001100011110110010100110111101101010100100110000101110000000010111110110110010110101000000001100010110101000010111;
#1 $display("%b", po);
# 1  pi=207'b000000100100110110111011111111110000110011110011010010010100100010110101010101010010101010110000111010110011011101101001101110101001111001010110110010111011010011011100010000010101001111000011110000001100000;
#1 $display("%b", po);
# 1  pi=207'b000000001100101100111010000100011101011010101011010110010111010101011010010110000000000011011001100001001100110001011011010011110111111000000000101101001111011111010110011111110011111011001111011010110111111;
#1 $display("%b", po);
# 1  pi=207'b000101001010101110011110011001000101101101010110100001001100100100101010100101100001010100000000111011000101010010000011010010001101110010011011101010101010011001010100011001000001111100111000000101011111010;
#1 $display("%b", po);
# 1  pi=207'b010001010001111101100010101000000110010101101100100111011000001001001100011111101011010110110011011101111100111001101000100011100110011111101100001111000111111010001111001001001111111010000111001101010110111;
#1 $display("%b", po);
# 1  pi=207'b101011011101110001111100111110110010000000001001101110000001110100001100101110011011010110010001110101110111010111001100101101011011101101110001011010000101111011100001110101001101101100010100011101011000010;
#1 $display("%b", po);
# 1  pi=207'b011110010110000010110011000011001000100000001100010101010000010011001010101011011100010111001110111000110101111110011001000000010110000110111000000001000011111001110101001010010101010011001010011001011001100;
#1 $display("%b", po);
# 1  pi=207'b000101010010011001101001101100011001101110100100101101111011100011001000000010110010001101011000011101110000111001001110101111001011101000110110101010001101111001000001110110110100110011101110101101001001111;
#1 $display("%b", po);
# 1  pi=207'b001111001101111001110010111001101100011011101100000001011011010110000011010101010000010001000000111010000010001000111111111011111100010000110110110001111111110111100000000010001000001100100111110000010111010;
#1 $display("%b", po);
# 1  pi=207'b010010101010101100111101000010000000000101101101101011011010100110111011000111100000000101011111110101100000111100111100010100001010011000000101000110101000000110101100001000010000111110000101110111011001011;
#1 $display("%b", po);
# 1  pi=207'b100010110100011000010010001011011011011100101110001101110011001111101010101011111001111001000100101010111101101010011000000101000111101010000001111110101001011010111111000010101110111110011001100101110110011;
#1 $display("%b", po);
# 1  pi=207'b100001101100011011110100101001010001101110100101100011110000000101101010101001101000101111110101110111001110011000010010111001100010001100111101101010011101010010101000010001011100111001101111110100100001101;
#1 $display("%b", po);
# 1  pi=207'b001011100100010110101110110011100110011100001001001000100001110011110101110100101001111000000110110101010100010001111011101001100011110100100001100001111001100101110101011000100101110111110110111110100110110;
#1 $display("%b", po);
# 1  pi=207'b110110100100001011110110001100010000011100100110100001001111000011101001110001001010011110000000111010000001110010100001101001110110010011010100010111010111100111001011000001001111101011101000000010011001110;
#1 $display("%b", po);
# 1  pi=207'b100100011001011000010111001000100000111111001111111011111001001010010001011101010001100011101110111001101110011111000110001000010100001111111000110101110011010110101111100110010100010010111010100010101110010;
#1 $display("%b", po);
# 1  pi=207'b101111100010110011111010110010101101101110101010000111101000011011010111001111011100101000011000101100010010110011000110010001011110010011011111111000001000000101100101111101101001100110100100111000111001110;
#1 $display("%b", po);
# 1  pi=207'b001100110110101000001101000001001000011110101001000100101111000111001111111000011110011010001010101101111001111111101111110111001111001011011011100011111011010011110011110111010111011000010110110110010001100;
#1 $display("%b", po);
# 1  pi=207'b010011011110101010010100000100111011000101001101111101111000110101101100000100101111101111001111001101110010110011100111001000010000011001000001011000101000110000110100011101101111111110110011100010000011111;
#1 $display("%b", po);
# 1  pi=207'b000111101110101100101010010110100111001101001010001100011010101000110100010011110110011010001011111000111111100001001011001000100101111110010110110100010010001111101111110000000111011100010010010010000001110;
#1 $display("%b", po);
# 1  pi=207'b111101011010101111101111101100101100010000010111100011110101100110011011110001100011110001000000100110000010101011110010100011000010111011011001001110100001101001011110101101010001010110101000110101010111101;
#1 $display("%b", po);
# 1  pi=207'b011010110010101010111100110011001111011100000010010001110101111001001011001110110111011011101100101111110001111011010011100111101011010110100100000001111010000000000110111101000001010010010000001011010100010;
#1 $display("%b", po);
# 1  pi=207'b100001011010011100001000000001111010101000000110001001101001011110000011111000101100000100011110001000000010000100000100100100010010110100001010101111100101001000011100100110100011010010101100011000010000100;
#1 $display("%b", po);
# 1  pi=207'b000001100001001111101100000111010111000011100110101010000111111100011101101110110000100001100011101100011111010111111111010000111000000101111111011101111101010011010010101111101100010111100000110111101100011;
#1 $display("%b", po);
# 1  pi=207'b010100110100000010011011100010110101101101010010000110001000101011111001111010101000000110010101100000011010000011000100101000000111011010011011000110110000000110011101001100101010010101000001001110000011000;
#1 $display("%b", po);
# 1  pi=207'b011010001100001111101001101011101111001001001100001100011000011101101100011010010100110100001111101101101100101011100101101110010101110001011010101100100001001001010111111000101101111111100001000010111101110;
#1 $display("%b", po);
# 1  pi=207'b000011100111000101111000100101010011011001000110001011110101110101110101001000011000000100010111001011100000101110100100111010110011110001110010100001111110101101110100001011000010000110010100101001110100010;
#1 $display("%b", po);
# 1  pi=207'b000101111011001101111000010001100110011110101101111000100110001111011010001011010110110001110101111001100110101000010101001001101100101100001010010110100101101011010111100100000110101010101101001100001100011;
#1 $display("%b", po);
# 1  pi=207'b000100100100001110011000101000010110110100111011100100100001111110101000011110111010101000000101100011111000100001010010000001011010000011000010101001110101110000100001000011110011100111111101100100010010010;
#1 $display("%b", po);
# 1  pi=207'b000010000010110010001110010010110101010010100101111000010101110001100001001011001001001101000110000111110111001101111001100010000111010010001001011100001100011100111000000010110100001000110001010111010001010;
#1 $display("%b", po);
# 1  pi=207'b011111000000001100011111110100001101111110010100010001000110100000101100101011111111100010010000111111000110110001100001010110110010101011110001000001100110100010001000100010001111011101000001001000101010100;
#1 $display("%b", po);
# 1  pi=207'b001100111010100111011101011001010011010001110110000110010110100010101001111100100010111000110110001101010011011010111110100110101010100110100100101001011011111001100001010101100101110010111110011001101111100;
#1 $display("%b", po);
# 1  pi=207'b110110001010010011100101101100101011001011101011111010010010100111011011111000110001000010101010000101100001111000001100011101110101101101110110101011001011001101000110110101101110100110101001001001001100111;
#1 $display("%b", po);
# 1  pi=207'b101011001000101111110000001000101011000011010100100000100110110001110001011110011001110011110001110100101110000000111110010001110110100110000111000011010110000010010100110001101100000010000111000100110010111;
#1 $display("%b", po);
# 1  pi=207'b010101110000101100101011100010101100000011011101000110000111001111000010000111100001101011100110010011111011000011101011000001110101100111000111100110000100001100100100100110010011101011101110010001111001100;
#1 $display("%b", po);
# 1  pi=207'b100101100011101011111110110110110111100010101011011111000000011011001000101111111001110101010111101010100100111001000111100000011100011111000100000101011010101000110100011100110001001001101101101111101010111;
#1 $display("%b", po);
# 1  pi=207'b001111110101011110000011100101010011111110010010111110110011010111101110001110010010100110001010000101000110001111111001011100001101011010111110010100011101000111011001101101101110001011001101101101001010010;
#1 $display("%b", po);
# 1  pi=207'b111011101111100010001001100101101000101110010100111010100001110000111010000010100100111001000100010110011000000010100001111111110101011111111100000110010101100111001110010100110001101010111011101001010111011;
#1 $display("%b", po);
# 1  pi=207'b000111001100001001100101111001111010011111010000111111011111010000010101011001110001100010001011010000100010100011000000011100111010110000001011000000000110100001000001101101101011100111001000011101100111001;
#1 $display("%b", po);
# 1  pi=207'b010101101100100000000111110111010001001000010101001110110010001110110101001110100101010101101110011000010101011010111110110100101011101001001100000011001111111001010111001011010001110010111011010001011110000;
#1 $display("%b", po);
# 1  pi=207'b000001001100100000011110001101010100011111101010001000100111110010101010011111110110101001010010101110001001110101001110000011101010011100010100101110111001000000101111111111110100010101000101000010000101110;
#1 $display("%b", po);
# 1  pi=207'b000000100101011111110110100011110100100100100111001110011110100100000101100101001010101101000110000101110100111110110100011001010001000100111101011001011100101111010100011000001010011111101000100010011010000;
#1 $display("%b", po);
# 1  pi=207'b010001100001001111100110101111010010100000101011010100001100111100101001010101111101001010010000001101111011000000110010100111110110010111110010000011000101001101010101000111010111000111010110000001001000100;
#1 $display("%b", po);
# 1  pi=207'b011011010100010111111111001101011100001110110101100010001000110010110000101011011010001101011111010011010011101111001001100110010110010001101000101101000010010110111101101101011000001111010100101101111110010;
#1 $display("%b", po);
# 1  pi=207'b000111101101000001011110001000111000000110101011001010100001100011000100111100000011101110011001100100010000000000001111111001100000011111010000100110011011100001101100001110100111001001000011110110111001110;
#1 $display("%b", po);
# 1  pi=207'b100011000101000000001011101011000101100000101000010000110001001011000010111000000101111111111001111100001111001101001001101010010000110001100001000100111010011101001100011011100100001010100101001100011001011;
#1 $display("%b", po);
# 1  pi=207'b011001110010011101000011010000100010110110010110011000001011111100111000001001000011110001011110000001010011111001010010100000110111110011001001101111111010010001100111101010010110100011111000010100000110110;
#1 $display("%b", po);
# 1  pi=207'b011101011110011100110010010110011100001000010000101110110010010000110111001101010010001001110000111110101011111011101110011100001010101001010100010111110101010100100111000111101100011100111111101101001100000;
#1 $display("%b", po);
# 1  pi=207'b110101000100011100011100000011000111001101100001001101111100000011000011100000010011011011011110110001010001111001011100111101110010011001011111000100111111110111110010000000001010011000110110000111011101101;
#1 $display("%b", po);
# 1  pi=207'b110111010110010100011110001011001010101101000010011001011001011110011000111110010010101110011101110111010111001111001011101111011011000101011000111011110101011001101111000010110101000111101011011000100000101;
#1 $display("%b", po);
# 1  pi=207'b110100010000111011111011110000010001101111001111010111000011111000110100110001111000010100001000111110011100100000011011000001011000111011010110110100101111001001111010110001001110101110001010010001011010101;
#1 $display("%b", po);
# 1  pi=207'b011111001011010001110100110111000110010110110011011111111111101100110100101100100101110110000011101110001000010101100111110110100010010011001100000010101011101010000010001010000000001000111011000111001010001;
#1 $display("%b", po);
# 1  pi=207'b110010100110010010000011000001110011001101111110100001111100000000111001001011111000101001011101101011101100000010110101110101100000000000011001000101001110100100100110000110001000011000000111011011001111011;
#1 $display("%b", po);
# 1  pi=207'b111110110100000111100110110111110101001100011101011000001111010000010000100100100101110110001000000010011011110000101110010101000010011111000111111110111001110001100110000100011100001111100011000100111001010;
#1 $display("%b", po);
# 1  pi=207'b011111110101010111011011100001010001010100101000010011111001110000111011101010101111000100011111100100101111111110101000010111011110000101010011001111001101011100110111101001000011010001001001010100010100110;
#1 $display("%b", po);
# 1  pi=207'b101010111000001111110111100100000100010110001111010000001011011001001011110111111001111111001101010000100010000100001111111010100011101111001011000011110000111000101111101110100001001110100100011011000011011;
#1 $display("%b", po);
# 1  pi=207'b010111100001111110101110001111110001110100011101110000011100110010011101010101011010100011000011000010111110000011101011110000001101011111001010111100111011000001111110111111001000111010010000000000101110110;
#1 $display("%b", po);
# 1  pi=207'b101110101101110000001111011110111110110101111110001011000111110101000101100110100010111111011101011100101100000010101011000000010100011111101111111100011101000001000101100000100101001101011101111110011100011;
#1 $display("%b", po);
# 1  pi=207'b101000000010001101100000100110111001100010100001101100110100111111001101010111000000010000100100011100110101000110100011101100110010001111101101111101100010001100001111111101001100000001001010011011001100011;
#1 $display("%b", po);
# 1  pi=207'b100000100101111001111010111001111010111001101001001010110110100110111001010111001111000000100001101100001011011100000101011011100110100000101100111100001111001111100001101010100010110110100110010000011110001;
#1 $display("%b", po);
# 1  pi=207'b001111000000100011101111000001011100101111001011011111111110001001101000001111100000011001101000010111101100001001111000110000001111110010000010001011010010011011101110111010010000101101011111101010101111111;
#1 $display("%b", po);
# 1  pi=207'b011001101100011100010100110001011010011010010110000100111101001100000000100110111011000100010001010011001000001000100010000001011100011000001101100010110001111111000101111111101000100100101111101000000001101;
#1 $display("%b", po);
# 1  pi=207'b111111000100001011010111110011101011001100111011110110011100110111111100000001010100101001011110101010101001001000101110000110001001100010010010001000000010100010010101011000000000101011111000011111111000010;
#1 $display("%b", po);
# 1  pi=207'b110000000010110111011101101111110010011110001001000010110001111100101010001110111001011100100101000000110101000000011111111001001111010011000101101100000001001101100010011010110101110001000001100110010111101;
#1 $display("%b", po);
# 1  pi=207'b101001000001100010001000100010100001001110010110110100010111001110011000110110101001100001011001110110100001110111100100100010111111010001100101111100110110001011100100010001111000111000100111001010010101111;
#1 $display("%b", po);
# 1  pi=207'b001111001101111100000011011001010001010111110110101110000101111110010111101111011100000110000111000101010100110101101100000110011100010001000111101110101010101110000010011111000011101101101101101011011101001;
#1 $display("%b", po);
# 1  pi=207'b100001011000110011111001001000010000011010101010011100100001000000101001111011000111000111001011001000010010010001110001000111111010000001111000010110010110001101111100001111101101100011110010111000000001111;
#1 $display("%b", po);
# 1  pi=207'b111000000010000101101100111000000110100000101000001011000001111111100010100010010111101101101000010010110011100001110001011011110000100000110101001000000101011100010001010000100101100011000110001010101110011;
#1 $display("%b", po);
# 1  pi=207'b011111010111010011110110111011100110111101101011100001000101010111010111100011100000011111001101101001101001101011110001001101111100101111011101110001001000101000001101111101110101001101001011111111110101100;
#1 $display("%b", po);
# 1  pi=207'b101111001110111110101001000110010100001010010001100101000011010010110111101011111000110010010110110011010000000101011111010000000011011101010100001010000001010011100010100001110110100010000111001001010000011;
#1 $display("%b", po);
# 1  pi=207'b100111000001000000000001101010111101111001011010001110011000110111101111000011001001111010111111000000010110011101001111101011001101010100111100000110011100011011110100011010101000111101011001110101011111110;
#1 $display("%b", po);
# 1  pi=207'b001000011011001001010000011000001011000100010111001111110110111100110110000100001011110010111111101100011111111001101011011111010011111011111011010011111010001111100010010100011111001111111110101111000101100;
#1 $display("%b", po);
# 1  pi=207'b111101101101010000010101111000001000100110101000100111110101100110001100001111111010001001010000010100101000111010101100100101100001001101011101010001101111001110000111010001010111010100110101110011101110001;
#1 $display("%b", po);
# 1  pi=207'b100101000111000011111110011010011000110001111011110101011101001111011100010000010001100110001111001001001011001110001011000010111100010110000011111011111000110100100100000111111100011101111000111000001110111;
#1 $display("%b", po);
# 1  pi=207'b101001011011111100000011000000011111011111110101111011011110000101110010001001100001001000111001101100011000100011010110100111010011000011001111010110100010111100001111001110110000001001110011000010111100101;
#1 $display("%b", po);
# 1  pi=207'b010110010010010000011011001100111000110111110001011101010010011110100100011010111010111011101100100001011101001000010111000000100100111010111001100011001100100010111010001110100010100110000011010111101111100;
#1 $display("%b", po);
# 1  pi=207'b011100010011110101100110011101101011110001110011011101001011111001010010001000000011100000110011100000010001001001001001010010110011100011011000000101001000000101110101011111010011001001101110111010000100110;
#1 $display("%b", po);
# 1  pi=207'b111111101111100110100111101011000100010011001111110001110100101011010001110101100110101010110011111111110011110000101001001011001111110000111101001001111100100010011111010001111010110101011110001111100000000;
#1 $display("%b", po);
# 1  pi=207'b100011111101010011000001100110110110101011000001001100111100100101110001110000111110000000011010100000010000111100110000000110000000101110111011000101010010100001011001000110011101011010011011010010100001111;
#1 $display("%b", po);
# 1  pi=207'b101000000010011110110011010010100101011110011101000011001001110001111000111101110011000100000000011001110111101001011000111110110111010001000100001011111001101011011100101010111000001100101010110111101100000;
#1 $display("%b", po);
# 1  pi=207'b010000111101101011011011011101000011100101010010011001011110111011101000001101110000111010000110010000010000111010011111011101110100111101011010011100010110111001011111100101001001101101011111010101000001101;
#1 $display("%b", po);
# 1  pi=207'b101010101001100111001100001100111000110001011010100100111010001010101011110101010011000001001111011111101010101011110010000010100101100000110101101011111010010110010010100000110100101100101010111011111111101;
#1 $display("%b", po);
# 1  pi=207'b011100100010100111000101111000111000010000010010011001100101111011000010010100111010101111001001100100101111011111101001001101000101101110111010011110110110011011010001111101010111000111000001001111100001000;
#1 $display("%b", po);
# 1  pi=207'b001110100010011000010101101110001110000011101101010001011110010010010001001101001101011110001010110000110011001001001011000000001010010010001000100010100000110101110101111010111001101110001110011110101100100;
#1 $display("%b", po);
# 1  pi=207'b100111010010100001101000111000011001110111000110011100001001011111001100011100110101010100100010001110010100000110001100001111111000011000001010101100011111011000100000100101101010011101101111101111001101111;
#1 $display("%b", po);
# 1  pi=207'b111010111010100110101110101110110100001011011000101010100001111011000010100001110101010001111001100000001011001110001011001111000011000000100110110001100100010111101011111000101001001011101010110000101011101;
#1 $display("%b", po);
# 1  pi=207'b010000101011110000100001010011100001100010111000011010101011101111010110110100001100110001111110011110101011000101011001100101110011001111111110010011011110101000110100010101010101001101111111110111101000101;
#1 $display("%b", po);
# 1  pi=207'b011010100011111011111101111001110100011110010110001010101101001011101110010011000100110101001110001011111000111000110110001011111011001010010111000010101110111110111101010001001011000110110011010110111001111;
#1 $display("%b", po);
# 1  pi=207'b010001010011111001110010111000111110101001010010101100011100110011111001101000001011000100011100110011111100100110111101010101111100000111001000100010100011011011011100000000111111100001010101101110101011111;
#1 $display("%b", po);
# 1  pi=207'b000110010111110111011110100011101000100011001001010100111110111100111001110000101010101011100001111000100000010110101000011010111110001010101010100100000011111001011111100110101110101000101100011001111101110;
#1 $display("%b", po);
# 1  pi=207'b100011011001011100111001010111101000001100011101010110011110011000110101001001110001001100010100111000011110101111110010001011111111101110001111100111000101011111100000111010010100000111010001011010110110010;
#1 $display("%b", po);
# 1  pi=207'b000000011110001010011000011001011110011001001000001001001100111101111010111011010110110010110011001100010011100101100000010010111011100111011111100011010100000011110110001100011001101001001001011110111100110;
#1 $display("%b", po);
# 1  pi=207'b100110010111110110111001101111101001000100000101000001011001001000010110011111100101001010100000111111010111110000000111100011110100000111000010100011110101001011101011010110001100010001111101001101111100100;
#1 $display("%b", po);
# 1  pi=207'b100011111100011010101001101100000010010101111111101110100100011011111111001101111100000001011100110011100110110000000100101110101010011010101111010100101100100000100110010101100010100011101110101101110111110;
#1 $display("%b", po);
# 1  pi=207'b101010110011101101100001101101100101011110110000001001111100001101001110010110001011101101101010000101011100100000110100101010011110100110011100100000010011100100100000011110110011100110101110001110010000000;
#1 $display("%b", po);
# 1  pi=207'b001010101011100010110000111101000001000011101111110010001010010101110101010110111001101010110110100001000111001100010110010001111011100101010010010111111000101010010000001110110011011111010110100101011001001;
#1 $display("%b", po);
# 1  pi=207'b011111101111100011110100001001011010101110111010010011100100100010111111001001000000100001010111101010000010101110000111000100010110011000101001110000100100010011111001111000011111001111111100101011110011101;
#1 $display("%b", po);
# 1  pi=207'b110101010000110000100111111100011110000110011110101011011101100000110010110011110101111011110011100000110110111100101010111000101101100101100111101110011100100000011110000000101110100111000000111101011100000;
#1 $display("%b", po);
# 1  pi=207'b111100000011111001011100111001101101100101111001100001000010100110101000011101000001100101011101000011000100110001001110100000101000000000101001101000011100001110010001010001110011101011011111001110110100000;
#1 $display("%b", po);
# 1  pi=207'b110100110100100100000100111101101011011100110001001111001001011100110000111001010001100001000011100111111000111011101101001011011110100101011000011110001001101010001010000001000100111001011111001100101100101;
#1 $display("%b", po);
# 1  pi=207'b010111000100011111001001111111010001010010010101001011101000000011101101010010111000110100000100010111010001000001100010011010010110010010101010100001100111010011000111010011101010111010100011000101111100111;
#1 $display("%b", po);
# 1  pi=207'b000101110010000100101011010101100000111001001001010011101010000110001110000100000101001001110100100100100011010101010010001101101110101001010101001110101000000000001011010000000110000110001010000111110000111;
#1 $display("%b", po);
# 1  pi=207'b101101001010100110110111000000110101100101000011010101010011100111000010001010000101001001000100100011100100110100100010110010010011100000101110011101101111110111001001110110101110010100000011011111000010101;
#1 $display("%b", po);
# 1  pi=207'b001001100011110010011010100111011100111000011011001100101001110111110001010100111100111010110011010010101010011110111001000111000111000100011001010111010011000011001010101001110010000110010000110100001001100;
#1 $display("%b", po);
# 1  pi=207'b101101100101000011001011100011010000000011000001001100101111111110000000001111011001111110001100011100000101011110101001000001001001000010001001100111101010110011011011111111000011001000000110111000100000001;
#1 $display("%b", po);
# 1  pi=207'b001011100010101111011110000011100111001000011000110101010100111101101110111111111101000101101000111000011001100001000101000001100100100101001111111111101110111111000101011001101110111010011010101001011011100;
#1 $display("%b", po);
# 1  pi=207'b110111101011011111011001100000110010101110100101000000010101110000100000110101000011011001010110100010111000100010110011101111100011010011010011110100110111010101111101000110110000010001110101011010000001011;
#1 $display("%b", po);
# 1  pi=207'b111011101010101110111111011011000001100101111111011111001110111000100001001011101011000010111010000000000100101111001000011010001101100000010001110100001111101100110000111100000111001000001001000100100111001;
#1 $display("%b", po);
# 1  pi=207'b111000000110111111001010000110110110100111111010110011111111101100010101011011010101011011110101101111001111111000011001110100001000011000011001000101111110000111110111001001100000111111111000010101111011111;
#1 $display("%b", po);
# 1  pi=207'b001010100001100001110001111110110110000001111000000111101111100101110011101101110101011010101101011011000110001000111100010000100101100100000101001111100110111101100001011010101100010011000000111100101000101;
#1 $display("%b", po);
# 1  pi=207'b001010000100100101011100011001011000101110010100001110111001010000110111110111111000101001001100000100101100000100101000100111001110011000110100001001001010111110010110000100101100000001001101110010010100111;
#1 $display("%b", po);
# 1  pi=207'b010101011100001100101101100111010001001001101110010011111001110001010010001101101111110101000111100001111010010011001100000011100111110100000000010000010100010100111010110111110010011000101100100000110101000;
#1 $display("%b", po);
# 1  pi=207'b100000111001101100111011000101100000000100111111011110101110100001110010001011010000011010011000101110101101111111101110101101110010111110110000100000110010001111001110111011110100000111110001111000110111101;
#1 $display("%b", po);
# 1  pi=207'b100010110000111010100010011100110000100101001011100100011001101000101011011101011111001110111011000110101001101001111000001010011111111111010000100101111011100101100111010100000111010100101010110111011111000;
#1 $display("%b", po);
# 1  pi=207'b111011001101011100000001010111000011100010001100010100011000101001000101110111111110111000110000111111101101101111011101101110011110100010101000101010111110111011001010110100101010100011101001011011000011101;
#1 $display("%b", po);
# 1  pi=207'b011110010001111110111000101001110101011101001111011010010011110100000000111101101111010011001100101110101000010111110000101011100010100000101100111100000101111100100001110000011110100000011011101110101100111;
#1 $display("%b", po);
# 1  pi=207'b101011001011101110100110010000010111100101100010111001100010111011110110110010001001010111001101011000011000000111011001010111100000100100111110000111111101110001010100111000111001101110100110001010010011101;
#1 $display("%b", po);
# 1  pi=207'b000111111010000010110010011101100100111010110100000010001010110011111100010011000001011010011010010001100010010100101110011000001011111100001011000000011010010011000111111101101110110100010001101001110011011;
#1 $display("%b", po);
# 1  pi=207'b001010001011011101010011011000001001001011111011111010010101011111011011100000101011001000110000001111001100011000110010111100010110001011011111010110101010110001110001100001011111100101110011111111010000110;
#1 $display("%b", po);
# 1  pi=207'b011001100011100110110110101011100110011111001000000010101010010110001110010100100110110100100010101010010100110110111111100011001100111001111100010010001010000001101010100101000000100100111110111010010110000;
#1 $display("%b", po);
# 1  pi=207'b101111101000100111111110100000010111010111001011110111011110001101001111000011100010001011100100011100001011000101111100100000110000000111110010100000010000111110000101001010101100111100101110011110010010101;
#1 $display("%b", po);
# 1  pi=207'b000111010111111000001101111100110000001100101001011001000000101011001011101111011001111111000011001000111000101110010000100110101001011111001111010111100111010000001111000110101011011110111011001000011101110;
#1 $display("%b", po);
# 1  pi=207'b000100001101100001001010001111100001010011001001111111011000111101110110001011100110001010000010110000000001011000100010100101011011110001011000011111101110110010011000101001000011111011000011100111100001010;
#1 $display("%b", po);
# 1  pi=207'b110010011110110111010011001100110100010110010010101011000000011000101100100010101101010111101000110011010010101000101110011000111110101000001110000110010100010101101100001000010001100010101000110001011010000;
#1 $display("%b", po);
# 1  pi=207'b111100000110011110001111000111100000001111010100010110000000000100100111001101111000100000001000011001111001101111001001011110001011000011010101110110101000101100001101100000001011001011110010001111110101110;
#1 $display("%b", po);
# 1  pi=207'b001100111100011101001010011111111110100111010000001100011101110101000000011000001011010011101001110000001010011011100100110111010010100011101111100111010000111010001011011111011110001010001001100011111111110;
#1 $display("%b", po);
# 1  pi=207'b011101000111111000100010000111101111010011010110000111010101110110100110111110001010001011111101011010110100100011010011100011000011111110001011011011001011101011001100000001101100101111001110101100111110011;
#1 $display("%b", po);
# 1  pi=207'b110111011100110011001111101111001011111101100001011100001011010111010100111011000011001111001101000110000010111111100000101111000111110001001111011101001001111011010001001111101110100001001010011111100010001;
#1 $display("%b", po);
# 1  pi=207'b001000100011100011011001101011110110011000011001111001010110100111001000100001101100110101111011000010110010010100001101001110001001100100000001101000010101110001011111000000011000001011000010010101110011010;
#1 $display("%b", po);
# 1  pi=207'b100000101000110000101101101110101010100010111010011011100011111011100111100111100011111101011100111101101100001101011110110001110110001111011001110011101101100011000000001111001001010111001010011001101011101;
#1 $display("%b", po);
# 1  pi=207'b111001011101111010111100111101000111011010010111100001101011000110000011011000011111111101000110100000010001011100100010001010011011011100101101011110111011101101000100010111011111000011101111100110111011110;
#1 $display("%b", po);
# 1  pi=207'b000011101111010100110111001100111111011001110001100101101101111001100110011000000000111100100010110000100001111111111111011100100110111011010001110011010010100011110111110010101001110000000000101100001000110;
#1 $display("%b", po);
# 1  pi=207'b011011101110001001101010111101111010101010000001101010101100001110111001010101100111111001100100100010110101011100101111010011111000110000010101010111011001000010000111000011001000011001011110100011110100101;
#1 $display("%b", po);
# 1  pi=207'b010110010011010101011000000101110001001111000011111110001011011111100110100000000011010101110010110111010000010111000110101001000101111101110001110101101111110111111101100011100011100000101010111100100011110;
#1 $display("%b", po);
# 1  pi=207'b101101001111010110011011111001001110110000100110111100001110000001010100000000110101001111000010101111111100010011001110011000101101110000000101101110111000100101001100001011101100111100000000001011001111001;
#1 $display("%b", po);
# 1  pi=207'b100011101001110111011011110001010000010010001011101001111001011101100010001011000110010010000001111101110000100000000100000101010001100110000011111101110011001100001010101110001011011110000010111000000111101;
#1 $display("%b", po);
# 1  pi=207'b010011011001011011100010000111010111001001000100001001001101010101110111100100101000101011100100110111111110000101101101010010010001111000110010010010101110001111110001000110101101001101110111101111111000000;
#1 $display("%b", po);
# 1  pi=207'b111110011110100110111101111000110010111010010110001110000100001000100011110000000110010100110101110011001011001011000100001101000011001101011111000000100011111011010000100100001000110000111011001011011101110;
#1 $display("%b", po);
# 1  pi=207'b000000000001110000101100100110101010101000110000111101001001110011110000001101101000000110000110001000001001011111010110100100011000011110110010001101010101110101110011000000110011110000101000010101100101111;
#1 $display("%b", po);
# 1  pi=207'b001011111001011001100111001000001000010101101001100000100011011010101001010100100110000010010000101000101001111101000110000000110111010000100001001101110001110111110010011110011110111011101011001001010101100;
#1 $display("%b", po);
# 1  pi=207'b111100011001011101011010010011001110100110111001110100010001111100011101101100111011100101101011100010010110001001001101010001010101101001010110101101101100010010000000001011011001111000100010000100111011111;
#1 $display("%b", po);
# 1  pi=207'b010001000101001011001110111110010011100011110011110000111111111000101110001110110101111110000111111001010100011100110111100011111010010111110000110001111101110101001011100100000011101010101010101110001110111;
#1 $display("%b", po);
# 1  pi=207'b111011011111110011011100110001010011010111100011000111100101100111100001101000100110011111001010100000000110100111101001111010100011011111100010100110000110001010101110111011010010110000111111101111010000100;
#1 $display("%b", po);
# 1  pi=207'b101110110110100001010011011000101100001010101100101110110111111000110010000100000101111001110111000111010101011001000101100111010001011011001110010101110111111110110100011100101110000000000011001100111101110;
#1 $display("%b", po);
# 1  pi=207'b110010001100001100100111000000100011011011100110100001001010000100111010010001010000001111000110110000010010110001101010111000010110011000101111001011010110110011110101000110110100001010101010111000100100011;
#1 $display("%b", po);
# 1  pi=207'b001010001101100010011111010101110100111101001011111100010110001100000111101010110101110000000001111000001101001000111001100110101010000001011000100011001111110000100101010111010011011110101011010101100001110;
#1 $display("%b", po);
# 1  pi=207'b101100110111111100100100000001110001110110001111101100011001100001110000100111101110101011100111010110010010011101111011100011101100110001101000011110101010001110011101000100000001101110001110010110110101101;
#1 $display("%b", po);
# 1  pi=207'b111001111110001101111100100000011101111011111110001110111001111101011000101111110001101111011111101101001101000011000011001001100001011110100110111010011101001101010100110110100000111111001110111110010110011;
#1 $display("%b", po);
# 1  pi=207'b111000111001101001111110011010000001101110010001011011110011011011000111001000111101010111001000001110010111101010000101111110110101011101111111001010100101011111110001011100001101001100010100010011100110010;
#1 $display("%b", po);
# 1  pi=207'b001101111010000000010100010011011001001100000101000011101010001010110000110110111010110101011000010001001011010011001100111100100111100111011100100101010001001101001111011011010000000011101011100011011110011;
#1 $display("%b", po);
# 1  pi=207'b100101110100001000110000101001000100011000010001010111100011011111011110111000000011110010011100011101100100111001011100110001001111100110010110101000000101100100110000110011011001100001110101100010101011100;
#1 $display("%b", po);
# 1  pi=207'b111010111111100000111011110101100011011010111001101100100100101110110010011000010011100100100000101101001011110010010100000110110000111011101001000111100001101010001101001000111001011001111011000101101100100;
#1 $display("%b", po);
# 1  pi=207'b111110001100100111011100101111100101000011000110100101110001010111110010100011011011101011001100111111010001001101111000101101011111100111010001000010100101100001100000011001101110101001100000010100010010011;
#1 $display("%b", po);
# 1  pi=207'b001010011010111010001000000110010110111111000010100100011110111010011100111001100001100011010011010001000110100011001010011011111111110001001001011010101111100000010101011000100010010010100000101010011111011;
#1 $display("%b", po);
# 1  pi=207'b000101101100010011100010001011001100001000001011111100110100111101110011001111110011110101100111001011000110001010100001110110000001001000011000001011001101010001011101101101010100111101111100111010101010101;
#1 $display("%b", po);
# 1  pi=207'b001000110100101111110100000111010110000110000001101101010111001101110111001110001100111000110100101000000010000110000111010101110010110110111000111110000111000110100111010010111111100100010111001010011111110;
#1 $display("%b", po);
# 1  pi=207'b100110011000101010101100000010000010001101101100111101100010011100111001101011101101100111100011110000001000011101001100111111111010100000111110001000111100101101100011111000000101000010001101101001001101010;
#1 $display("%b", po);
# 1  pi=207'b011010100001111110110110000010111000110100111000010111110000001001011001001101111110001100101010011010000111001101101110101101111101001000110111100110111001101100011101000010001010011101100100100100110111100;
#1 $display("%b", po);
# 1  pi=207'b001101001101101101101110110110010001010100000001011001011011100000001011010101110101011010101000000111000001111010111011001100101011111100001010011100010001001101110100011000110101010011110100001001001101100;
#1 $display("%b", po);
# 1  pi=207'b111010100100100001010110010001100110011000000011010110011001000010000001110011101001010000101000000110100000100101001100010000001110001101010101100000001101101000110111100011100011110011000100011101011010010;
#1 $display("%b", po);
# 1  pi=207'b111010101000110101100111110100101111001000100000011000110001101010001110011100110110000000001111101001111110100111110111101110010111101001101110100110000001000111000011000010100010001100101100000110111101000;
#1 $display("%b", po);
# 1  pi=207'b110011011111100011000011001010100100010101100101011000111000110111011011000101100110011111001101110110000100100000001000011111110010011001011010011101000111010100110011011110010000101101001111001011010000110;
#1 $display("%b", po);
# 1  pi=207'b111000011001011101000111100101110011000011110111011000100101010000010001011111110101111110010011110101000110101111000001001100110100110010000101000000100001001110010101100011010001011101000101110100010001100;
#1 $display("%b", po);
# 1  pi=207'b110001001101111110111010011011110000011111010010001011111011110101100101010100100111011011110011110001010111111001001110000110011100000101101010010110110000100110011011111010110101011011111100001101001111100;
#1 $display("%b", po);
# 1  pi=207'b111110011011010100100101110100011101011010101110001011110111100011001100111111110010101100100010000000100001100100111111011110100110001110110101100010110011110100100010111101100011110111100101001101011111010;
#1 $display("%b", po);
# 1  pi=207'b011010101000100001111110000101000001011100110010001110100000011000100101001010101111110001110000100010000100101011011000010101110111001011010111100110110100001001101010011000101101100000001000001001101000111;
#1 $display("%b", po);
# 1  pi=207'b100110100100100010101110001110000110110001100000011011101001001000111011001110101111011111010010010000010101110000111001000011001011001110100001101010000101100101110101110011101101011111100111111010011011010;
#1 $display("%b", po);
# 1  pi=207'b101111011100100101000010101000111111111110100001111000101010101111010010011011100010111011000110011111010000100001101010000110010000001000000000100101011101101001000110010011100110011101100110100001100010110;
#1 $display("%b", po);
# 1  pi=207'b011101100100101001000111001011011101101110110000101011100011000010101111000011010100010011011111111000010110000111001011000011100100000000001010010010011011110010000000010001111100100101110111001101001000000;
#1 $display("%b", po);
# 1  pi=207'b100110000100110110001001010011010111110000100011010000011011100010101001011100001011110100111101011010000000011001100000111101110011001110001001010101010110100010110100001110001110000010111000000000101010110;
#1 $display("%b", po);
# 1  pi=207'b110010001100001011011110101101000100100010010001110011011010011000110010010110101101100010000000100011000101011100101000111011011011001100111111101000101011100010100100111101001111101000001101011100000010111;
#1 $display("%b", po);
# 1  pi=207'b001010100010101001000000011111111011011110001101000011101001111010011111010100011101010001001111001110101100000011101101000111101101000110110100101000110110101111001111011001000000001111100111101100001110110;
#1 $display("%b", po);
# 1  pi=207'b110100101110110010010001000000010010010100011101000111001111011100100000000010000000100111111111000100111001000110111011110010011010001001001100000001100110001000001111011000110111110110111011110000100001101;
#1 $display("%b", po);
# 1  pi=207'b101001010111101001110110101010100000001110101011101010011110100011010011111000010001010001100100111111010110100000010001011100101100110100100001011000111100101001111111100010111001100111010100111101101110001;
#1 $display("%b", po);
# 1  pi=207'b110001011101000101001110010011110110100110011110100000001100000111101001111111110110001010000000110110100011111111010100110010100101101101000110001111101010110000000111011101111011010001010010100010001111110;
#1 $display("%b", po);
# 1  pi=207'b010100111011111110111100111000010101111111110111001001111111011000101001011010010010000100100101111011100011011111110000010010110101111001010010110000000111011000100101001111001100011100110111110100101010100;
#1 $display("%b", po);
# 1  pi=207'b111011110100011011110100111000101100100110011001000010111100010000011010001101101001001001001000100010111101101101000010100111111010011110001000000100101011110111101110011011110000110101111100010000000111100;
#1 $display("%b", po);
# 1  pi=207'b011000001000001101100101001011111000111010100001010100101011010100111100101110111110100001100111001101010100111000011110010010000110010011011101000010101011000101101001111101000101101010000101101110111110110;
#1 $display("%b", po);
# 1  pi=207'b111111010001111010001101100110101100011010010100010011111001010110000100011001010010001010010000010111101010111111101111011000011001001110111011100111111001100000001010011100100100001111000001010010110100001;
#1 $display("%b", po);
# 1  pi=207'b001010000111001101010110011000101010010000100001001101011100101100111001001010001111010110100100011111111100000111111111111011000110110000100111001000011111101001000000010000011001101111111001110100001100010;
#1 $display("%b", po);
# 1  pi=207'b000111110111111000101001110110101110101100110010000010001010101000001001011010101110111011110001001100110100000000100001100101011010101111001000010101100001010100010110111011100101101101001010011010110011010;
#1 $display("%b", po);
# 1  pi=207'b100100110010001111000110000001001000100011010000011100101100000111011001110001111000101000001010001000011101001101110010010111100010000101001011001000110011111000100010100010101011101101000100011010111010010;
#1 $display("%b", po);
# 1  pi=207'b111110011011000010010010110100101010000010100000001101000111010001100001101001111100110011011101010101110010101011110001011010011011000010101010001001011100011011000010011101111111100100011100001111100001011;
#1 $display("%b", po);
# 1  pi=207'b010101101111001000001111110101101110000001100111101001001010110011001000110100000101010001101101110100101101011001100001001011100010001001110001100111110111111101101100001100110010111011110101101010001111101;
#1 $display("%b", po);
# 1  pi=207'b101011101010010101111000001010110111100111011010110001011100011111111011001000011111110101010011001010001101111011000011100001111001100100001101110001000001111111011011001010111100011001010010110110010111100;
#1 $display("%b", po);
# 1  pi=207'b100011010000110010011110011010011111101011100100010111000011000010011101001001000000001000101010010110111000001111011110110111010001100001011000001110011110100011111011111111110111010110100010011111011010011;
#1 $display("%b", po);
# 1  pi=207'b001100100000101100000001001100111000111011010000001000100001010010001011011111111101001110001100101010011000000111001011111100001011110011011100110001000000101000101001111100001010111100110000110011010011000;
#1 $display("%b", po);
# 1  pi=207'b001001001101111110011010011010101100010010010000001001110000001110000111101011110101101100010101100001101111101001010010101000111000100000001110010100110011111001010011000010110111111011010100000000100101110;
#1 $display("%b", po);
# 1  pi=207'b011000000110101101111101110001000001110011101000011000110011010011101111101110001111001110001101000100000010111000001000000100000110111001100110000101110010000000010001000110000101011010010001101101100000110;
#1 $display("%b", po);
# 1  pi=207'b111011101111000111011001011101010000110100010110011100110001001011000010000111000110010011100001111101110000011001001110000011101111001101101100111001010000111000011111111110110001100100100100011101100100100;
#1 $display("%b", po);
# 1  pi=207'b011001111011100111100101111010000110100100001011100100110100111111011110001010010110101001011110010110001011011000000100000010000101111100111011001100000011101011010001001001011100010001100010000001010000100;
#1 $display("%b", po);
# 1  pi=207'b110000011011001101110001101010011010010100011100110100001100011011000101001001000111101011000100101110101001011110100101001011010100001010001110110100110001010001001000110010101001100001010111011010101111010;
#1 $display("%b", po);
# 1  pi=207'b101111010010010100001011010101011001111110110001111100001101010110110111101000000011101101011110010010100100001011010010010010111101110101001011000010111100010100111000100001000111010011111000000000101000001;
#1 $display("%b", po);
# 1  pi=207'b111000011110101011101110011010010000101111011010100001101101101011010000001001110100100011001000111000001011110101101011001101111100110001101001010100011111100101010010111101100011001001000011000011110101000;
#1 $display("%b", po);
# 1  pi=207'b011011011011000100101111010101101110111010100010110110011101110111101100001000011101011010100101110100010010001010011011010101111010011011011100110011111101111001000100111111011011101000101111000100101001000;
#1 $display("%b", po);
# 1  pi=207'b001111111111000010001100111110001110101000101011110110001000010001100110111111100011010011001101100010001110000011110100111110011100011010000010111001001000100101100111100100011111100000110101101111100110111;
#1 $display("%b", po);
# 1  pi=207'b000010011000000111001001101111100001101011011101100010100110111110000011000001110110111001110110100101100001100101000000101000010000111111111010101010101010000010111010101101001100110010010111011111100111110;
#1 $display("%b", po);
# 1  pi=207'b100011111100111101110011010000001010011101110010110011111011001000101100110110111010000110111111000010110011000000011111001111101100000110100001001011001001010011100010110000111101010101000100010111100001010;
#1 $display("%b", po);
# 1  pi=207'b010011001010110001000110010101100010110011101101100110100001101001100000010111010001001011100100001111101011010010011010111100111111101101000001011101100010100100111110000001111111011100101101110101100001001;
#1 $display("%b", po);
# 1  pi=207'b100000000101100101110110001100111101010101010000111101001111010010101001011011101010101010101011001100111001101011001100010011001001001010011001100100011010000100000010000101111000001100100001000101000101101;
#1 $display("%b", po);
# 1  pi=207'b010001111111100011100110111100010110010001110000000100101101111010100110001111111100101111110011101110101000110111000011111010100100111001000011011001100111110001111000010101010110010011111011010101110110011;
#1 $display("%b", po);
# 1  pi=207'b111001000011111101111000011011110110111010110100000101100111001010011000111010100111111011010000101101100100100011011111110001001111000100111111010010111100101101110011110111010100111110010000011101011000110;
#1 $display("%b", po);
# 1  pi=207'b001010111011000010101101100110011001001100001100010101000010101100100110001110000001001110001101100000010010010111111110000001110110101001101001101010100100101100100011001110101011111011111110000011011000011;
#1 $display("%b", po);
# 1  pi=207'b001101000100010001010100011001011010111011100110000111110000001000110111011000111001111000110100010111100001111001111011011101001001111110011000111000100111000011010011010100111110111010100101011110100010010;
#1 $display("%b", po);
# 1  pi=207'b101101100111010110111011000110011100101100111010111001001110101110010000100001110111111000101001001011110000101100100100110100100000101001101101001011111110101100101101010011101111011110010110100111111001101;
#1 $display("%b", po);
# 1  pi=207'b110000110110010100101011110001111000110011110100101011011100111001001000110011010110100111001111110111101000111110001001000111101100100110111010111011001010111011000100001110110011110111010100010100111100111;
#1 $display("%b", po);
# 1  pi=207'b100110010111101011111110010100101101110001100110110011011011010100001110101100101000010110011101000100011101100111011101100111101111001010110000111111010110111011000101100000110001110110010010001010101101000;
#1 $display("%b", po);
# 1  pi=207'b111111010001110111111011000101000001000011111010110001000110000001011100001010101111111100111110010011111101111100000010100011111011010001010001000011110100000101010100011001001100101111000101110110100100010;
#1 $display("%b", po);
# 1  pi=207'b000010000011011110110010111011110101110111010100001101000100010011110101110001011000011101110011100001110111001100111111011110111010100010011000000000010100000000001001111111001100010001110100011101100100110;
#1 $display("%b", po);
# 1  pi=207'b100100001000101110101111100110001010010000001101100101010001100100110101001111100010000110101001111011100100110001000011110011110111111001101010011000011001000111111011100101011101010110000101010000111111010;
#1 $display("%b", po);
# 1  pi=207'b011111100101111011100100111101010000000101000000000101011000111001000010001011011100100100110001100000110100010011110111110111000100101001011010100001010000001101100001101001011101111101001010010000110000101;
#1 $display("%b", po);
# 1  pi=207'b001110100001001001101101011011100111011010010110110110001011101111101001101001011000000101001100001001001000110011010001011100111111010000110010110101001100010011100000011010100010010011000010000100001001100;
#1 $display("%b", po);
# 1  pi=207'b000000011001101000101000111010111101111010110110001010001111010100110000100101001110101000010000110011101101111110011011001001011010100110001011101101101011010111000110111101100010011111000011100010010100100;
#1 $display("%b", po);
# 1  pi=207'b000001010110111011111000001110101110110010001001001010000100011010010011011011100100101000000010110000101001101011100111011010101000010011000010001100101100011000111101100000101100000100110010101101001010001;
#1 $display("%b", po);
# 1  pi=207'b000011101100000110100000110100110111011001011101000110000111010100011111000101001110001100000000101111110100111001111111000000110010111101110011000100110110011000001111101000110001001010110100101011010000100;
#1 $display("%b", po);
# 1  pi=207'b010011000000011110001100001101101111000101010111010111101100101110111100110101110110110001101101001000011011001001110001001111111001000011101100101010010011010011000111101101110001001001111111011111101101011;
#1 $display("%b", po);
# 1  pi=207'b010010011100010110101111001010100011110001011001000101110000111110000011101000001010000000010111000011101100010100110011101010111001101100000101010111001011101110011111100101100111011000001100011001111001110;
#1 $display("%b", po);
# 1  pi=207'b100000100101011100111100001000011011001001011000110101110110000110010000111011110000010111010100111001010000011010000100000000100111001110011011110011010001010001111000100111000010000101000100000101101110001;
#1 $display("%b", po);
# 1  pi=207'b101011110111010011011100110110001001101011011001010100110111111001110011000011010111111111010110000110000110101000000001010000100000000111110000001000000000011101101111100110000111100001100010100110101101010;
#1 $display("%b", po);
# 1  pi=207'b101000011011010100101011000100001000110100111000101010111000011011100011110011101111100101110101110011010001001100111111101110100010100010000001000110100001110110111100111100101010110000100111111111000101110;
#1 $display("%b", po);
# 1  pi=207'b000010000001001100001001000011101010001000111011101110010100001000000011010100001110000101111000100011110111111100101011010100000100000110110001000101101111001100110011010010011100011110000110110000101000000;
#1 $display("%b", po);
# 1  pi=207'b000000001110011100001110101010111111000100000010000001000100010100001010010101011100010110100100011101111101001010111110001010111111011000010101100011010110111000000101001011111101110100110101011110011010101;
#1 $display("%b", po);
# 1  pi=207'b010111111001110001011000000010110010111000000100110111100010111000000100011001110010111001011100001101000000011101010101010101001010001000101010001101000111111001110100011110100011110000101111101000010101101;
#1 $display("%b", po);
# 1  pi=207'b101101110000010011101101001101011010011011000000100100011000100100100101110001110100111110101001011100000010010001001001101000000110000011101101000010001010101100110110110000110011000010101001001100110100101;
#1 $display("%b", po);
# 1  pi=207'b100000011110101101010110001100111000000001100000001101100101100101111000000001010010000100110000100001111100101001100110111011000100010001100100100011111011110001011101000110110000000000101110110100011110100;
#1 $display("%b", po);
# 1  pi=207'b011010100001110110011111011111010100110100011000110011000000110011110110001000011100010001011010001010111001010011011111111001111001001110100000001101110101000101110101110000111011000001001111101110001010111;
#1 $display("%b", po);
# 1  pi=207'b010110110011110101111000101001111100100001100111111010010111101110001110100010011100000101110011010001110001100000001010001101010100000101110011011100011011110101001110000111110110011011001011110100111011000;
#1 $display("%b", po);
# 1  pi=207'b001110010110011111100000111110011101111101101011001011110101011000110000111001011100110011011110111111110001101100001110010110100101111011110001111100110110000011001100011000011101011010101111001001000010100;
#1 $display("%b", po);
# 1  pi=207'b001011000010100011010100000011011011100010110011100010110111100000110110110111100000010110100000100001010111010101110110100000000011101111111011001000000001101000101111010110110001101111111010011011111100011;
#1 $display("%b", po);
# 1  pi=207'b100110010000000010100110011100011111110111110111111111100000011011000100101001001100001001110110101100001000001101100011011010110100101111001000010011010011000110101100010011100011011100100001100110010111100;
#1 $display("%b", po);
# 1  pi=207'b011101000000100100001000111101000001011111000000010010011001101001011110001010110110000101010010001100011010111101110110011110110111101100000100110001110001101111111101000011001111101000100011011000110000100;
#1 $display("%b", po);
# 1  pi=207'b100101100100100101011111000110101110101010010111011001100111011011001101100101111100001010111011010011010000001110110001001000111001001110111110011101111100001000001001010010000001011010001010101101100001110;
#1 $display("%b", po);
# 1  pi=207'b010110010001011111101110010101010000111110000100111100000011111000011011001010101000101010110101001000111110101000001111010011011100001100011110100111100100100100000000111111011101101010100000011111011110101;
#1 $display("%b", po);
# 1  pi=207'b010000101000101100111110000001110000011111111000111011000001011010001111101110100100101101110000000001110011011000011110110101001010001111100100011011000101000010100101001110011111110000111101010101100110101;
#1 $display("%b", po);
# 1  pi=207'b010011110001100001111010101000101101011101011011111010001011100000111000001110110000001110101011101011111110101101001101011100111100001101101101011001111111010100001111101111101000101100010101010010000000010;
#1 $display("%b", po);
# 1  pi=207'b101110000011110010001000110101011010001111001110001001011000111001001111111011001011100001000100100001100011000000111001100111101001101101001111110100010111101010010111101011100010110010001111011101111011100;
#1 $display("%b", po);
# 1  pi=207'b110011100110111001111000000111101001000111011110010100111010100000001101001001001110000010011111000010100101101101011011001011010110000110100100111101100001011110100101001000101011110111100100011000001111110;
#1 $display("%b", po);
# 1  pi=207'b000100101000010100101000001010010010001011101010000010011010001011110110110110000001111011011001110100001101000000100111111111110101011001110110111011111110010101110011000000110010010001111111111101000110101;
#1 $display("%b", po);
# 1  pi=207'b010100100010011110110111100010010000001001101000101111000010101101111110001101101010010110100100000001110001101110100000100000111001011000001100001111110101100011101110111111110100010011001101100011101011110;
#1 $display("%b", po);
# 1  pi=207'b000100111010101101100010100000110001110111100011111000000001111000011010011011111111010001101100100010100100010101110101011000110011010110100001010010000010100000011010001001110010001011010000011101001110110;
#1 $display("%b", po);
# 1  pi=207'b110110000111111001111000111101101000100000000111001011011000001011110000111001111110110111110011001000100110011010101010100010101000101110100101100011001110000110000001011010010011010001101101111111100110100;
#1 $display("%b", po);
# 1  pi=207'b001001011001010101111111100101101101001111010111111001010011100000001111100001100001111010010110001100110101101101110010011001100100111110101111111001000101100011111000111100000110100101100110011100101010101;
#1 $display("%b", po);
# 1  pi=207'b001011100010101010100000011101100011110111001000010000110111100000101001101110110110110001100000001011111010110111111100010111011100000100011101000101011111011011101101111111111110001111101010001101010100000;
#1 $display("%b", po);
# 1  pi=207'b111000111101110111010100110101100111101110100100100100111100110000011011001000000010100001011101110110010010001111010100110110000110010010101001000111100000110010101011011011010010111100110100010101001101001;
#1 $display("%b", po);
# 1  pi=207'b000111110000000100010011100100001100001000001001101110111111010100010100000111111100001111001110011000101000111101010101011101100111110001011100111100111011000100011101001001001011101111000010111001110111010;
#1 $display("%b", po);
# 1  pi=207'b000001101101100001011011110101101001100001110000000110101100111101011101010111101001000001010111001111100111111100011001000110000000000001101111110001000010110111110100000110001100001111101001110100010100011;
#1 $display("%b", po);
# 1  pi=207'b000010111001011010011110111110010011000111010010100011110110100100010000010010010110000001100001010101100101100001011100010011001001110101110010110000000001111001100010101000001110100001101101011001010101111;
#1 $display("%b", po);
# 1  pi=207'b111001001101100000010101101110011010100100110110000011001001100110011101111000011000111000010011001100010111110101000111000100001111111111111110011000000010010101010010100001001100110111001000010110110111011;
#1 $display("%b", po);
# 1  pi=207'b100111111101101110010111101100111111001110010010010101111000011001011110111010010111110010001110101010011100001000001101111101110011111010000110000110001010100100000110101100100110110000101111010001010011010;
#1 $display("%b", po);
# 1  pi=207'b111001111101001111100011110110001011101111101111010001011000000010110000000100011101001011111111110110110011010110101010100111000000011110010001100110111100101101010011000111100011000101001001100100110001011;
#1 $display("%b", po);
# 1  pi=207'b011100110000011011010000101001101110110000010011100111000010111100110000010000010001110101111011011000000111001011010100110010111111111011111101101010110010011100111100011001100001101110011001110000000111001;
#1 $display("%b", po);
# 1  pi=207'b011111011000011110000110111011100001011001001011011111000101100001110100100010111111011010010110011010110010000011001100101111100101101111100111000111111100100111110000110110101101001111000100000100000000101;
#1 $display("%b", po);
# 1  pi=207'b110100000110010101111101111011101000110110001011011100100110001110111111101001000100100111011001010011111010011010010001000011001110111111011111100100100010010111011001100001001111010001101110100110000011110;
#1 $display("%b", po);
# 1  pi=207'b101010011001100101010100000011011001001110110101110001000001001111100010100001100111000101000011011001100110001000110110100010101000110011000010000010101011011111010011001111111010000000010110000001110001111;
#1 $display("%b", po);
# 1  pi=207'b101111011110010001000001111011111110001011000011101110110100100001000101011001000110111000111010001101111001000110110000110010001100001101111000110011110110110010100101110111011000110011000000101011111000010;
#1 $display("%b", po);
# 1  pi=207'b010010110011011010110010100111101110111010010101001010100101010101111000100000111000101110001100010010100000100010100011101100010001110011011000101100001101100011111111011100001100010110011110110111100000100;
#1 $display("%b", po);
# 1  pi=207'b011111011111101001010011001001011100100100100010001001000010010011101110101010111010011011110011110011100001100101110000101011010100000000111000010100101111111011011100111010100000010001101110110110111001110;
#1 $display("%b", po);
# 1  pi=207'b101011001111010010110000011110001100011010100011101100100000111001101101101000010011101011110010100101100101111111110101101010111111100101011010111110001001100100011101010101100101110101101011111111011000101;
#1 $display("%b", po);
# 1  pi=207'b100001111110001011010101001001001001111100100100010011100011101000110101000110010010000011110011110011011000110010111001000000100111101010101001011011000110111100011111000001011110001100111110111100110110000;
#1 $display("%b", po);
# 1  pi=207'b110111110101101000100110001101010011101101101010110010101000111101101100000100100001100001101100000000111001100010100100100110100001110000111110111010110010010000000100001001110001011000110110111000001010010;
#1 $display("%b", po);
# 1  pi=207'b101101100010001100110101100100010100100000111111100110001110011011110000011101111000110110011001001100100010110000010110001001100101001110111100111010110011100111101101011111111001111110011010010110011101111;
#1 $display("%b", po);
# 1  pi=207'b101001101011000101011011101101101100000000001011001010010011000001011101101001111000111001001000101011110011010011001101010110110111101101110011101010111000110111000011001101010111011101110100101100010111101;
#1 $display("%b", po);
# 1  pi=207'b101111001000001110101100001110110011100000110100010010011010100011000100011111110101100101011111011111010010111101001000001011011100111110100001001011110111110011001110110011001001000000011111000011001111011;
#1 $display("%b", po);
# 1  pi=207'b111101111010000000110011111011110010000011110111010000001000110110000101011010011111101101011010011010000000000100111010000100001101100011001101011010101110000010000001000100000000000110001110101111011111001;
#1 $display("%b", po);
# 1  pi=207'b111111111011011101111110011000000100111000111100111110000000100001001111101010111000110101000011100001010000100111110010001111000001111101011110001101000000100101010010100010001011110000011111001110110101001;
#1 $display("%b", po);
# 1  pi=207'b011111111111000100001110001100110000001110001110110000000010000010010101001110100011000101010000011100001100111001101101000011000001111011101011111100110111011010101011001001000111101101001101111000110001100;
#1 $display("%b", po);
# 1  pi=207'b101011000111000110110001110011100001110100100010100100001100110011001100011111111001111000101010110101001100110000101101010000110111001100011110001010110110001110110000100110011111010101100001011010001001001;
#1 $display("%b", po);
# 1  pi=207'b000101010000111110010010000001110000011011001001101011011000010101111011010001110010011111000100101010111111101010000000101000001111100011001010010110010111010011011010011111010101001000110000010011010010010;
#1 $display("%b", po);
# 1  pi=207'b010111000011110111111001111110111011110000100011110100011001001111001011000000010100101011100110100110010110000110101000110110000000111110000111000111101110111101110100111110001111000111000000101001001110010;
#1 $display("%b", po);
# 1  pi=207'b110110001101110010110000101011001111111000101001111000110000111001100011011110000010000000110111111110101101000100000010011000110000011100000100100000101000011111010111010010101001111010101110011000100001100;
#1 $display("%b", po);
# 1  pi=207'b101110110011110001001111010110100010101010110100101111001011111011100000100011001010101011000111101010000101101000100010001111010001100101101010011110111110100101001010011000111100110010010001110010100100011;
#1 $display("%b", po);
# 1  pi=207'b100111011001011001011011101010101100011101010010000110000111000000100110110001111001100110001111001111111111001101111011010100111100110001101100110100011001000101000101001101100001010010000011010101000011001;
#1 $display("%b", po);
# 1  pi=207'b000000010100100011100101001101111111000010110010101001011011100001011010011000000111111111111010001000000111011011111011011101110011000001000001001110010110100101010010010100001000110000001100111111111100010;
#1 $display("%b", po);
# 1  pi=207'b000111110010100110111111000110101010101011100110010101100100000100111011001000110010110100111100111111100111100010110111000111000111000110100100000111000111000000000101011000100011110011010100110100100000100;
#1 $display("%b", po);
# 1  pi=207'b110010000010101011011001110110010111110101110000100011000101010000010101000101101110100001010011011010101011101100010101001000010001101100010010100000001001011010111000101101101000011111100010000010010001001;
#1 $display("%b", po);
# 1  pi=207'b001010100110110011010000110110010001100101001101100110000011011011110111110001110000011011111010010111110000001011110001101100010011011110111110000011111010100010001011010010011110110001001000100101001110000;
#1 $display("%b", po);
# 1  pi=207'b110111101000101110000110001000011101000011110111011010100011001100000110101010001011010100001011010001100010001111110101101000011101100111001101000100111101111010011110111010001010100100010011101010101101101;
#1 $display("%b", po);
# 1  pi=207'b110111111111100111000011010010110001010010010100100001101011101011011000010100101000011000010111101001100000010101110100100110100001010000010101011000100000110001001100100101100100001011011000011100111101111;
#1 $display("%b", po);
# 1  pi=207'b011101010111111011100111100011111110111100000011010101001000010010011010010001000000010110101000100101001010000010110111110111111010100110001000001001110000011111001001100011010110010010010010010111100010101;
#1 $display("%b", po);
# 1  pi=207'b110000001111001000000100101100000001100111100111101000110000100011010011110110011011100001110000011110000110001101110001100011001100100010001111000111010010010011010010111111101101100110111100110100011101001;
#1 $display("%b", po);
# 1  pi=207'b001101011010110001000101111010111001101001000110010101101111000001010000110001010100111001101101001100010000011100010000011110011100001010010010010000110100000100111110101001101000011011011101100110110110101;
#1 $display("%b", po);
# 1  pi=207'b011100000100011111011111001011011011110010001000001111010101011100111100010010100101011110011001111110110100100010111101101100101100101011111001001001110110111101011010101010000011100100111000101011101000000;
#1 $display("%b", po);
# 1  pi=207'b101110010101000101011011000100001001101010111100001001010111111000011000101110000010000100100001110001010001111111001111011111010000111010000001101110000000000011110111101000101100110001100011000100101001110;
#1 $display("%b", po);
# 1  pi=207'b111111011011110010001011000100110100100000100100100011001111001011010101110111011101100011001100100010010110101110100100111000111011000011101000011011100011110101101001111100000101010000000010011000001100110;
#1 $display("%b", po);
# 1  pi=207'b110101011101110001100001110110101111100111111101111110000001011011011110101000000001101100101110010100011110111011001101110100010101000100110010111000101110001100101000011000001000000100000101011010100000111;
#1 $display("%b", po);
# 1  pi=207'b011011110001001110101010001000001111001011110101101100010001010010100110001111001001000110110100111000110101001100100110001010101010110010001000111000011000100000010110011011001111111000011010100100011100010;
#1 $display("%b", po);
# 1  pi=207'b010110100101100111001110110111111101011000011001010100101110000100000100110010010011000101010101000010101101101011010110100111000111000011001101101110100101101000111011110000001111111011011000000110101011101;
#1 $display("%b", po);
# 1  pi=207'b101101000100001010011111011111101110001110010010101110101101011111110010101111101100000010110011001000110100111101111111110000110100110100010110111001001010101101000000011100100010011101100111000000000000110;
#1 $display("%b", po);
# 1  pi=207'b111011011011001110010010111110110011110011110111001111111111000110011111100100001101101110111010011111001011000101011000101001100001011111100011011110101100001110101100100011111001000001110100001010101000111;
#1 $display("%b", po);
# 1  pi=207'b010000010011110010010111101100110110101101001100001001110111011100111010101010011010000110001111001000110010111101010001100110011010000000101001011111110110111100010101111100000010011011110111001100000111100;
#1 $display("%b", po);
# 1  pi=207'b000100101000111110000001010110001100101110010100110110110100101000101011110011100101111011100011111100110111100001001101100010110010110010110010000110001010110110001100001111000001010010001000100100111101011;
#1 $display("%b", po);
# 1  pi=207'b111110000101011100010000111010011010100101110100110110001001100010001110111100100101110111000110001110010101001000111101100101111110101000011100110101100010101100001001001010000100100101000111110011100011111;
#1 $display("%b", po);
# 1  pi=207'b110100111110110111011110011010100011010100100011111100111010010100111011100111000001010111111001010101001100010001001010000000100110001011011000000111100001110001110001010111101010001111111101100001101011101;
#1 $display("%b", po);
# 1  pi=207'b100001011100010111000011011011000110011000100001111101100010101011100011010001100111111110010101110101110011110000000000001101011110100100101101110001010000111110001110011011100000011001010110011111101000010;
#1 $display("%b", po);
# 1  pi=207'b001100110111111001001100000100101000110010011000010010001011110010011110111011100110110111110010011110101011000010000110100000010110011100101101000100000001010110100101000000101111110010000100011101101110100;
#1 $display("%b", po);
# 1  pi=207'b001011100100011100110011001100101010011111101110100010011011100001011010011011000100110111110101011000000111010100001000000011010110001010010100011101000100100101001101000010010010011101111110111010001011110;
#1 $display("%b", po);
# 1  pi=207'b101000011010000001000100001011100010101110100100011100000101111010100000111010010010101000010001001001110011010100101010010010101011111011100000000101111101100111010001101000101001001001110101000000001110010;
#1 $display("%b", po);
# 1  pi=207'b010100101001001001110111000111111011111000101011101100100011111101100111011000010110100101000101100111010101000101001000100010101100000001010000000011100100011110111011111001111000000101111011010111000100000;
#1 $display("%b", po);
# 1  pi=207'b000111111111100000011001100001100000010010011011000100100101001101000110000010100101100000010011110111100111110010010010000001110010001111110001100110110110111110110101010001011111111010000101110101000111001;
#1 $display("%b", po);
# 1  pi=207'b101110111010100110001011111001101001101010000101011010010101110111101110101101001010001001111001010001000010001101111000000100010001110110000011001101010010101011001111101111111100000111110011000110001101000;
#1 $display("%b", po);
# 1  pi=207'b100010101000001110011010011011111110010010010110001110010010011110000010111110111010101101110011001001011111100111010000110100000111101010100000111110000011111000110001111010010111110001010011110011100110110;
#1 $display("%b", po);
# 1  pi=207'b011010111100110100111011010001011011111010100010011111000011101110100110110011100000010000001111001001110010100001000111110001001011100001111010100100101011101010010111110000010100111000111010010110101100000;
#1 $display("%b", po);
# 1  pi=207'b110111110100111101110001100000001010100010100100011101011100100000101111001110000101111110101111111100110101111100000111110000010100000100111000000000001000111100110100111101011010001101010001101000110011101;
#1 $display("%b", po);
# 1  pi=207'b001101011010001101001100110000001000011001001101111001011011010110110110100010101011111010010000010111110011110110100011000011111010111100000000010000000010000110001001110010000000110101001100111011011101111;
#1 $display("%b", po);
# 1  pi=207'b100110010111110100011101100101010101001111011010001110111010110010110101011111001111101011010110101001111001011001101000011000111110100111111011101000110111010101101010101111010000001100010010010100010111111;
#1 $display("%b", po);
# 1  pi=207'b011110001001001100000110101100011110011110010111110111110100000011101000000110111111110111001110011000111000011010110111010111011000100011000101111011011111100110001000101010100001100100101001111000011000010;
#1 $display("%b", po);
# 1  pi=207'b000110011110000000101010101101111011110111011010100011000001110101111000110111000000111001101101100110011100000100111101011000110110001110111110000100111010111101011110111000111010000100001010010000100001100;
#1 $display("%b", po);
# 1  pi=207'b001011100010101001010001100100011001100111100000100111110000101011011110101111100100101000010000110111010000100000111100100011010110010110010001101100101011110000100001001000110011001100110000000011010101110;
#1 $display("%b", po);
# 1  pi=207'b011011111001110001001100110111010001101001010000010010100111001110001110110100100101000011110100011011111001011010100010001100011001110101110000011001111110111011000111111010110011111110110111011110011111001;
#1 $display("%b", po);
# 1  pi=207'b110100000011100100001001110110111110010111001000100010100110001001100110000011101010111101101111110101010101101110110010011101011000101101010101001011110010000111000100000010101110111100100010111010111000011;
#1 $display("%b", po);
# 1  pi=207'b111001110111100110011111110011100000110011010100001000001001100111001001101001101111110001101100111100001001100011010000101000011111010101011110000101001111010100010011111001101100010001011110110100011000011;
#1 $display("%b", po);
# 1  pi=207'b101011100010001011001110101111101001101011001101110111100010001110111110111011110010101110101111011011000000011100100110110110111111000001101100010110110000010101011011100100010110101100100011111001000101000;
#1 $display("%b", po);
# 1  pi=207'b100110011111011110101100001111010110001010000100100101011111100001111001000100011011110011100011001010001111011001110011001011011100011001111101001101110111010001101010110010111010111000000010010001111011100;
#1 $display("%b", po);
# 1  pi=207'b001101010100100100000011110011010100111110100011001111001010001110100111101010001100010011011001100110001001010011011011001100111011111101010111010101010110011010111001001011100100111111001011101010010111101;
#1 $display("%b", po);
# 1  pi=207'b000111100110001001010111110000010011011111010010111110110001011011100011111011000010101100011101110100001011110110000110011001001110000000111001010111000100000111101101111000100001010001110011010001001110110;
#1 $display("%b", po);
# 1  pi=207'b001110101011010100001101010110001000110010011110101010000001110011111010001110100001111011010101110000010111011000111100110110000000000111101011011111111111001010001010001010001000110000111011111111101010101;
#1 $display("%b", po);
# 1  pi=207'b111100101000001101110101000000100001000110000101010100100010000111011011111110010010000101110000000110101001100100010101011110001010111101010001011000011110100101010000110110111110110000110110000001011101011;
#1 $display("%b", po);
# 1  pi=207'b111101100000011111110010011111111000111110111100100111100010110100000110010010100100001000010110010100101110110101101100101000101101011111110001101111111111101011010000110010110110111010000000010000111111000;
#1 $display("%b", po);
# 1  pi=207'b100100001001000011101100000010100001111111110000010011101101011110000011100111001100111111011101100101100101100010101001100011010001100110100101001000001111101101010010111010010110111100110001011100110000010;
#1 $display("%b", po);
# 1  pi=207'b101001101011010000011111101110010100111101100101010010000000100011111010011001101001001010110010000011111000110010111110001100101011000000010111100101000011000111100111001101100010100001010100100001011101100;
#1 $display("%b", po);
# 1  pi=207'b111010001110110100001001010111100100100011000010000001111110100111001010100001011011000011010110110001000101101000110110110010111111000100100001100000000001100111000010110111001111011000001000110100100101001;
#1 $display("%b", po);
# 1  pi=207'b001100010011111010011111011101001101010010010000010100110000111110101011100101111111101100000010011011100101101100111100110000001010000001001001010011011000011100001001111111111001000111100101100101111110011;
#1 $display("%b", po);
# 1  pi=207'b011011111100100001001011011101100001110111110111100010110101110110000001001001010001100111111110011110010011000110011101100110000100111111100100100000001101110111001000000000010000111001011100100010010100000;
#1 $display("%b", po);
# 1  pi=207'b110110111110000101010100101101010111110000100111101001101011011111101101110001101001111011001100111100000001110111101010110000100101000110010010001111101001011001010101001010011101001000101111000001111100110;
#1 $display("%b", po);
# 1  pi=207'b011111011111000101111000100110010100110010111101110011111101110011110111000010011100111110011000110100001010000001110000001000010011001010010100110101100000101000001110101000011010111100010000001000000011100;
#1 $display("%b", po);
# 1  pi=207'b101000100001111111010001111101011110110001001000110010111000000101001110101010000001000100101101010011100110010101011010110100001101100001001000000110000010010110000111111001010000110000111111100100101111000;
#1 $display("%b", po);
# 1  pi=207'b000100110001011101100000101001110101110111000110010010000011110110111010101110010100110100101010101000100110010011010110111111111100011000001001011001111011001000000011000111100110001101011110011000111101010;
#1 $display("%b", po);
# 1  pi=207'b100111100101111110010010001110010001111001011000000010001111101101111100001101101101101000101100000001000001100110011001001011110101101101110101100101001100111100111101010100011001001100011101111000100001000;
#1 $display("%b", po);
# 1  pi=207'b100010110100001111000101110001011010100011000010011100110000010110100111011010101010111110111011011011101100011100110011100101111011100101001011010101101011011101011101001000001110101111001000100110110010110;
#1 $display("%b", po);
# 1  pi=207'b101110101110101000101100010010101010001001001001110001010001010000101011110110011100111100000100011011001011110011111010011111100111010101010001110110010000101010110110101010111111110001011100000101100111011;
#1 $display("%b", po);
# 1  pi=207'b100110110011011000110100001001000011011111011110110111010110011111110111110010100110000000111111000001001001001111110011010001111011111000101011111100101001001011011000001010111001101111111011100100110111011;
#1 $display("%b", po);
# 1  pi=207'b110111100001010101100110111001110100111000000001110011110011111010101100111100011110111110110000100000110110000001101111101101001001010001111111110110101011111111110000110011110110111010101011010101110001010;
#1 $display("%b", po);
# 1  pi=207'b001011101011001001101011110000101111011000111110101110110111110001101111101111000010111110110001001011000011101110101001101100011000001010111000110011001111010110011011010101000100000010001001000001110101010;
#1 $display("%b", po);
# 1  pi=207'b111101011010000101011100001100001101110010011101110010101000010100101110100001111111011101011101011001100011111011111010001111001001100010110101000111010001101010101111111100111100111110100011010100000111110;
#1 $display("%b", po);
# 1  pi=207'b001101101110100011110111000101000000110110100110011110001100111010011111011011011100100000001110101110000110100111000011001111010101111011011011110001010110100110000111001001101001101010100101101010001100110;
#1 $display("%b", po);
# 1  pi=207'b001101101011001101011010000111011000110001101101011100001101011011101111100111011101100010110001011110110000001111010010011001011000000011001110111001011011100011110101000111101111000100101000001000100011110;
#1 $display("%b", po);
# 1  pi=207'b111101001011000000011100001111010100110001111000011100000000010011001000010000000010011111110010001110111111101010111100111110110110011100010111101100010011010011111011011011110101101001110101110101011001011;
#1 $display("%b", po);
# 1  pi=207'b110011011110000110010110000110111001110000100110101011101111010110110110000111100010010101000000111001011001101010001101001011101000111111000011111000000100001011010111111110100011110111000111101001111001011;
#1 $display("%b", po);
# 1  pi=207'b111011001100101011111010100001110110100001001000111101001000011000101110111001001011010000000101101010100111101111100111010101111111000000111010011110100111000000010101101011110000101111101011001010010011110;
#1 $display("%b", po);
# 1  pi=207'b111101010011110000001010001000000001101110010001011111100100100000011100010010110000111110000110110011110101010110001100011010100010000100110110101010110111101111110111000101101011001100101001011110101110001;
#1 $display("%b", po);
# 1  pi=207'b011010100100000000111001010010110000001101001010001101101000001001111001000101100111001010010111110000100101000110011111111110001010111111100000110011000110000101011000010001000100010000010000101110011110100;
#1 $display("%b", po);
# 1  pi=207'b011100100101000100000000001001001110001011000010111000111000110111001100111011001100111011010001010111001111111110000011100101111110000000111110101101010111011100001111001000010111101011011010101010110111110;
#1 $display("%b", po);
# 1  pi=207'b110000000011001111011001110111011110010010110000010001110111111100111000101010000110011100111101010101111100011010101001110001000100010011110000010101111000000001011011000010010101111001111101011100010111111;
#1 $display("%b", po);
# 1  pi=207'b010110001111001000100101011100101100010010010010010111011010010001010000001101100010110000001111101110110011111110000010011101100011111100101001111001000111000001001010111001000100111001111111000101111010111;
#1 $display("%b", po);
# 1  pi=207'b000111111111001111000111001010101011011101111101000110100000011101101010001110111110100101010110011010100001100001010010001111000001000011000111111010110111100111101010001001011100001101100000010111001010100;
#1 $display("%b", po);
# 1  pi=207'b111111111110111100011101010110010011111001001100101111110011011111101001110011011100110010001000101111110101111100011000010101000101000010001111010011010110101010010111101101001010100111010011100100111001010;
#1 $display("%b", po);
# 1  pi=207'b101001111100101001101011111111101111000000010110110100010011110111101111001010000001011001100111001011000011000000101100000111111000011001011101111011000111011001110010000110101110101001111110100100100011011;
#1 $display("%b", po);
# 1  pi=207'b101010101111110101011000011000011010000010001000000110101100110111001101001100101100100000010100110001110010000100001101000000100001111101000000001000000100001000111010001010000100100101101110110010101001111;
#1 $display("%b", po);
# 1  pi=207'b010000101101011000110000010010011110111111101101110100000110101000111001010011001111010000111101111011011001110010111011100101100100011011100000110100010011001111100011011101010111111101111111010110010110000;
#1 $display("%b", po);
# 1  pi=207'b110101000101001011100111101011000111010101111011000000010101000001100101011011100111010110001001001101110101111011101101111100010011101110110110110010000010010011101110111001101011111111011001010001100011000;
#1 $display("%b", po);
# 1  pi=207'b011100001111010111001100111101101011000101010001000100000100001101010010011000100000000010011001010100100110011000100011011000101011100000000000001110101110010100101111001100110111010101000011000101101000001;
#1 $display("%b", po);
# 1  pi=207'b000111101001000001111100011000100001010110101100111011001010000100011000101111101000110001000100110001101010001010010001100111101100000001100101011111001010100000000001000100000101101100111001010101100111000;
#1 $display("%b", po);
# 1  pi=207'b010001101011111110010011101001010101011110100111101101010100110011100010010001000101001010100011101001101001000101100100011010010101110110010000111101110000001011001010010010110010001000000011000001010110011;
#1 $display("%b", po);
# 1  pi=207'b001111001111000100100111111111111001000111101011101100000000000011011000100001110101000110110000110010101000111110001010001110110011101001001110011101000010001101101100000101011011100001101101001100011110010;
#1 $display("%b", po);
# 1  pi=207'b001100010111111001100111000100111001001001001001101010100010100110100110001010111100011111111001010111001001010011001001001111111001110100111110100111111000101011001011111000011011100110100111110000111100001;
#1 $display("%b", po);
# 1  pi=207'b100000100000010001101001010001001110001001101110000011000111101011110011011000100100100011000001010001001000110110000111000110011011110001010101110001100101111000010111111000101001011101010011100111010010010;
#1 $display("%b", po);
# 1  pi=207'b110001101111100111101010110100001000011110110010011011101101000110101100101011011100000010001100101000100011110010111110011000010100101111011011001111010011111010001001100100010111101100110100101100001101001;
#1 $display("%b", po);
# 1  pi=207'b110000001000010110101000110110000000101101101001000011101001010111010001010100001000101100001111100110100011010010111000010001011011100101101110101100001100001000000111110101100001100101101011010010100001010;
#1 $display("%b", po);
# 1  pi=207'b111010110001111100100011100001010000100010011100110100001101100101011001111000011100011011011111001011111011001111111011011101111001011100011010101000111111100100011000110100000101010010111101111100000001110;
#1 $display("%b", po);
# 1  pi=207'b000101100010111000110110101111000111010110110100000110101111011011100000110010010110100010011001110100001110101000111101101101001100011101101100101110100010000011110001001010100011001001010000001001001000001;
#1 $display("%b", po);
# 1  pi=207'b101110001010011000110011000111101101101111000111011001101111011011000110011111001001010011000100000001100010101011111101001000100100001111101011111111101110011110010000000100011011001111101010010000001100001;
#1 $display("%b", po);
# 1  pi=207'b111010001100000011111010110100001001001011110011001001110001000100101001001100110100110010011111001110001110111001111101010101101110111001101010001110011110001110011101110111100101011111101101110010101000101;
#1 $display("%b", po);
# 1  pi=207'b111011000101110111011111001101111011001110101111001100001111011000111000101011111011111000100000011101000111000111011110110110111101011001101001011100000110001101100111111000101111110100010101100100001011000;
#1 $display("%b", po);
# 1  pi=207'b100000100100100111100100010010101011001110000011100010101001100101110101100010110000011010000001101010110111101101001101001111110011000111000000001100101001101111111110000110001111010110011100110011101100001;
#1 $display("%b", po);
# 1  pi=207'b000101001111110100101100101000110010011001110111010101110010000101101011011110100001111000110110101110010101101001010011111000111110101110010101000110100010010110000100111001000010001001011010111010010000010;
#1 $display("%b", po);
# 1  pi=207'b010001111000000101001010001010101011011110000111100110101011100011100000001101110000001000100011111011000111011000110011110000101010100111110111101000010001001000110010001001000100100000100100010000100000110;
#1 $display("%b", po);
# 1  pi=207'b110101110100111010000110100110010111010100010101101000100101101101000011101111100011011110000000101111010100010000100001101110011011110000011001101010010101011101011001101001100101110111001110111010111011010;
#1 $display("%b", po);
# 1  pi=207'b011101110110100100010110110101110101100010100101101000101100110011011100110110011011100101000000010010101100001111000011001010011101111000100111100111101001110111111101100110100100110101111100110111101011111;
#1 $display("%b", po);
# 1  pi=207'b100011110011011011011111101011110111011101011011000000010001101010011000001010011101000111100110110001001011001010001010101010011010000101100000000101111100000111101011111011011100101010111101100101000100111;
#1 $display("%b", po);
# 1  pi=207'b100110010101110011011101000001011110011111010001000010111111000011011100110100100001011011101111110010011010111001111011000110101000001000101011010111001111100101000101100100101000011101011110100010100011010;
#1 $display("%b", po);
# 1  pi=207'b111101101011111011111001000110010000010010101010011101001111011000000010000101000110001100100101110000101000011000000001100100101100100010100010101001011110111111111011001001110100101001001011101101100011110;
#1 $display("%b", po);
# 1  pi=207'b010010100110101010100001000000110100011110100011100110001101011011111010011110010011011111000110101010111110010001110000000101111110010101100010000111101010110110111110000101011100100101101001001100100111101;
#1 $display("%b", po);
# 1  pi=207'b110101101101011101010100110111101000001001011101111100111000001101110110010100010010111000010000101001000110001011010010000100111110000100101000011001100001011101010110101111101010101111011010101011110010110;
#1 $display("%b", po);
# 1  pi=207'b001111011000110000000101110001010101011110001110001000010100010101001000011111100000001100001001011101100010101000110100101001100011100001000101101001111111101101111001110000111100010110011110111010000101101;
#1 $display("%b", po);
# 1  pi=207'b011100101110100000100110100001001111001100111011000010101001000111000101001101000011101101110111110110000011001101000011100001010111101101010001000000000110000101001110000110001000000010101011011110111011000;
#1 $display("%b", po);
# 1  pi=207'b100101001101110001101011000010011011001101101111001001110000011001000010000011101001000000101001110000100000101100011101100010101000010110011010100001110001110011011010111000110001100110110011010101011010110;
#1 $display("%b", po);
# 1  pi=207'b100110110100111001101011001011010010111110010011010001010011001011010000001011010111100001011101001101011111111110010110101001100110011001010111001100101010011010010111010111010000101011101100011000110001011;
#1 $display("%b", po);
# 1  pi=207'b001001000010110001000111000010011000110011011110011100011101100100100001100111110000111001011011100110000000110001000010000001010000000010101110101000110010111111001100000001001011010011100111011110000011101;
#1 $display("%b", po);
# 1  pi=207'b111110010100100110010111100110100010011001101101011000110011011011101101011110100111110001000000111110011010001101111101001001010000100100111100110101111110000110010101000000010001000111001011110011011001100;
#1 $display("%b", po);
# 1  pi=207'b101001110110111111000101001000010010001010111110101011110011111110011111000001011101101011111110000001011001110111110010100100001000011000001001001111001001001000111101101100010000110010100000001110100010110;
#1 $display("%b", po);
# 1  pi=207'b000110000011011100100001111010101011001010111110100100101011000110101011100001010001101001101000011110111010111111011100011110000101101000011010001000001111111011110001011101011101100001101010001011001101100;
#1 $display("%b", po);
# 1  pi=207'b001110001010110110000100011111100011000000000010101001101101100000110011100111111100101011100011011010001101101110100001111011011010111010100001010111110101100011000101000001101101100011110101001110001100000;
#1 $display("%b", po);
# 1  pi=207'b000011001010101111110011101001011110111010111000110111101100010101110001001111111110001100110101000110011110010010100010100111101110010001000110111001101011011010101111111110010001000100010010010001101000101;
#1 $display("%b", po);
# 1  pi=207'b111001011101110110001100010101110101001010000110111000110111011101101111010110100101111000100110001010111001000110010011100010010010011100000100011010101101110000111111110001100110010001010100000010101111111;
#1 $display("%b", po);
# 1  pi=207'b110110010110000101111111000101110111010001000110010011000100001111010100010011010101011011001010010110010000000111101100011100101110000010101001111101111110101110111001101000110001111010011011110011010111100;
#1 $display("%b", po);
# 1  pi=207'b110001001100000000100010110101101111011100101010100011100001110011000100000100101011111100001100101111101110101111111100001000100011101110010011011010111111111101111100001001101101001100001111100101001100111;
#1 $display("%b", po);
# 1  pi=207'b001100110010111011011011010011101000100101110111111011111011100011100000010011111111011110011100101100100110100011011101001110110010110001111011100001000010001100111100010101011111111110110010010001101111100;
#1 $display("%b", po);
# 1  pi=207'b111101110011000001110010111101000101111000110111100101001010110001101101110011100000000011000101100111110111110100011001011101100110001011110100101001011111110101101110001111110010110011110010101110110110101;
#1 $display("%b", po);
# 1  pi=207'b010111000100011111111011100101011110100011101111010100101000011101100110010101101111001111111100101111110000000100111011101100000111111011011100111110110110111101111000110101000010101011111010111000100110001;
#1 $display("%b", po);
# 1  pi=207'b101100000011100011001100111010111111001101101001001111000111100011000100100101010011110000000000101100000100011101110001111011100100011001101101000000000110011010110111001111101010011101000100000110110110011;
#1 $display("%b", po);
# 1  pi=207'b100000000110111101001010111101101111110001000111101111111001111011010101001000101100111111100110000101110001110101011000111110010100100110110001001100001111000101111111001100110101001110100110111111111111110;
#1 $display("%b", po);
# 1  pi=207'b001100000000010100111101110110110110100110101011110101011110111100101101001111000100001110101011101110011001101110111111001011010101101110111100110110100111011001100010111001000111111001000110100101101001100;
#1 $display("%b", po);
# 1  pi=207'b101111111111101101001111111111110010000101001010110111101000001000001000101101100011100010011100101110111110010101000101101010001000000001111011011111000111111000000000101110010100000111101110010100010011111;
#1 $display("%b", po);
# 1  pi=207'b110100010010011100111111110011011100100100001100010001111111011100110001101010100100011101000011000101010000000101001010001100100111000000101110111110100110001110100111110110100010110000101000100111001111011;
#1 $display("%b", po);
# 1  pi=207'b101011001101100110110000111010001101001010010110110000100111011101100110101111101010000101100001000001011110001000001101111000101010001101010010000001000101110110100000110011000111010010000100111001001111001;
#1 $display("%b", po);
# 1  pi=207'b110000000011010011000111010000000111010110011100000011101000010001011010000001100001110000101011000111100100111100100100110110111110010110111000011001110100010000010111101011100010110011010100110001100011011;
#1 $display("%b", po);
# 1  pi=207'b001110100010000101001011111011111000000000000110011001010101100110110111010010111111110000001100000111110010001110011000000110111110001001010111011101100111101100110011110110010011100010000101111111001101001;
#1 $display("%b", po);
# 1  pi=207'b101011010000110101010111101110100101110100111111001111010001101000001101000101110101100001011000110110010000010010000100010001000011001100001111000110010010110001111000101010001010001110010010100010110001001;
#1 $display("%b", po);
# 1  pi=207'b100010000010011011011101010001101101001011011010111000111100000101111000100011110011100111101111011011011001001100101100000111111101110111001011001011011000110010101011011011010001100110001010000100000001001;
#1 $display("%b", po);
# 1  pi=207'b110011100111000101101010101100110011110001001111110000110110110000100100001110001000000001101000111010010010000111001011000000001100010011000101100100010100100100101010101111011000110001011010000000011111000;
#1 $display("%b", po);
# 1  pi=207'b110010101100001001000100011101101001100010011111111101000110011010110101111001010100101010110000001011011110000010001000101001110110010111000010100111011100001010101110100000011111100010100000010110101111100;
#1 $display("%b", po);
# 1  pi=207'b111000111110001110111000110011001001001000010110011001010110001111110111000011101101110110001000011111111111001101001111001110011100001100000010010111011111001010100011010001011010111100111101001000011011111;
#1 $display("%b", po);
# 1  pi=207'b010001000100111011011010011000101010101110101001010110001101110010010100001001010100100011011111100000101011001001111100100011110000010111000011000001100111001000111001100111001100100110000000111010000110101;
#1 $display("%b", po);
# 1  pi=207'b000011110110011010111001010011010111000100001100111001001001110010101010001110001000111001011000001011011010001100000011001000111101101101011001110010110011000001011000110000011111000010110101110110100000001;
#1 $display("%b", po);
# 1  pi=207'b101000100111001111001100010000000011010010011001111101101010110100000101010111101101001111010010101010000001001110110101101101011011001101110010000001101000110010010111001100000011110011111110001011111010101;
#1 $display("%b", po);
# 1  pi=207'b100100001110100010000011001011010010010111111110110111101100110110001001101111010110010100000110001101001101010111010100010011101011010110001110001010100011111100100001001010001010011101010110011010010010101;
#1 $display("%b", po);
# 1  pi=207'b111010001111010010000011011100000111111010010111110000101111111010000111100100101000000000011100110111111110011001100100101011001010101100101101100100001101100101111001110100110011101101111100000011100101100;
#1 $display("%b", po);
# 1  pi=207'b111110000111101101100100001001010101011001011011110011000001001011100111000110000101111111101111110001110001110000110110110101010101101001101011001001101100110111010001001011011010010111111011100001011111011;
#1 $display("%b", po);
# 1  pi=207'b110101000000010100100110110100011101111101001111101100111111001110001010011010001011001100100011011101100001001010001011010101110010101110011000001111001000001100010101111100010000110001000101010001010110100;
#1 $display("%b", po);
# 1  pi=207'b000111111111010011111100001111010010111101101001100011000000010000010011101000011000101000010111110101001001011101111111110010001001010101101010001110010100110010110110110110010011100010100011100110010001010;
#1 $display("%b", po);
# 1  pi=207'b111101101100001111111000100101100111111001100001011100011010101111111100100001110110100111111101001101001000110011111110011000101101100100101111010111011111011100110111100010101111011111011110010001101011001;
#1 $display("%b", po);
# 1  pi=207'b011001100111011100101000011101101101000110000101011001010111101011110101100100000010101100101111111000011000001110110100100111100101010000001001111011001101100010100101000111101010010000101111100101100100001;
#1 $display("%b", po);
# 1  pi=207'b111100010101111110011001110010101010101110101101010000110111011101010100011110011100010000101001101100110011011101010101001110100010100100001000100001000000000110110011000111110100101110111000100000010110010;
#1 $display("%b", po);
# 1  pi=207'b011110100110110011010110001100011111100110001001001111011110001101101011100111101010001101001111001010011010100111101001111111101111101101010111110000010111101010111110010010000100010111000010011000011011001;
#1 $display("%b", po);
# 1  pi=207'b001100000010111000111101000100011111011010010100100100111111011001001011001100001000110101101010110001000010111001100111001010100011111101110000111010010010010001101000001010000111011001000111001110001000111;
#1 $display("%b", po);
# 1  pi=207'b011000001101100100010010101010001011100000001001010100000100110000110100001111001010011010110001000110111001001010011111001011101000001000110011111011000101000101101011000011011111000111001101001101101101000;
#1 $display("%b", po);
# 1  pi=207'b000011111010000110100110110110111011011010001110001110111001011000000111001110100000010001111010111001110000110000110001001111001010000000000101000111011010110101110000100011001111011100000111011111101010000;
#1 $display("%b", po);
# 1  pi=207'b110100110110100001100011111010110010111000101110011001110101001000101000110000100011011000110100111101101000111101011111100000101011100101001101010101100110001001110000101110010010000011010100101010001111010;
#1 $display("%b", po);
# 1  pi=207'b110000100011011100100010010000110101101001010010111101111111100111010011011011100110011011011010010011010011110001110100111001000010100011010110011010000111011100101110001010100000100000011011110010000010000;
#1 $display("%b", po);
# 1  pi=207'b111010101101111011000011000110011111001001011100001101111001111110100010001001110100100011101011011110010101010011101101100011010100001010111101001100001010000001111000100111011100110111011111011101000110011;
#1 $display("%b", po);
# 1  pi=207'b111100111010110001000101010010010001010100101011110011011111100101010001101110011100000001000001000010111100111111101001110101000110100111001001011010100011011100001110111110110001000011100101010000111010000;
#1 $display("%b", po);
# 1  pi=207'b110110011010001001110111111010001010011110011100001101100110100011100000001001001000101010101101100111000001011000101010001100100010001101111101101110111010101100010000000011111100011110100110100110100110111;
#1 $display("%b", po);
# 1  pi=207'b001101101001100010100101001000111010001111011011010000111111001110000010011001010001110011100111000000010110010111010000000111010100011111010100101001010110111101111010100010001101110101000011110001101100100;
#1 $display("%b", po);
# 1  pi=207'b101011001110000011011000000111001001011100001010101011101101001111010110010000010100011101000100110001001001110010101100010110010001100111001110101100010110100101000010010111101010011110011110011000000000011;
#1 $display("%b", po);
# 1  pi=207'b010111011010000101010110111001111011000001010010110001010101001010001001001111100010111010101001111000011011101010111110001101100010001111010100010011100001100110101011011101100101001111110111100111101100100;
#1 $display("%b", po);
# 1  pi=207'b010101101000111001101010011011010010010010111010010101000100100000010011110001011001000110100011010111110011110101001110110010100000110101101011011111010000101110110100001110011010101010111000111101101100000;
#1 $display("%b", po);
# 1  pi=207'b111011101101010010010000001001100000001010010100000011101010011100111100010000100010100110101101111000010111000000100000011100001011000111100010011111100101001000010000011011110110100111110101001100010010010;
#1 $display("%b", po);
# 1  pi=207'b101101100001010101111011100001101001011101110000101101011011101010110010010101000110000001001110111011111000010001000110011111111110001010101101100010101111000010011010111100000110010100011110011101011101000;
#1 $display("%b", po);
# 1  pi=207'b110100110111110011111111010011010101000100110000111001101110110010111001110111110001111001101010101010100001010010011010100000011110000101011000100001001000111000010011001000101011000000111001001000101001100;
#1 $display("%b", po);
# 1  pi=207'b101001010011111010011101110110101010110010111011111001010110111101011111000011010011000110101100010101101110010010101101000110110111010001001111100000111011110110011100011011111101101101001000011100110001110;
#1 $display("%b", po);
# 1  pi=207'b111000011111010100110000100101111110010011101101001011000101000110110100110001110011100011001011000111000001100101100011101011100001111011011010100111000000101000111100100000000101000000000001111110000111001;
#1 $display("%b", po);
# 1  pi=207'b000101110101110100101100101101110111110000101000110110011000010001000000100001001000111110010111101000110001111011111100000010011101011011010100100001111111011110100011100101100010011010011111011010010001101;
#1 $display("%b", po);
# 1  pi=207'b000010110111100000100000010110001010010111001011101100100000101000010101011100111100011011110101011111100101011010110110010101100000001010111111110010111011110010110000110111111000110111011010010010010111110;
#1 $display("%b", po);
# 1  pi=207'b100001001011000001000110010000111011100101000011000000000011100110100110111010010111000001000110001111101010110100000111100011100101001011111110111000100100000101111001000011010011100101110111011110010001101;
#1 $display("%b", po);
# 1  pi=207'b110010101101101001001001010010001011101000101100110101000001001111000101010111100000111000001001100000010101100001011111000000100000011110001000001111001010111011010011010010110101100000010101101100010101110;
#1 $display("%b", po);
# 1  pi=207'b011100001111000000001000001110010010111110111101111100100100011100000111011011111010100101100111001111011111010000000101101010011101101010111000111011111000111100001001101100110010100011111100100010010010011;
#1 $display("%b", po);
# 1  pi=207'b000111101000110100001110001111010111110011001100010100111100101001100110110011110110010110011111101101111001111111100010111010000110001110101000011011011110010010001000111000111010000011010111001100001100100;
#1 $display("%b", po);
# 1  pi=207'b010000000000100000111011001101000101100000010001101001111101100001110001010001011111111001101110101111111110110011111100101111100111101001111101000000101101011010111000111110110110101110100000000101101101001;
#1 $display("%b", po);
# 1  pi=207'b000100010011111011011101001111111101010100101111110011101100010110111101010101111101101001001010110110110011100111100000100111001011010101011110000100010100101000110101001000001110110110111011111001101001011;
#1 $display("%b", po);
# 1  pi=207'b101101000011101110111110001101010110100110100101100110100110110100110110010011001011111001110011110010001100101100001110101110110111110110110101001111001000010101101100000001110000001101101011010010100011111;
#1 $display("%b", po);
# 1  pi=207'b010000000000101101100100011111111010011001111010010110100001101000101111000010110100011110011111101110010001100001011111001111110110011101110010000111001000111100100010010001001000110010001010101011100010000;
#1 $display("%b", po);
# 1  pi=207'b110000001001011110000011010101010101010111100111110011100010010011101000110000110100111010110111100110011010101101011101010010100110001100100111100000101011000100110111100100000010110100111011001000000010100;
#1 $display("%b", po);
# 1  pi=207'b100110100110101001001100010010011101100011101010010100011110001100000001110000111000011011000100110000000011010010011001110011011111101100100011000101110001010101010110110001111111001101010010001100010011001;
#1 $display("%b", po);
# 1  pi=207'b101011101100110110000010101110011100001100011110100100101000010111100110010000001110001000111000000100000011001001101001010011010110111011010010010101000011000111101111010101101101100000101011110111101111001;
#1 $display("%b", po);
# 1  pi=207'b000000011000101101110100111001100101101100101100001010101010000101011111000110111110001101101110101110011101111010110100010100101010000101100010101110100100111110011001110011111001010110110101111011010100111;
#1 $display("%b", po);
# 1  pi=207'b111011011110110101001000100111000100001100000110100100010100100110010001010101111011000011101001010001011010100110000010111100011011000001011111001000110010111101101000100010100100000001011101110011010001111;
#1 $display("%b", po);
# 1  pi=207'b001111011111000101011001110010001100011100110011011100001100100010000100000001101000001100101110100001110101000100001110111010100001011000111111101011010111001011110010000010111111111101001001101001000000110;
#1 $display("%b", po);
# 1  pi=207'b011111101101010001111111011000010111010011110010111110100011000110111110111010011100010010111101111010101110011001001100101000100110100001000110011010100100000011100001011001001110010010010001101100000101000;
#1 $display("%b", po);
# 1  pi=207'b101101100000110000101101111011000001011110101110100110100011110111101110011011001110011100100100110100101101110011001111111001010011100001011111011111001101011001000000000100110111010011100111011111101011011;
#1 $display("%b", po);
# 1  pi=207'b100110000101110000111001011001100111100010100100001001111111110100010011000100100010110010111101101001000100001000100101110010110110011110000100001010010000011010101101011001101010010010101111000000101111001;
#1 $display("%b", po);
# 1  pi=207'b100101000000011011011011000010010101001110010101101111101100001011011111101011010010011001000001010001111100111011111111101011011110111111010101100100100010110010111000001011101101110011110111011001010111000;
#1 $display("%b", po);
# 1  pi=207'b100110010010001011111111100010001101010001000111100110001000110111111110111000110111101101100111111000011101001000000010000110001011010111100010110010011010100110010111111100110110100110101010001000110000111;
#1 $display("%b", po);
# 1  pi=207'b101101011110010001100111110000100100110011100001100111001111000011110011110001010100111110110111110010011000000100100101110010100010110111000001100100000011100001001101000001011100011011100100101001001011100;
#1 $display("%b", po);
# 1  pi=207'b010111101111111100001101111010110110010001111001101101111101011110010010011100000010110111010011110110100101011100111010100100100001101000110110101010000011000101101111010111011101101111110011110010000101001;
#1 $display("%b", po);
# 1  pi=207'b111011100110000110111000111111010100001000101111101100011111100000110101011110111000011110111010010111101010010111010111011111001011010001000100011001111011011110000100001011111100110000010000011011101100000;
#1 $display("%b", po);
# 1  pi=207'b000010001011001011001110011110000101111110101011111110010001010111110001101100101001100110011100100001011111100000101001000011110101101011101111011010011110010001111001111000000011101101101010111001011101101;
#1 $display("%b", po);
# 1  pi=207'b010011110110010001110111011101111010111110101110111111100010101100000011101010000111001110010010100000001010110111101011011100111010100001100101110100100010010100011011000011010110111100011000010010001110011;
#1 $display("%b", po);
# 1  pi=207'b001101001101101110011110100010011100010100101110100000111101011110111101000011111111011011110110111100100111101100001101110011101101110001010100110011100111101000000100011110000111001001011001000100011000101;
#1 $display("%b", po);
# 1  pi=207'b010011001111111001001001110101000111110100101111111001111011111111000000001000110011100101101111011010111110100001110011001000111101000101011100101100000001100100100011100111101010101010011011100000101100101;
#1 $display("%b", po);
# 1  pi=207'b010001111000100111010110000010101110100010001101001010010100010101011000000110100000010010010101001111010110001100000101110010010001110010110000110011011100011001100111100101010010010010100010001100010010000;
#1 $display("%b", po);
# 1  pi=207'b011100101101111010111111000111101001010110000111111001101100100110111010111101000100011100101000000011000110110000111011110100001110110010010100110101000010010011101000110110000111100101111011010111011000000;
#1 $display("%b", po);
# 1  pi=207'b011001011010110101110011010101011111000100111001011000011101110111111000010110001111101111001001110111111100111000001100010000100101001111011010010001010110111000011100111101111010110101011001011110100100100;
#1 $display("%b", po);
# 1  pi=207'b110101000100100111110001000110010111001001000011101100000110101010110101111100101101011101100000000110110001010000000000101100101000011110100001100101100010101100101111110111110100110101001001101111001111001;
#1 $display("%b", po);
# 1  pi=207'b011000101111000110100110011111100001111101110000100100100110010100111101001111001111011011001100100101111111011101000011100011111000000001100001010111111000001110010001001110010111101000110000010100101011011;
#1 $display("%b", po);
# 1  pi=207'b100011000000001100010100000100100010001101111101110001001010000111000111110110100011000010010010111001001111000110101010101101000100010000000111010101101101011100101110101011011000001000011100110100011011101;
#1 $display("%b", po);
# 1  pi=207'b101001001011100110001011111110100011100111111000101110011100110010001010101110110100100000001101011011110100010100011000100001011100011011110000110100000000000101110010000111101001000000111100000101010111111;
#1 $display("%b", po);
# 1  pi=207'b011011100010010000001111000010110110111111001110101100100111111010000011110011011101111111110101010100011110011000000001010000000100110001010011101001101011000011011000100010110000000000011011001110101000111;
#1 $display("%b", po);
# 1  pi=207'b011010110101111111100010011011111010010110001100110110011010010110010010000010110000100001011001001001011111000111100101100011100111110001110100000010101001111110100001111001000111110010001001110011000001100;
#1 $display("%b", po);
# 1  pi=207'b010000100110100010111000110001111110100101011110111100011111101100100110001010011100100110110100001111001001010101001101100101000111011110111011000010110100011010110011110111111101011000000100101010111101101;
#1 $display("%b", po);
# 1  pi=207'b011101000110100100110111000101100101110111001111100011111000001100001110100000000011110101110001010000110100101000000100010011000111000010100000101101001011001011101000101001010111001001010111000000110111011;
#1 $display("%b", po);
# 1  pi=207'b111011011101011011011110111001010010010000100111101001010101100101001000100011101001010001101000010000000111111101100111100010011100111010010100111111111110100100000010011111111000010000011011000001011010001;
#1 $display("%b", po);
# 1  pi=207'b010101010110010100101011100010110110111000011101010001110110000100101100011110100111110110011100110000101111001100110101001011010101000101101111010110111110010100110001110001101110100001111010110001100110010;
#1 $display("%b", po);
# 1  pi=207'b111011111001100101100010100101000111111101001111100100111111110111001001011001111101111010000011010011101010111001001101001110010110100000111100111100001011011110001100000010010110110111101000011101100100000;
#1 $display("%b", po);
# 1  pi=207'b011111000011111100010001001011001110110000000101001100111101000001011010010100001010000110110001000111010000110001101010110111011101010100101111111010111111111000000001100010011000101110111110100111011000010;
#1 $display("%b", po);
# 1  pi=207'b011100110111111001111000111110111100011110101111000010001100000001101111101111010100100110110110100001001110101011011001110111110101000000010000101011000011111000011111010011010111001100010000001000101011100;
#1 $display("%b", po);
# 1  pi=207'b101101110000110001010010011110010010100010101111001110110010000000101000111100110011001101101001010101111101000110011111101111000100101111000010010110011101001010000110101001110111010000000001011110010011101;
#1 $display("%b", po);
# 1  pi=207'b000101010001011110110110001001101100100000000001110010110000010100111101110101001001001101110000000011000101111101101000011000100100011100101110001110100110101111100101101101101101000001010010101111111011000;
#1 $display("%b", po);
# 1  pi=207'b001011101110110011100101111011011110100101100000101011111111111111100111000010011101000100010100011011010101001111001011101010100011000110110001100110100001111001100010011110001011001111110101111110011010110;
#1 $display("%b", po);
# 1  pi=207'b010100000110101111000110100001001001100110001000100010000001001001010101011100111100111101001010101101111001101000011100110100000111010001111101000010111101000000111110011001001010010001110100011111011100101;
#1 $display("%b", po);
# 1  pi=207'b101111011000011101011100011001100110110100010010110111110000010101101001001010001001100010111101100101010101001000110101011011101100011010110010001001111010000111110000111010110011011000010101011000101010000;
#1 $display("%b", po);
# 1  pi=207'b111011011111001001100110101110001100011100101011011101011011111101010110001000110000111011010000011110001001100100100100011001010000000010001000100010100001100010010001000001111100111111100001011110111101001;
#1 $display("%b", po);
# 1  pi=207'b011011101011011010010101101001110110001001011011000100101100010100111011011111111110110010010001010010100100110110000110101010000001100111011001100100101010000101110010101101011010100010010001110000101100011;
#1 $display("%b", po);
# 1  pi=207'b000000100001000111000000001110001100010101010111101011101111101100001101110111000101000001101101110011100100011111000001111100010100101101100101110001000110110110111010000110101001010000111010100110110010101;
#1 $display("%b", po);
# 1  pi=207'b101001000010111100011000100000001101110110110100000001100100001010110010011010100111011010110111001100101000000000010101101101000101010111000100011001000110111001000001100110101111011010000100000000011010101;
#1 $display("%b", po);
# 1  pi=207'b011100000100101001010010100000101010001101010101110100010000000011010101111100011100101010100100111010111111110001011001000000001100111111000001110011011111100111110100010000111100111111011111010011101001000;
#1 $display("%b", po);
# 1  pi=207'b110111000110010000001001110110101011110010010101000110011010011010010011110101010111110110110111011010100110110001011101011000000100100101100101110011100011100001001010001011010010001001010111000000010001111;
#1 $display("%b", po);
# 1  pi=207'b101010111110111111000110011110100011101100111110110101100000010011011100110000010010101101011010000001110101100101011000011101101000000000001010111011101111111010001000111110100001010000110110100001110011010;
#1 $display("%b", po);
# 1  pi=207'b001100011001110111110010000011000101101110110110110001110010110010101001000011000010000011001010111010000011111101001000011001000110101010000001110111011111111101001000100101010110011010110110111110101100100;
#1 $display("%b", po);
# 1  pi=207'b000110001110111101111010000010110001110100000000011110011100101010111000111100000110001101011000011110101110010111111011100100010001110100110011001010111010110111001010110100111001110100101111101011101010100;
#1 $display("%b", po);
# 1  pi=207'b111001010011100100010101101101111011001011011000111111110000100010000111111011110110111011011010111110110011000011011100001011000001111101010001010011001111111010111111001000011010010000111011111100101011000;
#1 $display("%b", po);
# 1  pi=207'b010011111110011100110010010101100000100010100100010000010111101011100000111010011101000001011100001001000111110110010000111100010010100011011010011100011000111001101100001101111111111110011110100010110000010;
#1 $display("%b", po);
# 1  pi=207'b011111011000001100010000001000110111011100110111100101100011001011100000101101000100011010110110000110010100100001001101110011010110100001111001100110100100100010101100111011001010111110010101101010100011011;
#1 $display("%b", po);
# 1  pi=207'b100110011111000001110111110010010001111001011100100000101111000101111011111110101111101010111110111011010111100101010110000110111000010011011101101111111100111110100010010011000101011011011101100001100001111;
#1 $display("%b", po);
# 1  pi=207'b100111010110110011100100000101001110011111001011100111110001110100100011000110001001010101011111011110010001001010111110000010100010101000100011000011010101011110011011111011011110000100111000111001110110011;
#1 $display("%b", po);
# 1  pi=207'b101011000010110111010111001110100111110101101101100001110000011011000111100111101000001100101111011001001101110111000000011011000000110000111100001101111110100010110001010001100111101000111110010000011001011;
#1 $display("%b", po);
# 1  pi=207'b000100010001010111100110011011110101000100001010001010010111010101110101000010111101010111011001010000011111000111100011000000011110100110000010101010011010111011001100000011111110100010111100011111101001111;
#1 $display("%b", po);
# 1  pi=207'b100110111010001101001010110001011111001101011101101110000010011000001000111010001111111110011010101110001001101111000000011100001011100011000101111100010100011000011000100000001011100001000011100010010010110;
#1 $display("%b", po);
# 1  pi=207'b111000101100000001011000001101010000001000010111100011110101111111011101010101110111000010101010111000001110110011010011110101100010100010110011100111100100111011010011110000101011111111100110101101011110000;
#1 $display("%b", po);
# 1  pi=207'b111011010011110101100010100111100101100010101010100101011111001111101011001010011011010111011110000110100000100110101001010100100010011111011000110000000001010010001100101111101101000010100111001100001101000;
#1 $display("%b", po);
# 1  pi=207'b100000110001110000011100111101010111010100001101011101100101010101000110110110010111000010010011011010101110110101000111001011010110010000011100010101101001111110110111011111010011100011101100111000000111101;
#1 $display("%b", po);
# 1  pi=207'b011011111111100111001000111100100011101110010101010110000100010001111110111110001010101001111111001111110100000110011010000000100100010101100101010100101111100110100001001011000010110011110111010011000101001;
#1 $display("%b", po);
# 1  pi=207'b111111111010111111011010001111011111000101001100010110111101000001111010101010000001100101001000010101011011001110011000000111001010000011000001000011011101010100101101111101010011111000100101010000001000001;
#1 $display("%b", po);
# 1  pi=207'b011110101001111100010101111000011101001010001010011110001011111011111110011111100111000010011111110000101100111000000010010011010101010001010010001001000001100110101001010011111111000100010010111000010100001;
#1 $display("%b", po);
# 1  pi=207'b011111001111110100111100011111100001011010000010100010000010001100011011001101010000001001101011111010111000010111101001111010101001011000110001111010010110100100100010010011111101010101111111001111011100000;
#1 $display("%b", po);
# 1  pi=207'b110001110110001111100101111010100100000101100110001110110011100110000110010010111110111101101010111110001101111001011001010000001011001111001000000011110110011010011111100110100110111001001001111011001111001;
#1 $display("%b", po);
# 1  pi=207'b001000000001010000111110100111011000101111101101010011011101001101011100000001100101001100010000100001011011110010000101110111011011000110101111111011110001100110111100110100110111010110100100100011000110000;
#1 $display("%b", po);
# 1  pi=207'b111011111111000001011100110111110100000111111110111101011100101110100100000100100001011111110000101001000010011000000010011000011110111101110000000110101000000011010110010110101010110101111110000111110001000;
#1 $display("%b", po);
# 1  pi=207'b110111101111000111010010100100100111110001101110001100110001010111111001001001111110110110000100000000011101011101011111001000001110101100011001000110111101011011010001111011111010110011011000011000101010010;
#1 $display("%b", po);
# 1  pi=207'b000110101011000100100101001000001001100101011100001001001101100010101001111111010111111100110010000110010011001011010100011110010000110111010010110100110010010011010101110101010001011111100000000010001101011;
#1 $display("%b", po);
# 1  pi=207'b111101111001011101111010011110101101110111101100100010111100010010000101101101011000111111011001111010010011101011010101101110110101001001000110011110011101001010100001000010100001101000000000001001000100011;
#1 $display("%b", po);
# 1  pi=207'b111101001010100110111100011111101100110001000011010101010110110101110000000000110001011010001000100110111001110100011011011100101011010110001101011101111011011101111010001010111010110110011110010111110001101;
#1 $display("%b", po);
# 1  pi=207'b010011000000100001101110100111101001001011000001110010001010101000101111010111110001000110000010010111101111011001000101011011001110011000101100000111101111001101010111100101010100010010100001101000110011010;
#1 $display("%b", po);
# 1  pi=207'b101100001001001011000000001110001101001011101111011100111101011110010000000011101001010000011111001010101111010100000100011101000011111011110001110110000000010100011011101011011100011010001100001011000010010;
#1 $display("%b", po);
# 1  pi=207'b000101001010110111000010100001110111110000110101101000101110111010001010011110010010110111000011111111100011011110011010101111111100010011001010011011100101100001000100010001010000111101010010000011110001101;
#1 $display("%b", po);
# 1  pi=207'b101000011001101110001011110101001001101100111011111010101101100010001011101110100010011010010010101001101011000011001001011101000010110011011101001001110111101011110001101001100111111011010000000100000111100;
#1 $display("%b", po);
# 1  pi=207'b010111011000010011001110100010101101111110100000100111001100101010011110110001010100100101110100111010101000100001101111001010101011100000001010110001001011001001010110101000010110100111111000010010000111010;
#1 $display("%b", po);
# 1  pi=207'b011110101001111010100000110100110110111001010001111000000111011111101100001101110010101010011100111000101011001100001101000100110100001110100001000010010111111001100110001001010010010011000000011101110001000;
#1 $display("%b", po);
# 1  pi=207'b010001101001101110011000101011010001110001000111100111010011000000101000100101101100100010000001111110111001000000010001110001101011000100101010001100001110100011110011010001001100010111101111101010011111010;
#1 $display("%b", po);
# 1  pi=207'b101010011100010110001110101001010111100011010010100110011001111011011000001100000010000000000011000000010000000110001011001101110100000011111110110011111100001011010000110001001011010001111101111001010110101;
#1 $display("%b", po);
# 1  pi=207'b001101110001110010110001110101011010011011011100110010111010100000000100010000110011111111001011011010011010110010001011010011110111001001101111100100010111010111101000001011110010011000011111111001111101100;
#1 $display("%b", po);
# 1  pi=207'b111010001010001101011101101011110001000111101100111001011100000001001010110011010100001000111000110011110010000100110001110000101111001010000110100011100011011111111000110100010000111110111111110110100101100;
#1 $display("%b", po);
# 1  pi=207'b100111011000100001011011000100110110001101011110000100100001101000010111010011000100101111010111111010010111010010000001101001010011111010110101100111000101111111000100011110111100100111000110001000100011011;
#1 $display("%b", po);
# 1  pi=207'b000110111000100110110011110001010010011111010111111101100010000100010000101011011000001110000011111001100101001011100001110110000101101110110001000101001110011111000011100001101111010001101110100110011000110;
#1 $display("%b", po);
# 1  pi=207'b011011111100111001111110101001001101100001101100000101110011110111001010111001110111000001001010010110101000111100001010000111010111111010000100011000101110101010101110100110100110101011111110110111111000000;
#1 $display("%b", po);
# 1  pi=207'b110111000000100011101000000101100100110111011100010010001000111000001001100001100001000010010110001111101110010111011000000110011110101001011011101100110010011000110110011101101011101110011011010011101111100;
#1 $display("%b", po);
# 1  pi=207'b101111111101110100101000010111110000001001011011000001101100000000111000100110111011001110111110011001100101001001101101001111011100000001011001101110001011010000001001000111010010100111111100100001001000100;
#1 $display("%b", po);
# 1  pi=207'b110011101011000101101011101011000111110011101001101100100000000011011101101111001010111000010110000100101111111101000101010010110001001110010010101111101000110100010100110100110110010100010010110011000010100;
#1 $display("%b", po);
# 1  pi=207'b010010101000001010001100001101110010111011011011101100100111011001011111110110000101000000000100101000110001000110101010001010010100110111110100100111110001001011001111011001001001010011101011100101001000111;
#1 $display("%b", po);
# 1  pi=207'b101111011100100000101111111111001011111101111011011011110001011101011100101100100110011111011101010001111001001100110001010000010111100110101100101100101100101000010111011101110011110100100110100000100110010;
#1 $display("%b", po);
# 1  pi=207'b001000100001100100001110111010010100001101011100011010101010111000110111110101100100110111100100011100000010111001110011010000000101011110111101111110100011001110100011110101010100001001110011101100111100101;
#1 $display("%b", po);
# 1  pi=207'b100011101011100111011111110011110100011001111000011000001110001111011011111111110101111001001110011100101010010001100101111011111011110010110111110000101110110011110100010111111100101111011011100110110101011;
#1 $display("%b", po);
# 1  pi=207'b100111010000000110000100000111011111110001011101000101001001010110111110100010000000011101100111100100001000110101100101110111100111010101011111100111110000001010100101111101110110000010000111000000000001110;
#1 $display("%b", po);
# 1  pi=207'b111111100011011110110101111011000011011100101100010000011000101110001101011101101111101100100000111001000101101011001101010011111000110111100111010000101001100010000001000101110110010010110010110011011100010;
#1 $display("%b", po);
# 1  pi=207'b000000010101001100111100110111010011111100011000000001110110110100101011111011010001100010010101011110001001011000110101001110010100011111100010111010001011101011000000000011010011001110001011000110000100100;
#1 $display("%b", po);
# 1  pi=207'b101101100010001101000101001100100111100011100000111111110010100111100001011100001110110111111111010010101000110010100111110100110000100101011010101110001100110011011000001110110000010011101011001111001110000;
#1 $display("%b", po);
# 1  pi=207'b111000001100111000110100100000010001001011111110110100011001010101110010101111001010100111111101011001101010101101100100001001111111101101111000100010111011010000101111100101001001110010001100111000010011101;
#1 $display("%b", po);
# 1  pi=207'b110111110010100010000101110011001000001101001010101001010001000000100000001011000000001001100111011001011111110111011101110000001100101011000011110001110011100111000011111010101011001000010000000001000110011;
#1 $display("%b", po);
# 1  pi=207'b110110011000100011111101000110010101100010000010000010111011000000101000010010010110010110101101010101110101000111100000100111101100010100011011100010101100010100001101011101111001110010010010011101101011010;
#1 $display("%b", po);
# 1  pi=207'b111101101101001111111100011010100101011100000001100111001011010001001101100100110000110000110101010101010101111110000000011010000001001011110011100100100011111101011001011101010100011001000100110111110000111;
#1 $display("%b", po);
# 1  pi=207'b000001000000101010000110010101110000100110010011100000111000001111000111000100001111111010110010101010001111001010011011110010110110010101011001111110000010111101110011000100110001001000001110011010001111111;
#1 $display("%b", po);
# 1  pi=207'b111111111111000101000101111100110100100110011111001001010101101100011101001111110010101100101100010100100110000111010011001001111011011111010100000100011001111101111010010110100001110011000001011110000000001;
#1 $display("%b", po);
# 1  pi=207'b010011010001101101111011000110010100110001010000001111100111011011001110100000110010010001101000111000010101011000110101001110010100000101010101011110000011100100011111111011110010000000000000010111101001100;
#1 $display("%b", po);
# 1  pi=207'b001111101001000111101101101110100001010011011100100011110101000001000100010111110110000001101110100001000100001101101101000001001011001111100010000001110001100011011100000000110010000110011010011101100011001;
#1 $display("%b", po);
# 1  pi=207'b110101101101100001110011100110100001100101010001100100011101010100001010100110000000010010001100110000111011111110110001010110110011011011101111010001010001111111010000111101010100001001111100101000010011110;
#1 $display("%b", po);
# 1  pi=207'b110011011010001011011101101001110111100010011000010010001011010111001010001001010001010001111101110000001111001001101101010100001000100011000011110001100101010011110011101000110111000111010011111010101011101;
#1 $display("%b", po);
# 1  pi=207'b010110001000101000110001110000110111111110010110110101110101001101011100110100100000110000111001101011000001111111000000101111001010011100010000010110111101011000101100000001101010000000110001101101110110111;
#1 $display("%b", po);
# 1  pi=207'b111110101101111111011101011011010100000010011001110001110001001101001011011101010011101010011110000001101111111000110110110010110111000010001111110001111110010100010010011101101111100101011100011001011100101;
#1 $display("%b", po);
# 1  pi=207'b110011101010011000010111111011001100010110100101000101101001111001100011110110000100100100101110110100101001100111101100010111011011111111001111011100011010010000000011100000001000000100001110100110010010010;
#1 $display("%b", po);
# 1  pi=207'b101101010110000000001010101101000000101100111001111111011011011011110011010010110110100110001010101110011000011010011000111100001011000001010110101010110111010011010010001111000011110011101001111111011011101;
#1 $display("%b", po);
# 1  pi=207'b110010100101011001110100101100111110001110001100011010100101100110001110010010101111111100110011101100011100111010010010110100010110010110011010010011000001000010011111011110111010001001111111100000111101111;
#1 $display("%b", po);
# 1  pi=207'b010011000100101010110101011010111101001000010000100011100101000001110010101000110000010110111100110111100101001110110000101011001010010010011101010000010100100101000101101101110111010111010101001001101011100;
#1 $display("%b", po);
# 1  pi=207'b010110110010001101111101111100110010001111101001110100101100101101110110010010011110110010011001101001111100111000000111101011000001000000011101111010000100110110010010011010010100001111110000100000110001010;
#1 $display("%b", po);
# 1  pi=207'b111010110110110011011101000001000010001010011111101000001011011100101010111000010100000011001000101010010100001000100010011010011100001100101100110001111011000001011010100100101000111000011110001111010101110;
#1 $display("%b", po);
# 1  pi=207'b011110010001110001111101001000111000101001110010001011110000010101000100110100000101100110010011011001011110110001101110101011000101111110101010001011001100000111000010110101100000011010000111100010111111101;
#1 $display("%b", po);
# 1  pi=207'b011010101011101001011111001100011011110010110100011011011001111100001110001110110111011100010000100101110010111110011100001011101000000100110001110010001000100010000101110101000001001001011101011111100010011;
#1 $display("%b", po);
# 1  pi=207'b110010101011101101010010011100011110111000001100111100100101111110001010000010010010100011100100100001001111111011110101001110011000111101111111011011001001001001110101000100001010001010110010000010100011001;
#1 $display("%b", po);
# 1  pi=207'b000110011110000110011010010101101011101101010101011100100010110110100010011101010111011001001000101011101010101011101101011010010011101111010000001000000000001000110111100000100110010101010011100100000010000;
#1 $display("%b", po);
# 1  pi=207'b000110111100000101101000111100111110111010111111111110001110100101111010111001101011111001000111101001110010111100010111111010101111110110011000110110100001100111010101101001010010011101001011111111000011100;
#1 $display("%b", po);
# 1  pi=207'b000100011011001100011000010111100111000010101001011011001001011100010110011101001111010101011101010011100000110011100111000010110101001001100101111001010010010111001000100110000011110101001111110100000100001;
#1 $display("%b", po);
# 1  pi=207'b000101110100110111010110100111110110111000000001111000001111010001111011111001011101011000101100110011111001010000001101111011110110000001101111000010100111101110010110101010000010111110100010001000010101000;
#1 $display("%b", po);
# 1  pi=207'b010001010110011110110110000100100011001000110010001101101010000110111011011111011110000010110001011011000011100100111100000010001011100010100101110100001010100000101010001001110010111001000110101110010110001;
#1 $display("%b", po);
# 1  pi=207'b011001100111101110101110010101001001111001000100110111111011000000101000001000110101001101011000110110001101011101111010111001100110010011111010010011001001101111001010111011100011111010010100000101110000001;
#1 $display("%b", po);
# 1  pi=207'b111011001101101100101110000100000010010000111010011111110010011100100101100000110110110101010100001011100001000000010011010111010100010100110010111111011001000110000010101111100010111001010111000011011010011;
#1 $display("%b", po);
# 1  pi=207'b100001110010100001100110011110001001101111000010010101001010100001000000000010010101100100000011001101000100011100100001010101010011010110110111101110010010000011011101101100000101100001011001001000110000100;
#1 $display("%b", po);
# 1  pi=207'b110111110011001011111010111101100011000000001110010001100011100001111000100011101001111001110100101001000001011111101001111000101110011101111011011000110011101011011000000110011110110100010111110000101000110;
#1 $display("%b", po);
# 1  pi=207'b010001100110101011010011011110011110111000000110101011001011111010000110000000100110010101010011011110001010011001110101110000101000100010011100010111111101100001001110100110001110001010011100111011001001011;
#1 $display("%b", po);
# 1  pi=207'b001111101100010011111001101100011000101000110001101100001011001101011010011011100010100110100101010010110110000000110111101101000110101101110111011011000011110111100000010010111100100110101010101011010011011;
#1 $display("%b", po);
# 1  pi=207'b010011110010100001111010101001111011110101010111011010011101100010011101110000110101100011101011101111001101000000111110011000010100001101110011110111110000100101100001001111101001101111111011111000111001011;
#1 $display("%b", po);
# 1  pi=207'b101011101011101011110100110101000001100111001101111101100001110101110010010111101001001101000010101111110011111000101110000100101110001000110101001001000111110101010101101100100111011100100010111111011001000;
#1 $display("%b", po);
# 1  pi=207'b101000001100111000110100111101011011100000000110101010010110101101111110000111101000011001100110000110110011000111010011000101101111100010010111001110001000101000001000010011101010100100101111011000011101000;
#1 $display("%b", po);
# 1  pi=207'b111100111000011110011111101011001111011101111000111001001001100100100010111001001010010100010101000011101011000111101101010001000001011011011110000010000011110110101101100111110001010110110111100000011110101;
#1 $display("%b", po);
# 1  pi=207'b000010011100010110101011111100010100010001011010110111111010001101000010001000011001000011101111001110000010001111101001110101111001010111110001000111011000100001110100011101011110001001111000000011111011010;
#1 $display("%b", po);
# 1  pi=207'b110010101010011101100100001011000011111110100111000111111100011111101011001101001011011001000011101100000101110011011011001001110010100100110100110000010001101010000001001000110110110011011010001110101111000;
#1 $display("%b", po);
# 1  pi=207'b011010010101011100000001100011110011000010010110101011101001011110100011001100010010101101010110000001100101000101000000001010010110100001010011110110010101111101110010100110110111101010000111110001101110110;
#1 $display("%b", po);
# 1  pi=207'b110101001011001001100010011101110110011010100010000000000111101001101101010010001001010100111111110000010011111101111010110110010111100010000011000100010111010000101101010100110101000101110111111011100001101;
#1 $display("%b", po);
# 1  pi=207'b010101011010110011010001010011110000010110100000101010000110000101100011001000110010100100001101000101000110111111011011100011101100100110100100010000101110000111000001111111100101010010111000010111010111001;
#1 $display("%b", po);
# 1  pi=207'b011110011000010101110001101111100010001000110100110001111100010110101111011111001001110011011101100010010100011111110010000010111100100001101001110110010111100011101001100000011001101001011101110101110000001;
#1 $display("%b", po);
# 1  pi=207'b100011011010000100110111001111011001011001011010110000100110011010110100011010100011110001001011000010010101000000101001110011110010001011111000110111011101010011100011000100010001001010011100010110000010110;
#1 $display("%b", po);
# 1  pi=207'b000000011110111011111010010000110011011010111111110001100101010111010001111010001100100001110111010000100101011101110111101111011111111111100101110011011100010101110101111101010010101000000010100011011001000;
#1 $display("%b", po);
# 1  pi=207'b010100101010101001010010110110010001001101100110111001010111110110101101101111001101101110101011010001110110100011100111100000010100111011010101101101110100111011010101001100010001111001001100001100011101111;
#1 $display("%b", po);
# 1  pi=207'b010010001001101100001001100101110001101011010001101000100101010101001100000011001100011110101111100010111010111100100101100110100110100111001110010001001000111011011101110100101001101111100010000111100111110;
#1 $display("%b", po);
# 1  pi=207'b100010101101100001000110110110111010111000111011110000101100000011111101000010011110011100010101000100110100110011000010001000101000101100010100011011000100111110010011101000111110111000110111011011010011010;
#1 $display("%b", po);
# 1  pi=207'b101011000001000010000110110111011000000100111100011000010001101010111011011111110100101001101110110000000110110110100110011010100100110110011111010100010011010010001001010110100000110011110000100111001101011;
#1 $display("%b", po);
# 1  pi=207'b011000111000010101001011111101111011010101011010001000111110111111001110101111111010010110100110111001010110111100011111001001100011000010000110101110101001001000110110010100101111100010001000000110110100001;
#1 $display("%b", po);
# 1  pi=207'b000000100100000000111111001011111000100110000010110011110111100010111011000111011101000000010110001111000110110110001110101100110011100111011100101111111111001101111001110110110001101001000001110110110000011;
#1 $display("%b", po);
# 1  pi=207'b100000101100111000001111010101001000110110101111001100001000110110110001010011000101011001100100011001111100101110100000000110101011100011101100000011111011110101111011101100011001010001011011110000000011011;
#1 $display("%b", po);
# 1  pi=207'b010111001001010001110111100000110110101010110100110110100010110100011011001000110001101001000100000111110011001110000100100110001000010000101110001111100011100110000001111011101110111001011000000101001100011;
#1 $display("%b", po);
# 1  pi=207'b000101100001101100011000011111001101000000100010101111110101010001100011101000101111001001100000001110000000011000001011010010101100111101001000010100000110101001101011001111100000100110001101111001101000101;
#1 $display("%b", po);
# 1  pi=207'b100001110011000100000000001011000100100000000011110000111101011101100100001001001011000010010111110001101101001000100001100010101011011001101010001100111100000111000010110010010100011111110001000101101111010;
#1 $display("%b", po);
# 1  pi=207'b000101101101111011010010011011100011101110000010010111000110111110011001011001000101010100111001110001011000100101001100111001100110011101011000010010100010001100011000010010010101001101110000001110010100110;
#1 $display("%b", po);
# 1  pi=207'b100110100001010010010111101011000001110010100010101010100111111010011101001111010010111111100100100101110010111110011110011111001001111111100110000111111110011010100000011000111000111010101010100110010101000;
#1 $display("%b", po);
# 1  pi=207'b010000111110111001111101111111101101110100100110110101011101011110100100101111100000000110001111010111111100000110010101110000110010111101111110101110101111100101001101100010011011001111101100010111000010110;
#1 $display("%b", po);
# 1  pi=207'b100111010110101111010111100011100001110010111100010111011101110100011000100010011100111100100111110111100011111000000111011111010001101100100001100100101100010010001111111000010010000111101111110100001010101;
#1 $display("%b", po);
# 1  pi=207'b101001001100100100111011010101001001011100100100111011000101111010100010110111010100111001010110011000100101001010100010010000011111010111011100100100001011010110001101101001011010001001100101000110010101100;
#1 $display("%b", po);
# 1  pi=207'b101110110001011010001010000000110011010110111111011111111011100010011110001110000000000101111110101111011000010100001111010010100111010100101110101110110100101011101100100100000100110010101000101101111000001;
#1 $display("%b", po);
# 1  pi=207'b111110100010000100001011101010011111101000110111010010110001000011111101111110110111101111101011000010010001101111111100000001110001010101001100000100101010001111001001001001001111010110111011000000011001010;
#1 $display("%b", po);
# 1  pi=207'b100001111110101100011000110010111010111101011100100110111011010001101110110000111100001110011001100010100100000001001010110000010100100101100011110101110011011111100110110001011100110101100010101110011010111;
#1 $display("%b", po);
# 1  pi=207'b010110111101000010110011100001000010111001010011101001000010010000001100100100101011101101010110000010001100011111011101010001010001000011101011011001111010000010011000011001100110001100110010100001111010001;
#1 $display("%b", po);
# 1  pi=207'b001101110100010000001001110010011001100110111010101010100101110110001001011011000111110001011111001101111010010000011110100001100001010001011100101011110010100010111110101001010101010100100000001010111011101;
#1 $display("%b", po);
# 1  pi=207'b001000000000000100010110000110110100001000001001111011010111000110011100101001001000010001111010111111101001010001010101001011101001101101011110000111101000101001111111110100110110001011111100010000111100100;
#1 $display("%b", po);
# 1  pi=207'b111100011100011100100000101110001100100110001010000001101101110000110001101011011010001100001010111111000100100010010100000001101101100101100100000011110010011100010100010011011111100100001110101100000110010;
#1 $display("%b", po);
# 1  pi=207'b010010111111110111101010101000010001010010101011010010010100000101101011011110100000001100111110000000100101111011111000101001001111110001101010111000100101010110100110010001111110110101001111011110001001101;
#1 $display("%b", po);
# 1  pi=207'b101100011010001101001011011000010100000000011010101010001000011100011011100001110010000111010101010110111001000101110110010001100110001010010011101110110111110101100110101011001101100010011101011000001111101;
#1 $display("%b", po);
# 1  pi=207'b011110000001110000000011100011101011000111001100000000000000111011111000000001010100001101000001110010000100111001101111100100000011110111111000101101101001100000001100011010000001011001001100011101000010011;
#1 $display("%b", po);
# 1  pi=207'b101111011110010100001010111100110110001011011110010001101100010101110001101011111110010100011011011011001001011011100110110111111101111001010100011011011001101010100100001100010111100000100010101110001110000;
#1 $display("%b", po);
# 1  pi=207'b010110001101101111010010111100101010010101011100100111010110010101000101100001010101010010110000111101110000001110100000101101010111110000010100011001000111010001101000111100101100000111101111010001100010010;
#1 $display("%b", po);
# 1  pi=207'b100000010000111010011000101100110011010010000011000110001001011111110001110000000110111111001101010001100100101011001111000010100101011101001101001011010111110100100111100011100001001111001101101001001000001;
#1 $display("%b", po);
# 1  pi=207'b010101010111001010101011110010011011011011011101101110010000000111001000101100000110000000101110010000100110010001001001000001010100010100111001110000111111011001001100110001001010010110010111011100111011001;
#1 $display("%b", po);
# 1  pi=207'b110011000110001100101010000011111000101101010100101011101000011111101011101100110110000011011100100001111000001000110100001101011100000001001100111111101001011000110110011001000010010110100100011101001000010;
#1 $display("%b", po);
# 1  pi=207'b100011100010001110011101101100011111110010000001110111001001010101101110011100010110000010110011110111110111100010000011010010011001000100011100000101010001010101111111110110101000011000101100000011110110111;
#1 $display("%b", po);
# 1  pi=207'b000110100110100110100001111111001011010000111101010101101111101010110100010001011010001011111000101110100101010000110101001000111010100011011000111111100110000111100000111001001110011001010000001111010111110;
#1 $display("%b", po);
# 1  pi=207'b011100111001011000110000100100000011001110000010000001010011111011011000000101100010011001011110011000011010111011011000101111010010011110000100001100011101111101101111010011001001001000110001111101100110000;
#1 $display("%b", po);
# 1  pi=207'b001110100110001101100010011010000100001101011001101011110010100110011011010110011000110100101110110010000100001001101110101000000100011010010001110000101110101110101011011110011111010010011011011000011011001;
#1 $display("%b", po);
# 1  pi=207'b011010011110000100001111011001010001111000011000101010011001010011011101010000010000100101110100111001010010000110100001000010011011111000000111000010011001110111110010101101001100110111000111000111100001111;
#1 $display("%b", po);
# 1  pi=207'b110100100101001101100000100110000111111011111111011100001011111011111011001111101100110010100100011101101001001000100010010100011010100001000101101001001010100110001110001000011001100100010101100110000100101;
#1 $display("%b", po);
# 1  pi=207'b100010100101101010110111100001110100111011111000110000100001010100000101000011110101110000100100101111001100010110011111100001111110010110001010010011000011101010110110001110110000010011110101100000101001010;
#1 $display("%b", po);
# 1  pi=207'b001101100101011000011111110100111010101101001000101110111101001101010011000000010010010101000110011111111110011110000000100111001100000011100011100011101110110101001111001100111110110001101010001110111100100;
#1 $display("%b", po);
# 1  pi=207'b010101000000001001100011110110001011000110110010101101001000111001011101000110011001100110001101100011000000100111011110100100001000101011011111010011101101011011100001001001101000011101111100010111010011111;
#1 $display("%b", po);
# 1  pi=207'b000100011011010100001011110101111001010100111000000010000111011110101110100100100101001010011011110111111110111111111001010000000110010010101000100011011110001011110101011011011011011000111101001101011101000;
#1 $display("%b", po);
# 1  pi=207'b001001001100010111110110111111110110001100101000100110100000100011001100011010011001000110010100000110100001001110000110101110001001100101000001011000111100010110111100000100010011011101001111000101101001100;
#1 $display("%b", po);
# 1  pi=207'b111100101110101000010111011000101010000010001100011111110001101011000001110101101100010011010011010000100000100110101100001011011001100100010111000101110110100101001100001100000100110001111010111100001011010;
#1 $display("%b", po);
# 1  pi=207'b000100110111110110111011100011001111001110101100000010111011100011101010001111111111000001010101010001101111010111101010111001111000101110010011110000100000110110101001100001010000110011000011010100110100110;
#1 $display("%b", po);
# 1  pi=207'b100010010011010111110110111100111000111001111101111001011000000101000100111100111110100011110001101001101000011001011111001001000000010110100101011100001010100100110000111111110110011100000111100101010101011;
#1 $display("%b", po);
# 1  pi=207'b001111010010011100100010110110010000000110010101011100011110100010110000011001110010100011001110110100110110111101111000011010011110001010110111010000110010101101000101011101101001100101111111001011000001100;
#1 $display("%b", po);
# 1  pi=207'b001101011010001100010100110000100111011000000101011000000010100011010101110011100000000011111111000011001001010001000100011110110011100101001010101000101111110110011011010101100010100010010011011100010100110;
#1 $display("%b", po);
# 1  pi=207'b100001011100001011010110011000101011111111010100101010010101100101000010000111100000010010101101001101110001001100101100001000111111001000100100100111001011110110000110100000111110000001000110010111100011111;
#1 $display("%b", po);
# 1  pi=207'b000100110000101011110010100100110010100100110011001110010110011001101010001011100110010000010100000100000000011000101010010011000110000111011001101000100110010001001011101000010100101001000110101100110010111;
#1 $display("%b", po);
# 1  pi=207'b101100110101010110010111110111000101110011011010111101100010101110101000000100010011011101100110101111111000110011101011000000011010001100011101000011001101101000100010111010001111110001110000010101001111111;
#1 $display("%b", po);
# 1  pi=207'b010001011001110001011001100000110011101101011001111001100010011111100110010011010000111010010101111000010000000000000100100010000111101011110111000000001011011011011011100001101000000101010010111000110001011;
#1 $display("%b", po);
# 1  pi=207'b111111011000110100010000111001001010101110001001101101111010010101001001001100110111101010010111101111010010111011001010101110010100110011110001100011110000111001010101000110000000111101010101011001000111110;
#1 $display("%b", po);
# 1  pi=207'b011111110000000110111010010110000110011101000101000100011000110111100101110011100010000110101100110011110101011101100010011100010001111100001100100110011001100101101111010111100101111110100001110101000111110;
#1 $display("%b", po);
# 1  pi=207'b110101100001010111101011011011010110111111101011101001000010100100111011010010100111001000011000001111100010110010000011011100001010110000100111110111010001110110001011011100100001111101101111100111010011111;
#1 $display("%b", po);
# 1  pi=207'b010101001110111010011010000011100101010000010010011100000010001100000101001101011011101100101011000011000111101010101100100001101010010100101000110110011000000000100000010110010001100011111001100011111001101;
#1 $display("%b", po);
# 1  pi=207'b011101000011100000001000000000100100011010011101000010000011011010011110001011110110001001101001100010101100011001100111101000011010010111101101110010011010011101010010111000001010001101001101001110001100111;
#1 $display("%b", po);
# 1  pi=207'b110010001101110111000000000111110010100100011011010011110111001010101001010100100010001000101000001111101001100111110110110011001011000100001100000110001110100010100100111010000100001000110010101010011000110;
#1 $display("%b", po);
# 1  pi=207'b101111001000110011000000010010111101001111111100011111111110101001101010010100100010100101001111111010100110111001000001010100110001010100100101111100111001100001110011001101111011001000011101011111000000011;
#1 $display("%b", po);
# 1  pi=207'b110110010010101000000010000011011001010111100011001111101010010011000110111001101001000101011001100011001010001101111100101000011101010010100010000001011110101101010000110000011110110100111100000001001100001;
#1 $display("%b", po);
# 1  pi=207'b100000001110001000000111111000110111101001101110010100101011010111100000110100111000111100000000100010010001110110001010011100011011101110001101111101111010011000011001011001001101110101010111001011110111110;
#1 $display("%b", po);
# 1  pi=207'b001001001110111001101001100101111111010000111010110100100011011110100100110101000111111011111101000101000011111001110011011100100000000110000011100000110110110010101111000011010111111000000011101111001100011;
#1 $display("%b", po);
# 1  pi=207'b000001000110001000101100010001001000100001101110011110011010011110001110100000001010010100100100111111111011110101011100011000000011000101111111000010010011001111001001011110111100010111110000101000011000111;
#1 $display("%b", po);
# 1  pi=207'b101101111101111011001001101100111110010000000111010010010010000110010110011101000101011000011010011110001111100011001001101000000111001010011011100010010110111011010101000000101100111000110000100010110010011;
#1 $display("%b", po);
# 1  pi=207'b110111011100110000111101010011001111111110011111010000011011011011011000110111100010011101011101111000000011000011101111110101001101010101110110111010111111000100101011000010111100000001010000100110011110000;
#1 $display("%b", po);
# 1  pi=207'b101111110011110000111010100101110011111111011011111011010011011101000101010000010000000000000110110111000011011000111000111001001100100101001010101010111010101000011000100011101110001110101000110100100110001;
#1 $display("%b", po);
# 1  pi=207'b100110100011110100011001000110100000111001110111011101011011110010011010010110110011111001100000011111011110010000100100101110001100001100100011010000111010110000011001010010010100101110000110000111011100000;
#1 $display("%b", po);
# 1  pi=207'b101001100011010110011110100110011111111001011000001101010101010010011111101111110010101101010011100000011101001011111001110100110011000011010000110010110001010110100001101000101111011000011001011011010001110;
#1 $display("%b", po);
# 1  pi=207'b000011010011100110110010010011101011010011011100111100011101101010110110001110111100010100000011100010100011111100010011110110001001010110111100101101011110110111110011001100100100011001101010010000100100110;
#1 $display("%b", po);
# 1  pi=207'b100011100110010000110101100110011111111011000101101111000111010100110111100101010000111101101110111110001010110110011000011010111110111111000011111110100011111000100000100011111011000111110000100010110100110;
#1 $display("%b", po);
# 1  pi=207'b111100000001000101111111010000101011100010000101000100100000100011001101110001100001101100011001001011011000111010011001100111011110000110010100100000111101110001100101101100001011000111110101100011110100111;
#1 $display("%b", po);
# 1  pi=207'b110100101101100000000000011111111001010100110010100100100011100001111111101001110011010101101001101101110100110000110101101101010010011101001000110110001000101011110101010010100101100010111110101100011101111;
#1 $display("%b", po);
# 1  pi=207'b011010101011100111000100110001000000010010001101000010110001011001011011111101010001101110011111100000111101101000000001101010011001001001100100001111110010100101000100111101000101100011001110000101011011100;
#1 $display("%b", po);
# 1  pi=207'b011001111010010010101010110011101101001000010001111011100011001000010000001111111110110101000001111010011011110110100011011000000100110110110101000001001011100011010110010011010111011011001010011010010110001;
#1 $display("%b", po);
# 1  pi=207'b011000101011100110110101111000100011101011000000010010100101001110111000000100100010001001000010101101100011111001010011111110011010110100110101000101001010001010000010000100000111110000111100011001111010011;
#1 $display("%b", po);
# 1  pi=207'b001110100100000100000000011011010010100000100111001110111000010000010000101110011111100001111001001010001001101000010000111110100111011100110110000010111011101100101100011000101101101100010011001010001010100;
#1 $display("%b", po);
# 1  pi=207'b000110111100100101011001010011001010011011001101111001001101101110010111111111101110011110010100100010010010110001000111101001000110000101100100011001110101010010100110111011100110100011110000011110100001011;
#1 $display("%b", po);
# 1  pi=207'b101101001110111101001010101000010000010100001010110001100111101111100110001111011100010111001011001111110001010111111000100110100001100111101110010101111101111010110111000001110110110100101100100000000001110;
#1 $display("%b", po);
# 1  pi=207'b111000110111000011100011010011101101101110000110100111100100111011011000000100110000110011010010111010111000010001101111101101100010110110010101001110101001100001110111011000100100110111011011010100100010011;
#1 $display("%b", po);
# 1  pi=207'b000001100110100001010100010101101010110011101000100010010010010100011111101110110100001100101101111001001000100101101100111001100111010101101101000010110111110110111111010000100000101101100011111001111000001;
#1 $display("%b", po);
# 1  pi=207'b100110001011010111010100001001001100011110110111010000111110011100110000101000000100010011011101000000111101000111100100011010000011010001101011101110001111111111001110101000010111001011111101001011101010101;
#1 $display("%b", po);
# 1  pi=207'b000000101101000111100011110101000100111011101101000011010111011010010010000101011000111111001000000101011001101001010010110111010000110100011010110000011100000110101111101000010000010001100001011110010001001;
#1 $display("%b", po);
# 1  pi=207'b000111101010011000000100001010001111010000011000111001101110110100110001111111000000101110000001111110110101111101011000001011001010011001010110010010011010000111011100001110100011010101001001110110100100100;
#1 $display("%b", po);
# 1  pi=207'b010000111101000010011100110011111000101110110010110110111010000111001100000111000010011101110110111010100111010010101111010000010011100101110110011100101111011011100111101000101000000111001001111001110000100;
#1 $display("%b", po);
# 1  pi=207'b110000001010111010000000110001101001111011101010111101000100111101101100100101100011000100111011000000011011100100101000011011111000101010001111111111110111001000010011001110011011010001011101011011010100010;
#1 $display("%b", po);
# 1  pi=207'b110010011010010011110110010111011010011101001111000010010001001000011101001100011110101110000100100101010110111111001110111000111111001101110001011000011010011010010110110111101110110110011111101110010001000;
#1 $display("%b", po);
# 1  pi=207'b111000011011110110000100101010011010000000001100111001100101000001101010001101111111011001010110101010001011010110000000110011110111010000011100111011100101011001000101100011101100011101000110010101000100111;
#1 $display("%b", po);
# 1  pi=207'b000001111101111111011000111001001111101001010010010001010100001011011001101001001000100101011001110001111101100011110101010111001111000001100011011011011010001111111001111101010001011110101010100010010010001;
#1 $display("%b", po);
# 1  pi=207'b110101010001100010101101000000101110111100010001010101001010011001010011111000010111101110011100110000110001011011100100011111011010101001011111100001000100001100111101001010101100010010110110010010010011000;
#1 $display("%b", po);
# 1  pi=207'b011100101111001100010010100010110100011101110101110100101111101110101100011001101010100111101010101001100111011011001001000010101111100110100100001001100110011000110010010001010100001011010011010010111011110;
#1 $display("%b", po);
# 1  pi=207'b001100001010100011001001100100100101010011001011000011111111000011010100111010111010000011100100111101011110110110110001110000000010111111101101110010000010111100010011001100011101110000000101101011010010011;
#1 $display("%b", po);
# 1  pi=207'b010001010111110000000010011110101001100110010011101000110001010001101001100111001001110101011000001001111100001110001101100010001100111110111011101011111001011010100001111100101011100110010000100111000011001;
#1 $display("%b", po);
# 1  pi=207'b011101010101000101000100000100011110000110100110110010100110100111010000100110000000110110011011110000011011000100111111011100011111110000001100111001101011010010100110111011010100001010010010001010101100100;
#1 $display("%b", po);
# 1  pi=207'b000010110011011111001110111011111100100011001101110110111110001000000010011100111000100100011001001100111110001011111101100100001101011110000000100111110001111010100111110110101010111110100101101100001011010;
#1 $display("%b", po);
# 1  pi=207'b100011100001001111000010010100111101000001000111101100000110100000110001010100110101010111100001010111101111110001101001000001000101001100101010111101001111010011101011000010000100110001100001101100000011011;
#1 $display("%b", po);
# 1  pi=207'b111110111110010101010110010110101001100100001110000001111111111110001000011100000100001100010110001011101000001111001110111110010010110101111110110110011011000100100011000011101001110010011011111001101101011;
#1 $display("%b", po);
# 1  pi=207'b110111000100010111100101100000011101111111010110001100001000101010001111110010111100111000111000101011100111001000011110011100110011011111101000100100100101010010001010100110100000110101000001100110100101010;
#1 $display("%b", po);
# 1  pi=207'b100011000001110011000101101111011100001010111110001101000110010011001101101100001010110110000001100111000101000100110110000011101000111110101101001001100101110001111100000001011010000001000111010010000100110;
#1 $display("%b", po);
# 1  pi=207'b010100101000000101110000111111001000001000111000100010011010110110000000101101000000011100101100110101110000110101111000111010100011010011000110000110010011010010111110101010101101011010100101001011001010110;
#1 $display("%b", po);
# 1  pi=207'b110101011000111101100111101001011110000101000101011110010001101000011001010110000000011000110001010101110100100001111110000110100010100010010001011000010001110111010001111111000111110010100010101001110100101;
#1 $display("%b", po);
# 1  pi=207'b000001001110000000110001011010010100010000110110110001101000001001111101011010010011101010101110001111111011111000111111101010010001011101001101111000011110000010010011001100110001001101100000111000100101010;
#1 $display("%b", po);
# 1  pi=207'b101110011110001000111011101001000110011000000000000000110010100001011100110011010000010000101000010101100110001100000001110111011000000110011010110101010110110001101111100001111010000011011111010101000111000;
#1 $display("%b", po);
# 1  pi=207'b100101010110001010110111111010101110010010001100101011101110011010110010001001110000001000101111110001111101110110111110110000010101110011011111000001010010111101101100011000111100101110001001010010101111001;
#1 $display("%b", po);
# 1  pi=207'b101101001111011001100110111001000111000100000000001101010111100111001100011011000101010001110010010110110110110110001011001000111101000001001111101000110100010000100110101001110110010000001111110001010110001;
#1 $display("%b", po);
# 1  pi=207'b010111110111010100101001011101110110110100110101100001000011011010000101000011000001101001011011101111011111111110110011000111010110001111011011100010110110011010001110111100000010000101001111100000111011011;
#1 $display("%b", po);
# 1  pi=207'b010010101001111011111010110010101001101100110110110111110010011100000100101001100000100010111000110100110111100011000010001011000001001100101101000110111000101000101100100110010100000010101111011001110000110;
#1 $display("%b", po);
# 1  pi=207'b111100110001100101100100010011110000000001110000100111011000000000001011001001010111110011101100010111010111000011100110001111011010010000010000001011000000101001100101110010100010101000010010011000011001100;
#1 $display("%b", po);
# 1  pi=207'b011111110100001011010000101100101111100011011110111101000111100011111100010110100001110101000011101010011110110011001010101000110101101110111001011111110110001101000110010110011000111000110011101110000000101;
#1 $display("%b", po);
# 1  pi=207'b000100100111101001001010110111101010110001000100010010001001010001001110001111011010111110000000011101111001111010011110110111100101101111101011101000011000101100100111001000101101000011100101110011100010101;
#1 $display("%b", po);
# 1  pi=207'b011110101010011101011100011011111111011011000100011010011100101110101111101001011110100000001011100011110111110100100110101100110101110100100110011000010010001001111111000011101100110100111010101101000111010;
#1 $display("%b", po);
# 1  pi=207'b111100001001010011111001111000001101111111001001011010001011101100001011010101011101101110011001111101000011101001110010100100101111000100001100111110101110000110001110111110111111111010100110100101111100101;
#1 $display("%b", po);
# 1  pi=207'b000110001011000010111001100111001011101111100111110000011110011100010100111010111110101001111001011110000011000000000111101111000000110110010011100011100100111001001110100101010110111001001111110011000110100;
#1 $display("%b", po);
# 1  pi=207'b111110100110000001110101101111010000010100011111101101111001101100000000101101101110000111000000110100111110110101111001100111011110110010010101011000101100001001001110110011100101000000001000110110100111001;
#1 $display("%b", po);
# 1  pi=207'b000110111110001001011001101110101110111111011100111110011001001011100100100101011010000001111001111010001010010111010011101001011110110011101011000110100000111001110100100001010001101011011101100001100000101;
#1 $display("%b", po);
# 1  pi=207'b001000111011011110010010001010011111001000100011001110000110110111001010100011000101000100001100100100100011110110110110101110100011111010101100010011000111111100000001010110000010011001111110010110000101111;
#1 $display("%b", po);
# 1  pi=207'b001110110011000111101110100010110000000100101111101001111011111110101101101111010001000010100100100111101011010111101001010110110001101110111001111101000100110001011000100010100001000100111111100110100100100;
#1 $display("%b", po);
# 1  pi=207'b101000100100010100110111110001001001101001110010100000001100000111111011001010111111110000101111100110111110000111011111101000100011111110101110000001011111001101000110110100011110001110010010001010100000011;
#1 $display("%b", po);
# 1  pi=207'b100101110101011100111010111100001001111110000011001010001101010000011011110101111010010111110111110101101011110101001100011111000110111111100100010101101001000110100010110101000001100101110000111111110011000;
#1 $display("%b", po);
# 1  pi=207'b000001110110100100100011100011000000010110011011001011110110111000010110000101100001010010100011110101001110111001011111011111000101111110110111101010001011010100001101011100011111010100110111100001001110001;
#1 $display("%b", po);
# 1  pi=207'b000100001000110001010001010001110111011000101110000110100001100101000101101101011110110010110110010000100110000010101100110100010011110101011110100010101100001100000011010001010100100111100010111111011100000;
#1 $display("%b", po);
# 1  pi=207'b110100000111011100001100010111101110100011110111110110011111110000001110000000101111111110010100010001111010010110100011011000010101011100101001001111010110000100001101011000010010001111001001011110001110100;
#1 $display("%b", po);
# 1  pi=207'b011110001101100111000001011101010000111111111001001111001100000101010011001001001000011000010110000011000000101011100101101001110100100011001111010111101101110011001000110101011111100010000101000010111011110;
#1 $display("%b", po);
# 1  pi=207'b011010010110010101100100001011000000100111101011010101111100110101110101100111011111100111001011111111100101100010101010100001100111100111111000100110010111110000110101011110011000011011100001000101010111010;
#1 $display("%b", po);
# 1  pi=207'b011110100010010011100011000010000110110101101000000011101001100001001111111000110100000001010100010001110111101011100101011000000010010100111101110000011100100000001111010100110010011101101001110000001110010;
#1 $display("%b", po);
# 1  pi=207'b101101100001000101001000100100011001011001101101001100100011000010110000100000100011100010101111111001111110001011111010011100110011111111111101101010011111110000010100100010000101100110010000010011011011000;
#1 $display("%b", po);
# 1  pi=207'b111110001101111000001011010001010011010010101100000110100010101110110111101100110010010100100111100000101101000111001001000101110101001011101001001101001110111110001111101100011101101110011001110000111110111;
#1 $display("%b", po);
# 1  pi=207'b000001101011011011100011101111000100111000100111000100000010000100100010011110011101100001101110000100101100101000010011110101000100010101100010011001011000100000100111011001101000111101011111100101111100101;
#1 $display("%b", po);
# 1  pi=207'b010010111001000110110100101001111110110011010011101001110011110001011010001101011111000110100101001111110111100101011101101011000011100000001011010111010110110110101001010001000001110101100011111000000010001;
#1 $display("%b", po);
# 1  pi=207'b010000001110100100011110111110011010010111111111010101100110101001001111001111001110100011001100111001101101011001100100000110110010000011000011111010100011010101110111101010110110101100111000100010111000010;
#1 $display("%b", po);
# 1  pi=207'b101100111100100011010000011111011110000110110100100110100000010001110001010000001000001111100010011010000001010100010000000001110000111000100010001010111111011111111010111100111111011111110101111000101011000;
#1 $display("%b", po);
# 1  pi=207'b110110110111101011001011011000100100111000111011111011010111000111000000111110001001110011100101011111011110001101100000110001100111001110001010111010000101110110111001010111101110001011111100011001010111100;
#1 $display("%b", po);
# 1  pi=207'b000000101010000001010001000101110011010010000010011001011101011000011001101110001010110101001100101110110011100101110011100011011011110101101001000001101110011101011001001010101110010101111010111101011110011;
#1 $display("%b", po);
# 1  pi=207'b001001101000011000100001010001100001010001000011111111011101000000001111101011110010110101000000001100000010011011100011001101100011010101000000111111000010100111000110100111101011011010101011100001000001011;
#1 $display("%b", po);
# 1  pi=207'b110001100111100111011011111110110101100100010110001001001010000010000101100110101110010101000011110100101000010100100110000000010110100100101011101011001101010010111101001101000111110110000111101111100000100;
#1 $display("%b", po);
# 1  pi=207'b100110001011110101011101011010000101101100110111101110000000110100100001110101100110001001010000101000001010001001110011001100001111010001000110010110110111000001011010100110100100101001101101010011011001010;
#1 $display("%b", po);
# 1  pi=207'b001001010100110110110100110111000110100111100111100100001110010000010000010100000010101101011011000000010010000110111100101001001010101000100111001110101100111100100110111110000001011000000001001010111100101;
#1 $display("%b", po);
# 1  pi=207'b001000111001010000100010100111111100011101010101100001010101001111011001001101000101011011011001110111110100011001110110101010010111000110111111010110010110101000101010000111011101011100010000111110000111110;
#1 $display("%b", po);
# 1  pi=207'b000011011101011001100000011010110111010110001111111100010000101101110000010111001100101011101010011010110110110001101111101101110010010011010000101111101000110101011001011100000000010000111101010110110110100;
#1 $display("%b", po);
# 1  pi=207'b000001000100010100110000100110100010010011011010110010110101011100001010010010010010111101110111101001100100100110010111000100011001011100011011101010100001010001000000010100000111011100011011111001101111000;
#1 $display("%b", po);
# 1  pi=207'b100000011011001100010110011100011101000110101111110001110001111000001010101011010101111101111010100111100001000110110010111110101111010010100101111100001000001110101011000000010001110000000100111010111011110;
#1 $display("%b", po);
# 1  pi=207'b001101111111111100011001110100010011111010110101011010101110010110110001111101101100000101100010111000011110100111101011110100001010101000001000111010011010111101001010110111011101100111110001011001011100011;
#1 $display("%b", po);
# 1  pi=207'b001101101010111100000100001101100000101000010101100111111010111001001010010011010100001000100000101100010101011110111011011110111101011110101000001111111000101100101010110000010000101001011100001110110010000;
#1 $display("%b", po);
# 1  pi=207'b101110011110100101110111100001001010110101011010010000111100101111011010011100100111001000111111001100100000111010110100110001110110111100101100000010110011011001001110110101000001000110011011001111001101010;
#1 $display("%b", po);
# 1  pi=207'b011110101001000010110010101110101000100100100111101100011110111001001000100101110011110010001110111111011011110010110011110001110000100101010001000111000111001010111110011000111110010111110110010101110101001;
#1 $display("%b", po);
# 1  pi=207'b010101000110110101110110110000011101110111101010010110111001010101011010101100111011101001000110000001010000011011011111011000011101001101100001000011001101001111011111110010101011111001110101110011101100011;
#1 $display("%b", po);
# 1  pi=207'b100000000001101001000010101100001001011000110111100111110011001011110010101110110101100011001001101101010100110010111000000110001011100101011010000010010000010101010001111100000011101001110011010011111110011;
#1 $display("%b", po);
# 1  pi=207'b001011001010000010000110010100011100001010100000101010000110001110101101000111111000100001000000110011010111110100101101101011001111101100011001011010101110010110000000011001101100011000111110000011000010110;
#1 $display("%b", po);
# 1  pi=207'b111010011100000010010101010101110001110010110001101000011111011010010111110010111110011101111000010010001100110111001101110000000111100111111000101101110011010100111010101011000101000100011011100110011011101;
#1 $display("%b", po);
# 1  pi=207'b000111001110001111011000100011110010000000001111110110011001111111110111000011000110001001110010010101101000111110101010101001111100110011000011001011001010001110000010100101101100010110001111111101000111000;
#1 $display("%b", po);
# 1  pi=207'b110001110010110001001011001111010010010111100101011001010111110101000011011011000111001110111010010100000000111010000000001000001110011011101101000111010001101111001010101001110001100100100110101101110010100;
#1 $display("%b", po);
# 1  pi=207'b101100011111101000000100000110100110110000001110010011010000100110001101100010001110000100100110101101010010001111000001010011010000001101111011110110111100011110000000100010011111000010011010111111011000111;
#1 $display("%b", po);
# 1  pi=207'b100100110000000111110010110001000011011011010001101000010001111010111000011011011000011011111111100001011011111010010100000100100110110001111111010101111001101011011110010101111110110000101111110110001100010;
#1 $display("%b", po);
# 1  pi=207'b100100011100100000010010010110101011111010100010001000010000010101000010000101111010111111011110001010110010100111111101111101100001110100000110000101111011000000000111000000110000000010110011000101000100110;
#1 $display("%b", po);
# 1  pi=207'b111011111011010011010000101011001101000111000111100101100011001001101000011001011100010111011001100011000101000000011101110000010101010000101010111110001101100001111111000011000101010000001001010000111111111;
#1 $display("%b", po);
# 1  pi=207'b100011010000100101010110111000010010011100100010001011001000100100011001101111001010010101010110001111101111001000001101111101001101101100111001011001010011111001010101111010000011100010101001101000010110100;
#1 $display("%b", po);
# 1  pi=207'b101111100010011100011101011101011101010001101000000001101010101100010001110001010011110110000101011000011111101101111011001110101011001001011111000011110001100110110101001011101110110110100101000100101011101;
#1 $display("%b", po);
# 1  pi=207'b110010101010111110101000000100000010101000101010100101101001000001000111110011111100111110010101010101101000111000010011000111000100100111010000000101110100100101111000111011000001101010100001011000010000010;
#1 $display("%b", po);
# 1  pi=207'b100001001110111101101101100000110111110100111011111011011001010010111011010110001111010001110101001010100110111010001011010010100110111101011011100001010010110000110001100011111101101101010011000110000111111;
#1 $display("%b", po);
# 1  pi=207'b110011000010110100000100101110100011001110101110100101101100100010000111011101011000111110011111010010101111010010011001001011000011000000110111111101111100000101100100010011001001101110001000011100110010000;
#1 $display("%b", po);
# 1  pi=207'b110011100001100111011111001100100101000101100010000011101010000110000001011111101001010100100111110111101010011110000100111111010001100011110111100000100100101101011000110110000011110100110100010110110100110;
#1 $display("%b", po);
# 1  pi=207'b100010101110001011100100001010001101001111001010011011001011011110100111101011101100100000110000011110101111010001000001101101111010011001001100011111001100111001101110010100100010100101010011101111110001101;
#1 $display("%b", po);
# 1  pi=207'b011100000010001110000010111011110110110111110111010110111010101101010111101010111110100010101100100001001011101010000011110101010000000101001011010111000000010011101000101010000110000110101001111000010110110;
#1 $display("%b", po);
# 1  pi=207'b000101000001000001101100011110011010100111010110100111110110011101001010111111011110010001101101110001101100011001000011100100001011001111011011011010101000110010001001011011101010001100000010010100101101011;
#1 $display("%b", po);
# 1  pi=207'b111101100001111010101000101101101101010000010001001000011011101101011000010000111011011110101011011100011111001011100010011011101010101011101111010010110101001010101100111100010110111110001111010101010011110;
#1 $display("%b", po);
# 1  pi=207'b111100110111100110001010101001001011010000000111001011100110101000111000110000110110000001011110101011000000010000010001000000011111100110100111110011011001101101000100010111001001100110011110001101101100111;
#1 $display("%b", po);
# 1  pi=207'b100011000110000101111001011010001000001000011111000010111000100111011101001010100111101001010101001111000100001110111011010000000001000110101010000001110000100101001110100100110100110001111101111110011111111;
#1 $display("%b", po);
# 1  pi=207'b011001010010001011001101100011001101000010110001000010011110000010101000101000001110100111010110111000001001000011011101100011111111000111110000011000111100010000111001110101010111010111011111101110101100100;
#1 $display("%b", po);
# 1  pi=207'b101000101011011000111111110110001110101110110001001010111000101101000001010111011110101110100101001010000010011100100000000000011101110101001100101011011010011111000100101110001110000111010001001111100101110;
#1 $display("%b", po);
# 1  pi=207'b010010101111100001000100101010000110010011110100101000100010101010011110100001111010011110000000110111001011001101101101011000111100110010001011001011001011100111110101100001011000011111110000010010100110011;
#1 $display("%b", po);
# 1  pi=207'b010010001101001001011011001001011110000101000011100010111010100011010011101101110100011011001101001010101110100011011010010101000011100111010010110110110011111010101100110011010101001001010110010100100011000;
#1 $display("%b", po);
# 1  pi=207'b110011011100100000100001111011010011101001010110000011111110001010001011101001011100101000100101011100001010011010011000110011100001100110011011000110000000001010101010000101101010001001011111110100100001011;
#1 $display("%b", po);
# 1  pi=207'b000001100001100001101101100011111100000010011111101110110101110010010000010010011011000110010101001011100110110010001001000101010000010011111111110101010111110110010110111010101000110011001011110001110110010;
#1 $display("%b", po);
# 1  pi=207'b100110100011011111111000000000010000001111111101110011101001110001000010101101001011011011111100010110001100011000010111011110111101000011110000000001111111101010001001111010111011001010110011000101001110111;
#1 $display("%b", po);
# 1  pi=207'b000011001010001000110100000100101000000100000100011000011000111011011011001011100001011010111110110110000110100010010001101011010110000111010000101111001001111111110110111111100011011011100100000011110110111;
#1 $display("%b", po);
# 1  pi=207'b111111001100010011100101001110111100110011011101111110101001001000000010010101001101011001001101111001010110100111110101011111001000010001110001101110111110101000010001101001110100101111011110001100111110010;
#1 $display("%b", po);
# 1  pi=207'b111110110110101111001110110101010010110111001100001111000110010101110111110010101010100111010111000011000100010100111111010100100010111100011101111101010001000100110010011000100110110101110000011110111010110;
#1 $display("%b", po);
# 1  pi=207'b111101010110101011001010110010001011010100011100101100000001000000001100101101001000000111000111000011101110101100000111010110011000101110111000010110111110110010110011010101011100010110101010011011010100011;
#1 $display("%b", po);
# 1  pi=207'b110010101011111101100110001010010101111001100111000110101001110000100010101001011001000000111001100001101110101110100100001111100000111101000100100100011110010101011001011001110100110111100000010101101110000;
#1 $display("%b", po);
# 1  pi=207'b100000001011111110001110100100011000110011011000110001010111011101101010001111000000110101000100110000101111000010000101011111100010000101010101010100010000000111110111010110111011101000001110110100100110111;
#1 $display("%b", po);
# 1  pi=207'b111110010101010000100000111110010001010010100111110110110001101111100010111110110111001110111110111010000000100000100100110101111100000011110101011001101100110000101000100110110101001101101100001000010001110;
#1 $display("%b", po);
# 1  pi=207'b110010010000100110101101010011110011100011101010010111011000011110000111100011010001010100100001110010001001010000011100101001110101110101010110100010000011111100101101000010000001000111010100101111001111101;
#1 $display("%b", po);
# 1  pi=207'b110001010111110011100000010000000101111000010000111001000101101100100100001010011011110110101101100001010101100101011000000010111111001001101100011000001101010000000110100001100111010100101110110011101010000;
#1 $display("%b", po);
# 1  pi=207'b111010101010100001011101101101111011111100011010011011100110001001100000110110100101000001111001000010010101000111001110010110000111111010011000101011011011100000001100101000000100101000000000111101110011001;
#1 $display("%b", po);
# 1  pi=207'b001010011100110110101111100101001110010110101110001001011011100101000000101010111101111000100100000001101011011001000110010100100111101111000000000101001110001111010001001100010010010000000000110010000011010;
#1 $display("%b", po);
# 1  pi=207'b110111111101001111010011000000101101110011000110000111001001100101110000000100111101011011000111111110111000111101000110011000101001101000101011010010011001111101000110011110101101111101001010101010011010010;
#1 $display("%b", po);
# 1  pi=207'b001111001111001000000110000100111111111000010011011011111011110011001010000100001010011110100001010001100001000100010111011001000100000101110011011001110100111110100100101001111111010100100011100000111111110;
#1 $display("%b", po);
# 1  pi=207'b001100101101001110110011011111011011011111011010000010011101011000101100101010010011101111100001111111111101111001010111111011011010100111011101110100101010011111010010111000010100111001000000100010100001001;
#1 $display("%b", po);
# 1  pi=207'b101101111111000011000000010101100000100110010001011111110110101110111101001001111101000000100110011101110111101011100110001110100110001000001100010000110010010110101001001010101101111100000010100100011101001;
#1 $display("%b", po);
# 1  pi=207'b110111111100101010101000101100001100111011010001001001001000100101111001110011101010000010000001011101000110101101101000111101101111110110011011010000100010111000001101101011011111101110000010111111111010100;
#1 $display("%b", po);
# 1  pi=207'b110001100111011011010101011010010100001000000011100100011101110000110001010001110000000101001000001110011000001010101010111010001100111100111101001010100010101011101001010010011001010101001110101000001010010;
#1 $display("%b", po);
# 1  pi=207'b010100011000010000001110101101111000100000001011100101111110111010000101111101000010000000100110111011101011101010111101100011001010101001000000000110011000110011100001110100101100001011010100100100100111011;
#1 $display("%b", po);
# 1  pi=207'b110100011101110001010101011110000101110111110101101011001011000010111001101111101011110101111010100001110111111110100011111110111100000010111000101001000100011011010010101000010011010011010011011010111111111;
#1 $display("%b", po);
# 1  pi=207'b000000110110101101100110001111101101011110000000110001000101001011110100111101001011000001110100110010101101000010010001001001101001011100010001111001110110110011110111100001100000101100101001110000010111011;
#1 $display("%b", po);
# 1  pi=207'b011101010110110100010010100001010011100001111111100111011110100110101100101101001111100101010000100100100101101110101110010101010011011011110100111001101000101101001111010101110000011100100010010001011111011;
#1 $display("%b", po);
# 1  pi=207'b100000011010010001011010100001101110111010000100111010000111101010010100110101011010011000111001010100100101100100111100111110111011000100101001000110110011000001011111110111111000000100010010111100011011001;
#1 $display("%b", po);
# 1  pi=207'b101111100100110010100111101111010100000111001101011100110100001000010011100101101101110110101100001110011111110101100101101111000110110111100000110101010011111010010100001000100101010101000010110011011100000;
#1 $display("%b", po);
# 1  pi=207'b100001111100010100111100100100010111000000001100110001011000100001000111101000000110110000100011111001011011100011110000100110111111100101101001011100110001010000101100101110000000001100000110000011001111011;
#1 $display("%b", po);
# 1  pi=207'b110111110100011010101100001101000101110100101100011101010010101011110010111011001000000011011000100011011001010101101101011101101111100111111110110100001000101101110001011101010100100001000100100001000100110;
#1 $display("%b", po);
# 1  pi=207'b011111100100001001100111101101111011110000100000000100011001011111101010110100000110111100110101010101110110110110111111010110000011101111100001001100000100011111001101111110110001111011100110110011001111000;
#1 $display("%b", po);
# 1  pi=207'b011100011010000110011100110111100111001101000001001000001110000001110111111111000001000101100110110000110101111010100010100001111011101101111111110100110100111100111001011011100110110001110110101101001110001;
#1 $display("%b", po);
# 1  pi=207'b000000100110011110010110000001111110101001101000010111101001100011111101000001010011100001001011001001010011011000011010111100100100011101101110110011010001000000000000001111111111010000010010000111111001100;
#1 $display("%b", po);
# 1  pi=207'b000001110010000011000000101111101010010110101011001011100110100011111111011100111000111000011001000100101010111100001011101011000001010101011011100010011111010011011101111100110010010000110000000111001100011;
#1 $display("%b", po);
# 1  pi=207'b001111001011001111010001001010010111011001110111101000010101100010010111001111110000110011000110000100001100010010010101101000100011111110011110111101110111010110110001110010100100111100101111001001010010100;
#1 $display("%b", po);
# 1  pi=207'b001100101101001000100001100101010000001011010100001001010011100011100011001001010110000000100101111010100110100001010010010010010100101001010111000101111001001001100010110000001110110100010110111011110110011;
#1 $display("%b", po);
# 1  pi=207'b000100010101001111101110110100111001000111001101101011001101110100111101111101010011011011010101100010001110000110101100011101100101011000001111110011101110011111000100000011110110010000010001000010001001010;
#1 $display("%b", po);
# 1  pi=207'b111001000110000101010110100110100010011100111011001001101010011011101011010010110011011101000010000000101100001000010101111010001011001000111111110010110000100101011010111010110001110010000011000010110101110;
#1 $display("%b", po);
# 1  pi=207'b101001111111100101111110011011010101100011100111001000111101111000011100000011001011111110111100100011010110001011110100010110001111101000100101011010000010110000100010111010101101101000001100101001101101001;
#1 $display("%b", po);
# 1  pi=207'b101110100101111000001000001100001000011111011000101100010000111100000110100110101110110101100110111001010110110111101010110110010011011110000111111010010000010001011000000001000011010101010101111101110001111;
#1 $display("%b", po);
# 1  pi=207'b001000111001000000010010101000100011001111110110101010110000111011100001001101000101100000110110001010100001101011111101100010001110100010101010100010001101001001001011001111010001011011110100001010110010100;
#1 $display("%b", po);
# 1  pi=207'b011110110110100001100000011100011010110010100000010001101100110111011111000010110100100101011010101111110010100101001011110111000000101011100001100111011110110100010010001110101011111000110101100110111110000;
#1 $display("%b", po);
# 1  pi=207'b011110000001000011111011111001100011000100111011110011010101011001010111010011000110001011110101000100110100111101111101111101111000100111100010000000110000010010000111111011111100110000000110011000000011110;
#1 $display("%b", po);
# 1  pi=207'b011010110111010110100111100000100001110101000110011011000111101011100000010110011101010001110110100100001000111100000110111011111001010000110110111001010101010001001110110110110101100101000100000111111111011;
#1 $display("%b", po);
# 1  pi=207'b100110110101000101100111100111001011010111110010001011001011001110001010000001000101111101001110111111011010011001110001000000100110011101111000101000100100010001010011100100010100100011000101100100101111000;
#1 $display("%b", po);
# 1  pi=207'b111111101010010001111100110111000000100111001101101110111000101111110010111011101100000111000101101011010001110100100010000101010011101000001001011011100111001001000100100101110010010010110100101010000101101;
#1 $display("%b", po);
# 1  pi=207'b000010000000001111101000011010000111100101011000100011010111101011001000111001011110010001010010100000100101110010100101010111101000011001111000000011111011100001011101111000110111101101011000010001101101101;
#1 $display("%b", po);
# 1  pi=207'b000001000100101001111100101010101001100111100010000001010110110001001100000111111100110110011011100110110111110000110101000001000010110001010100000110011001001110101101110100110001011001110100011010011010000;
#1 $display("%b", po);
# 1  pi=207'b110101011110101101111110001000011010100011000000001111111111000001100010111111000110110100111011000111011010111100001011110010100110111010000111001111010101111011010010011101100011000000001101011000100100001;
#1 $display("%b", po);
# 1  pi=207'b111110110111111000001101000000010111011100101110000011010011100111000111101000000111101010000000001101100000101100011111010001100110001011011101100011001000110110101101000101001110100100000001110101011011111;
#1 $display("%b", po);
# 1  pi=207'b110111110110000001101000001110011110111000000000111001111110010101110111100110111110001011110010000110011111001111111010100010000111000011101111100100111000110110100000111100111011101101010100101110100110111;
#1 $display("%b", po);
# 1  pi=207'b100001001101101001001101100000010101101010010101000000000011110010101101100100101110000010010010100011111011000001111011000101001010100000110000111111110100000011000101101011010101000001100010101101111100010;
#1 $display("%b", po);
# 1  pi=207'b011001010011011101100001110111000111101010101001101001010001110000110011010011101001111011110000001011100110111111101001001001000100111010011100111100001000000101000101110011101100000000001000110001111001101;
#1 $display("%b", po);
# 1  pi=207'b010111010001110011111101001110010111111000001101100010111000111111110111011001110100101110001010010110111010011001111010110011111101101111100110011000111111100100101010000100000011000100101000011100101100000;
#1 $display("%b", po);
# 1  pi=207'b000101110011010000101111100101110011111001111001111000011111011101100111010110100111001111110111100111100100110000000010100001100001011000001101110011100011101101111010101011011101001110111100111101110110110;
#1 $display("%b", po);
# 1  pi=207'b101001001001000100010010000000110100010010000111000110111111000010111000000000000100110111111101100110111010100101010000100101111001110101000001111100110011011110101010010110000111000001001110111011010000011;
#1 $display("%b", po);
# 1  pi=207'b011100010000000111100000011110100100000110110000000100010010011010101011001010001000000101110010111111000111000010000010101111000111111011000111001011000110010011100001110111011011101111100011010111100100111;
#1 $display("%b", po);
# 1  pi=207'b100111000010100001000100100101111010001010111011100110000101010010010010000100000011000001111100010000000011000110100000100011000001101011100111011101100001100111110110001100000000101010101010001111111011001;
#1 $display("%b", po);
# 1  pi=207'b001001010010011001110001001011101011001110101001000001001010010100000111101101000010010101001000000101100000100001010011010100010001000001100010000000100111010101111011110001000111000111010101111101001000111;
#1 $display("%b", po);
# 1  pi=207'b000001101111100010111101100111010011110111101100000110000100111000011011011011000111000100010011110101010000001011010101100011110011101100101111111111111010100110101001110010010011110011010101101001110011000;
#1 $display("%b", po);
# 1  pi=207'b001101111100111101010001001101011000001101110000000000101000101100011011101100110100111010010101011100100010011101111111111100100010000010111000101110111111011101101011011100011101100110000001010111001111000;
#1 $display("%b", po);
# 1  pi=207'b110100101010010101000010111100100110010110001100010010011111111001111101101000011001110010101010110111111101111100011010100010011001111000000101100010011001111110010011010000110011011001110010101000010001100;
#1 $display("%b", po);
# 1  pi=207'b000111010000111000101000000110101111110110110101101010000000111101000000010000111001110111001000000101001100011111010101110101111000010101011000101011110010110100110011001011100000001001011011101110000010010;
#1 $display("%b", po);
# 1  pi=207'b100010001100101111001110101011011111011111001111000011100001101011101000011011000100000000001111101110101011001000001010111001101011011100100110011100011011010111110100101100100010100100000011010001010101010;
#1 $display("%b", po);
# 1  pi=207'b000000100100100001011001111000010010000100001111010110011011100001111000001000011101111000011111101100011000100000000010001000011111011010101011000110000111110011001011011001100100110110110011001100100000011;
#1 $display("%b", po);
# 1  pi=207'b110011001000011101101111111011110100110001000100001110100010000101000000100111000000110100111001101100000101011100001010101011110000011111000101001111110110011111011000001000110000110110101100011001000000011;
#1 $display("%b", po);
# 1  pi=207'b101011111011111100111010010011001100001100111001001111011011010000110000011111110101010000110001001010010000101110111001110111010000000100001101111011011100110000000000100101100010111100001011101001110110111;
#1 $display("%b", po);
# 1  pi=207'b011101101100100001100001110110011011000110111000010000110111100000111100000101001011000011100011000111111101100000011111011000011101001010000100001111110100001100011000110111010100101011101010111101010000111;
#1 $display("%b", po);
# 1  pi=207'b110011111010000011111010100010100110101001010000110100010010010101000010000011010010111101001100001001110100001101011010111100000111100101100001010001010110011000011000111100000100001011010111000100100111101;
#1 $display("%b", po);
# 1  pi=207'b100000111010011000111001111101110011100101110111111101101001101010001110011110111010100100100101001100100011001010000101001011011010010110100101100000010001001010011000101100000000101000001001111011010110010;
#1 $display("%b", po);
# 1  pi=207'b100100010001110111111101001001010010010001000101010101110001111100110001110011010100000111011001110101000011100011101101010101100101001111000001101000001111100011101110101101001110011111000110100110011110001;
#1 $display("%b", po);
# 1  pi=207'b000110010111100011101001001111111001101011001101110001110101110110101100110111000100011100100100010010100111000111010110000110110110001010110010000010001100111011101110101001001011011111111010011001010000011;
#1 $display("%b", po);
# 1  pi=207'b101100100111001001101111000000001110011000110000110110011100011011101001010011011110111110111100111010111110101000001010001000000111101001001010100111010101001011011100000101100001000011100000000011001001111;
#1 $display("%b", po);
# 1  pi=207'b001100001100000011001010101101010100011001110000100111100110010101011000111111010110100100110100100000101000010111111010001100101111000110001011111110001011100101011001010101011000110001010101111011010001011;
#1 $display("%b", po);
# 1  pi=207'b101011101000101101110000010100001000111100110000010010000110001010101110001011000001101101011000010101100011000000011100110010011111110011111000111100001101010010111110100011001001100001111010001110001110101;
#1 $display("%b", po);
# 1  pi=207'b111110100111100001110100010100010011011100111110011001010100101000110110101100011001000001100110000101100000100010010011011011110001001111011101110010110101101100010011001110000011101000111111000101010000110;
#1 $display("%b", po);
# 1  pi=207'b011001100111111000111000110110011000100011111001110110111100111110110101110101101011011000000101011000001000000011101111000101000100111100011101100101010100010100010110000110000111100101010010011000101110101;
#1 $display("%b", po);
# 1  pi=207'b110110011001001000001100111010100110100010000010011100001001101110010001000010111111110011000010110001100010000000101101001010110111110101001110111010010010011110011101100101001110001010010011011011010111010;
#1 $display("%b", po);
# 1  pi=207'b001110100011000000000001111100000010111000001111111101001010000101100010001001000000001010110000010101011100001100101111001010111010101000000101011000111001111000010110101101111100101101000010100011101101011;
#1 $display("%b", po);
# 1  pi=207'b111110100111100100010000100001111111000001001100111001100101011011001100101111001110001011100010101000001101001110000111100100000111011101001101100000111110000111001010100100111001110001101100101110111110001;
#1 $display("%b", po);
# 1  pi=207'b110001110100000001111110001100101101000001010001000110100010110001001110011000010000011001101000110111001010011000000111000110110101010011111001000001010001001101000110011000101101101001011000010001010000000;
#1 $display("%b", po);
# 1  pi=207'b110001011000001010011010010101101011011010011110111011111010111100101111100100100111010000010110000000111101111000101101101010100001001000001111110100100100001101100000111111111010000100011000110000101010101;
#1 $display("%b", po);
# 1  pi=207'b100010100001000111000100111100101101111111110110110101101110001001011001010010010110010100011101000001001000100001111000100111011100001110000100100011100111000010010100101100000001101111010100001110110111110;
#1 $display("%b", po);
# 1  pi=207'b111111000011000110111000001101111101111100001111011010011101001110010011101000101001100111001001111010000110010011010010111111110101010011101011001011111010011010011000110101001110101000001000110101011000101;
#1 $display("%b", po);
# 1  pi=207'b101111010101110100001111010000101011101100110000000000011010100110111111101111000010000100000011101001101010011111001111011110111010101000110001011001001100111010001001011101010011100110100110111010000011110;
#1 $display("%b", po);
# 1  pi=207'b001110011001100101111100100001010001010101110110010100011011001000001001101110101011011101110101110100010000110000101011100010001000000011101101001101100110011100000101111111111001001100110100010000011011011;
#1 $display("%b", po);
# 1  pi=207'b000111011000111001111100010101111100000011001000110101011100011001100111011001010110010000111111111001111000001011011111100111110010110110001010001000000011100101100110010001000101000110101000101011101011100;
#1 $display("%b", po);
# 1  pi=207'b001101111111001101001000101001111111000111110010110011010101001000101110010111010010110000010110010100011111000101001101111100101100001000110110010011000001010101011110000011110000111101100010001001001011001;
#1 $display("%b", po);
# 1  pi=207'b000111011100111000001101010100111100000011110011010110100100100010111001100100011110010001010011111110010111000101001010110101000011111101011110101110000100001111110001010111101111010000100010100111000000010;
#1 $display("%b", po);
# 1  pi=207'b000100010010100100000011011101111111110110100011011010011000000011111011011111010010100010111010011100000110011001110010101101110010110101110011000101000110001011000010011000011110100101011011111110000111110;
#1 $display("%b", po);
# 1  pi=207'b110110100000110111100100100011010010100010101011101100111010001001010100111010111011010001101100010010111000011001001010100000000101101001100000100001101011001001011000010001111011111010110111010011000100000;
#1 $display("%b", po);
# 1  pi=207'b101000110000111000100101011111001101000011100100101011100111010101111100001100111011100110101000001101001100111101011011001010011000110111010000111000101001001100100101110111110001110111101111100100110010010;
#1 $display("%b", po);
# 1  pi=207'b101011110000101111011011010101101101101001111000101001100111101100111001110001101100110101100011001110000000011000001111010000101101011011011011100110011001001100111100111001000000000101000100001011001011110;
#1 $display("%b", po);
# 1  pi=207'b010010111001001001010110101000010011110110101111110110110000110110000110001011000101001011000000000010100000001100100010110000111011100101001110000000000111111010101011010110110001010010001000011010001100101;
#1 $display("%b", po);
# 1  pi=207'b011110110010101011010110101011100010011100010001001110101000101101000111010000100101101001101110110111110011111001100000010111111010100111111010001011111110110010000000101011100100000100010001011001000100000;
#1 $display("%b", po);
# 1  pi=207'b101101110101011101110101010111111011010110111010100100111100110101000101010111000101101010011011111001111100011110101111100111111101101010001000000000111110101101101000111010010100001100110100100101110101010;
#1 $display("%b", po);
# 1  pi=207'b011000000101010100010010001010100110000011010111100000111001100101111011001010100111010010100010001110001110011110111110111010000110001000001001000001010000110110100100101111010101000101101111000100000010010;
#1 $display("%b", po);
# 1  pi=207'b000111001000010101101001011001101110110110001001111011111011101011000000000111111110101001011101101100101111001110110000100000101100011111110110101100100101110000011101110010110110001100000011111011111100000;
#1 $display("%b", po);
# 1  pi=207'b000011001010001101010001011010011100000101000000000100110000010100000000101100101100000000000101110010111100011101101111001110100000000111100010000100011010011001100100100110111000001111111110100001100001100;
#1 $display("%b", po);
# 1  pi=207'b100100001111111001000011100000111111110110110000011011011011000111111001101010111100011010011111010001111001100101000010000000100001011111010000011001101100000110100001010001110011111001100000011011111011111;
#1 $display("%b", po);
# 1  pi=207'b100010011101010000110001110110000101111110010001001001100101001110001000001011101011111001010101110010100101100110011011001011010100011010010111011110011110100001011100011110101001101001011011111000100010010;
#1 $display("%b", po);
# 1  pi=207'b000100101101111110111110110101111011100101100010001000000110110000110110010111100010000011110100000101001000000100000111100011000011101110010100010001101011000010011110000100100100010110111100110100101101011;
#1 $display("%b", po);
# 1  pi=207'b010011000011110100011100110000101101010010100110010111011010100101100001111100011001111110110000101000001010101110101110110001011000101111111001000001100100110100100110101000111010110010111011000101110100111;
#1 $display("%b", po);
# 1  pi=207'b101011010000010110001011011000111010101101100010001100011001100001101000011100111001110001100100101101110100010111010110111110110101110110011010100110011000101101101011100110111100100011101100100100110010010;
#1 $display("%b", po);
# 1  pi=207'b111011010010111110001001111111001100010111001011101010001011101111111100101000000110010000010010100001100011011111001101010001001101110101110110011011110000001100101011011000111111110111000000000101111100001;
#1 $display("%b", po);
# 1  pi=207'b001010110100111110111101001001010000111101110000111110101000110100011101110101000111111100010010111100110010010101011101000110010001100000011000011111010010101001000101110110110110010111101111110011111010100;
#1 $display("%b", po);
# 1  pi=207'b111000001100010011110100110010010111111111110010111001110101111010001100000111001101111101011010001011000111001101111011010011011011011100110101011000001001000111011111011000110000011000111100110011110001110;
#1 $display("%b", po);
# 1  pi=207'b101000110011101001111110001101000111100110111111100011001011101001001010010011110101010111101010110001000100010000111110010111111001000101100010010010111011000110101011111001010101100101100001111101100000100;
#1 $display("%b", po);
# 1  pi=207'b001010101111001010101101110101001110100110101110001010011001101010101101001001000001000111010010110110001001111000111111111010010111101001110111000100110100001101010011001111010111110000101001101011001110001;
#1 $display("%b", po);
# 1  pi=207'b001101111101011001101010100101110111111001101001010110101111111001110110100011100010110001101111001100110111010100111111100101111010100101100010111000000101001111010100010100011001010010010010011001101111110;
#1 $display("%b", po);
# 1  pi=207'b011001010100001100110010100011011100101100001001110100111000101000010100111001011011100101001110011011101010010100101011101101011110000101111100001000111111101010000010100110011100101101101111101111001100101;
#1 $display("%b", po);
# 1  pi=207'b101010110111010100100100001100001100110101010000010001001011010011011001010000000111000111111110000000000010110111011011000011000011000100101010011000000110010001110010010111000111011001000110110001110011010;
#1 $display("%b", po);
# 1  pi=207'b010010110010110000010010111101001101110000001010011111001110111110100000000011010100110001111110100111101110110000101010000001111000101111101110101000101100010100101010000010000101001111100111111010010001101;
#1 $display("%b", po);
# 1  pi=207'b110000001010011001100110001001100100010001000110110101011111110101111110111000010001101001000111101011001001011110011110011101100111000010111110110100011101001111011010110000101111101101101100000100010010011;
#1 $display("%b", po);
# 1  pi=207'b010011000110101000000010001010001101101010000100100011100010010000000101111110100000110110111101100011011101001100000100110001111001101000011000011001000011101000100111010111111110000110111101101101011000111;
#1 $display("%b", po);
# 1  pi=207'b111101000101101010101111000111011001111001011110110011011100010100111011111010010010101010000000101111011100100100101000000100001001111000100111111001110100010001110111111101010111010110100011010011101000111;
#1 $display("%b", po);
# 1  pi=207'b101011001010110101110111000001000001101000000001000101010110111010011111101110000011001110010000111010101101010000100111011101001111010000111000010110011011000101110100100111000011101000011010101101110110011;
#1 $display("%b", po);
# 1  pi=207'b100011010100011011101010111011100100010111110111110000101101011110010101010111111101011110001000011110011001100111000000011100011000000011000110011000111101100101101101011110110101000110010011010001001001100;
#1 $display("%b", po);
# 1  pi=207'b101111100111011000000010001000111110000010101011011101100101100000010011001111010111111101010011000101101001101010011010001011000111100011110000110011101011011001100100101001000110110011000111000010010011110;
#1 $display("%b", po);
# 1  pi=207'b101100100101010110010000111000111010001001101110110111001110111100011001101011010110111110000000000001000011111101100000110100011110001101101010001100110111010010100011010010101111000011010011011010010100110;
#1 $display("%b", po);
# 1  pi=207'b010100001011011010010001101011101000110111110000000100000100100010110111101110110110100111011100100000001000100001100111110111100100011100101011000111111010100000011000010001101000100110100011001100111000110;
#1 $display("%b", po);
# 1  pi=207'b000000101000100101000101100000011100100110100010010000110101010000000011111001100001111000110110001101101001011111110111011110101100101000010001001000001010011100111100000101110100101011100011100001111001000;
#1 $display("%b", po);
# 1  pi=207'b001011101111101100000000100011111100010000010011010011111101001000110110110110101001000001100111100101110011111100001001101011011001010000111111100110101111111101000110100011001001000111110111101101110001111;
#1 $display("%b", po);
# 1  pi=207'b111010100000101111010100111111111000111011111010001001111010111000010010101011100001101111101000001001010001110011101010101000011001011011110001010111111111100100010101111011001011101010001100111011100010110;
#1 $display("%b", po);
# 1  pi=207'b010001010000000010011111100110010101100100001001000110111010100101000100111011111000100011101100101110010111000001101110100001111110110000011110100010111011001100010111001101101100010001011111111011001110101;
#1 $display("%b", po);
# 1  pi=207'b011001110000011110001000000010000001101110011000011000010010101010100001110010110101001100100111011101001111011011100001101111100101101100111001101101111101110010001001001000110111000000110001001111110001110;
#1 $display("%b", po);
# 1  pi=207'b100101110001001001000110000010010001000011111100010001110110101001111101100000010000010101101101001111010010110011011001101101101100001010100001100110010110100011001000110000111000101010100000111001110011100;
#1 $display("%b", po);
# 1  pi=207'b101100010111000010111010100010111001110101011001100011010101011111000101101111011101011110000010010000000111110101010010000101101101110011010110100001110011101101110000110000111111001111101011110111010000111;
#1 $display("%b", po);
# 1  pi=207'b111010011110101101001111001001110001101101000000010111000111011101100111010011111100111011110111001011111011000110110011100010010011001011111111001010111001000001011011111011000100011011110010011011000001111;
#1 $display("%b", po);
# 1  pi=207'b010111011001110010110110100010110101111000111000010110110001100101000101111000110010000101111010001000110011111001000011011010001111101110011100110111101100010101010101111000110000001000100010110010100011111;
#1 $display("%b", po);
# 1  pi=207'b100001001010101110001000001000001001111101011010010100110010100110000111101001011101011110001010010000010101111011100100000100001001010000110101101001011000011001010011101001001100010110011010100111110100011;
#1 $display("%b", po);
# 1  pi=207'b111100010101100000010111010011100011110010110100010010010010110000000011011101011101001100111001110101111001000101000001010011101101101101001111100011101100001010001111101011101000100110110100010101100111100;
#1 $display("%b", po);
# 1  pi=207'b001000011001001001111001100101001100010011001001011110011000111010000011010101000011110110111000000011110000110111011001110001010101000111010011001000110100111100010011110110010111100101010010010111001110001;
#1 $display("%b", po);
# 1  pi=207'b011010000110111011011100100110101011111110001100111111110011000110000110000011011111101010100001010010010110111101110110110110000010101001010010111100111101010111010010000000110000011000000111110010111001111;
#1 $display("%b", po);
# 1  pi=207'b110000101100100010010011101101011100111000111110111001011101110101010100110110100001101010011010000101001101010001011111010101110101000011010111010000100101101110110101111010011101001000011011111110111111110;
#1 $display("%b", po);
# 1  pi=207'b111010000100111100010111000101110110100010000101101101101000000110101010100011011111001001010101001010111000111101001011110001100000010010101101000011001111101100000010010100010101010011111100010100011100101;
#1 $display("%b", po);
# 1  pi=207'b010100111001110000000111111110011010101111011010000010110101110110101011110110011001011011111100101010011010101000000010100010010111100001110110101000001000001000001011110111100000000110101000000001011010101;
#1 $display("%b", po);
# 1  pi=207'b111000011001100010101001111110010000000100001111101111000001001110110001100100000100100110101100011010101101010101001101110100001001110111110001000100000100111011110101010000001011101100100000110001101100011;
#1 $display("%b", po);
# 1  pi=207'b111100010000001101111000001110001110011011110100101100111010011101101101000111001100111000000100001001101111000011110010111000011010001100000111101001001111010001101011011100110001110010001110011110000000000;
#1 $display("%b", po);
# 1  pi=207'b110111000100110011111101010100111011110100011100100010111011100001111000001010111101001111110001001001001000111101101010111001010110111100100000001110100001110000000101000101100011001001000010010011010000001;
#1 $display("%b", po);
# 1  pi=207'b101010100100001000111011001100001010010100000010011111011011110010001011000110101110010101011010111111111011100001111000010011101101100001000010001011100001001111010111111010101111010100111001110101011110100;
#1 $display("%b", po);
# 1  pi=207'b010100000001111000101101010001101001110110110011011110001000100101010111000110111010111010111011101011111001010011100000000000001011100100111011110101111100110100100000110000010010001100001000100001111101100;
#1 $display("%b", po);
# 1  pi=207'b101110111000110000000001101111100111000110101010100011001010100111010011100101001100110111011111100011011001001011000100111101010110100011000010001110000010011000100100110011010110001111100011000100110000111;
#1 $display("%b", po);
# 1  pi=207'b011110111111101101001011000111000011101110111011010100011101110001001110001010110000101110100110110011110100000101001100001110111101010100000000100010111101101011100011011011001100111100100010101100100111110;
#1 $display("%b", po);
# 1  pi=207'b111010100111010101010000001011001100010011100101100011101110110011110001110110101011101000000000110110110101111110111000000001101111011000110010010001000110111111010011010011000101000010110101111010001000001;
#1 $display("%b", po);
# 1  pi=207'b110011101001111000100111111001001100101111001111101110111000100100111101110111011101001100011100010001100001110111101010000001111100110001010001010001001101001000011100001101010001110011100101101101000011000;
#1 $display("%b", po);
# 1  pi=207'b000111001000101111111110011101001000001100001101011111101111010000001110101011010100101011000010111100111011110011111011000110100011010110110011001000110101001111110111111010110001111101101001110001010010011;
#1 $display("%b", po);
# 1  pi=207'b111100010110101010101100000011110001100111101101000001101111100111001011110100111101101110111100100010100010001100010110011010111001000001101100011011011100001101011110011101111110100110110110110111111100011;
#1 $display("%b", po);
# 1  pi=207'b001001001000100100000010110110100011101111010000011110101011010000011001111111100101011100000110010100000110011110110011011000011010011000001101010100011101111111111110010111111101001011000000000000101011110;
#1 $display("%b", po);
# 1  pi=207'b100010101101111110011100001000100111000100110010101100101110101001010001011001100011001011000011111100011001011001100111011010011000001010111011101001010110111010100111010010011010101001011000111111001011001;
#1 $display("%b", po);
# 1  pi=207'b101111001010110111001010101001000011011101110011100011010111010110110000110000100101011010011100011111010011101011100010111110110110101111101011111101101010010110000110101111111010110010111111101110010001111;
#1 $display("%b", po);
# 1  pi=207'b000011101000110101001110100000001110011100001010111101100100111110010001110000111010111111100011111001100110000000100100010011011010000011000110010101010100010010011110000011001001001101000000000110100010110;
#1 $display("%b", po);
# 1  pi=207'b101011010011111111000101101111011001111111101101100110100101010001000111001001111001000010110011110010010011100101110100111010110101100001111100100000101001101111100011111100110111001001000110010000010010001;
#1 $display("%b", po);
# 1  pi=207'b001100110110100011110011111110111000001101100001001101110111110111100011000110110000010100010110001110011010110010101111110010110101100111000010001000010111110111110100110010011000101010010110110011000000110;
#1 $display("%b", po);
# 1  pi=207'b100100001110000010110111011000100001000100100010000000000100000111110001100101011000011110110101001111000101101111100010010010111000001011010101011111011001111010010111010101010110111010100110000010111001101;
#1 $display("%b", po);
# 1  pi=207'b010101011000111001111100100101111110001110011110011101100111110100011100101101110010010110011011000001100101110111011010011111101001000110100101010001000000000110100100110110101100100011000101000010101110000;
#1 $display("%b", po);
# 1  pi=207'b101110001111010000001001110100110111010000001010000101110111101000110111101110010000111010010011101000100000100011010100010110010001111010010111000100000011010111010000101111001010101000111100011000101111011;
#1 $display("%b", po);
# 1  pi=207'b001010001100011000111001100010011000011010010110101000000000011001111001001110101000000110100000110000001100101001001100001101100011000001010000100000110011111100011010110100001000000011100101001110101101111;
#1 $display("%b", po);
# 1  pi=207'b000011111111010100000001111000101100100000000100111010101000001110100101101000000011011100010100110111111011101000111100100001010101110010101001000011011000011111000100101110001110101111011000001101110111010;
#1 $display("%b", po);
# 1  pi=207'b111001110110100001000010101010011101100100011000111001101110101101001001001011110100011100000001111111001000010010011001011101100011000100000110110010011110111000101010101111011010000000100000010111110111010;
#1 $display("%b", po);
# 1  pi=207'b111011010011010000010100100010111011101100111111100000011010101101111010111111011100010000100100011101000110000011101011011110101100001111111110110011010111010111010010001000100101110101010000100000000011110;
#1 $display("%b", po);
# 1  pi=207'b100101010001101101010111100110101101110111001001001010101011111110000000000100100001100011101101101110111010010111101000011110110110110110001101000011110110010111000001010101100010110100001100111011010000100;
#1 $display("%b", po);
# 1  pi=207'b011010111011111011011011011110101001011000100101100010010000000100101001001010110101001010100011111111011010101100110101101101000001101101010100011110000101100100100011011100001011000001111100011110110000111;
#1 $display("%b", po);
# 1  pi=207'b001111010001011100101111101101001000101010101111101010010111110100100101110110011100011011101111010010010100101100011010010011001001000110001010001001011011100001011110010011100101111110110011001010000011110;
#1 $display("%b", po);
# 1  pi=207'b111011011100111111011110000000011000000011011101011100011100100111100010000111011111101101111010110001101010110011111000000000100000110011010101100100111001000011100001111110110000010000000111000111101111100;
#1 $display("%b", po);
# 1  pi=207'b000100000100011001001011000111001111100001010010001000010100101000110011000010101010000100001110001110110000100000101011101000111100011011110000101100010000001111100101011100011000010100100001011100110001011;
#1 $display("%b", po);
# 1  pi=207'b010011111011110110011110001010101101101000001001000010111111001001011100001011011010101000000100111010110111100010010001100101110101000000001101100101001011111000101101011101010010011101101011011001010010110;
#1 $display("%b", po);
# 1  pi=207'b111110000010010110100110100110100111101010001001110010010001000101000101010010010110110011011010110001001011101011100101001000111100101010011110111101011111110001111010011111100000001110111011011001010000101;
#1 $display("%b", po);
# 1  pi=207'b111000100000100110011111011110000011101010110000110011100110010010111010001100101001101000001101011101110011111100001100111110111111110000010011001011000010110110001000001000101111111111001010110011110011010;
#1 $display("%b", po);
# 1  pi=207'b000111110101100100101101011000111011101010110001000011110101101011010110011011001111000010101110011010001101001100100110010101100001110010000011010011001100011100111110111101100011110110100001100100011111001;
#1 $display("%b", po);
# 1  pi=207'b100001010010101001011111111110011100111000000101011010110101100011100010010010011010101111010110000110110111011110110000010001010011011001100101100010000110101011111101101111011110011101010000001101101011010;
#1 $display("%b", po);
# 1  pi=207'b000010111111001000100111000101010110011101000011111000011011110111000101111010111101010111100110001010110000001111100011011010111111111011100101000110011000010011101010000100101010001100111101011001111110110;
#1 $display("%b", po);
# 1  pi=207'b101111010001111100110000101011011100001101110010101010001101010110010010001000111100110011101011010101000000011011111000110000000110010010100001011111100100001000100110110110001101101000101110111100000010101;
#1 $display("%b", po);
# 1  pi=207'b000111010010111101011111101011111111100100101101100111011111011100110100100111110001111010110011000101011100110100001001110101110000001110010000101101011100100100101100010000100100001110011100101011000110011;
#1 $display("%b", po);
# 1  pi=207'b001001100100010110111010010100000100101010101100000011110010100000100110110010001001101001000110000111001011010110101011010011010011001000100011000110111010000000000111110100011000101111001010111110100111000;
#1 $display("%b", po);
# 1  pi=207'b100110101110011000011000010010001100000010101011110011100110110101100111000110001111001100110110000011101110111110110111101100110001101010010111001001101000101001010001010001111111010000011011011000001001111;
#1 $display("%b", po);
# 1  pi=207'b100001011100000001000010000100010010100101111101111111110000110101000101110110000010101001111111110010011101011010000010110011000101010010110000111011011111011100001100000001111100100110100110011111010011011;
#1 $display("%b", po);
# 1  pi=207'b010001011100111100001110111001101001101110001000011010010100000101010100001110111001110110001001010000110011111011101100111001011111100110011010101001001001111100110011101011110001000001010010101101011101110;
#1 $display("%b", po);
# 1  pi=207'b000110111000100010001000110100100010000110111000001000101101100001001011011101010100100011111110100011001110101100110011010110011001110011011110101110000001100010011111001100011000111111100110000110100101111;
#1 $display("%b", po);
# 1  pi=207'b100100011000101100001110100111001111000011110101100011100001111101111001000011011010000011110000110101101111110011010101010000110000011111011101100011110111001011111001100110101011001100011100001011100010011;
#1 $display("%b", po);
# 1  pi=207'b111000001000101000101010011010011000101010000111011100011011100010001000001011111101100101101111111000110000000000011100100111010101001100111011111010011110011000001001100110011100010001010000101010001101001;
#1 $display("%b", po);
# 1  pi=207'b101110100100010001000001101011100111101010000111011100101010101111000110011100110100000000111111100101001011001000001100101101110001001100101111011001000011010101001000001111111000100111110110101100111011110;
#1 $display("%b", po);
# 1  pi=207'b001100101011110100000010100001010001000000010100001000110010011111110011101001100100011101100001000101101001000100111010000000011100001100111010101100110101100111010011101100011001000110101000011011011001001;
#1 $display("%b", po);
# 1  pi=207'b111101011000011011000100101010010011101100110010111100110101100001110101001100010011001100110100011111101110110101110010100001000010001111011110110010000001000000001011011000100010101001001110000011101000101;
#1 $display("%b", po);
# 1  pi=207'b010010011101010010001000101100110010100010101001001001100110010111001101000000111000100011001110000111011001111100001000000000000011001011001010110010010101001100101001111010010001101000001010010000110000001;
#1 $display("%b", po);
# 1  pi=207'b010100011001000001000000100101000101010010110011100100000000110101001001100011110101010101101111101101011101011101011101000001001101011111111101101011100000000110100000000000011111011100100001110110111001011;
#1 $display("%b", po);
# 1  pi=207'b110110101110011110110101011011111011011110000110001110111001101110000111100011010101100111000010110101111111111101011000000101001101011110001010110001010000111010011010110010110010011001011101111101111011111;
#1 $display("%b", po);
# 1  pi=207'b101010001110001010111111111111100010000101010101000000100010111111111100110001011001000111111010101100001000000001011011010100100001010100010101011111001001011001111010111101001011011010000110101110101111000;
#1 $display("%b", po);
# 1  pi=207'b011100011011010000010111101111010011000011100011001101000011001110010101101001110110111000000010100111110010111011001100100111011001101010110100001011001011111111110010010111111101101000010011100111000101111;
#1 $display("%b", po);
# 1  pi=207'b000101010100101000010111101011001001101111111000001010101100100100010101100010000101101001100100010110100101010001100011100001110110101011001001000010000000011010011011001001001010010101010001111001000011100;
#1 $display("%b", po);
# 1  pi=207'b011100001011111010101100111000001000110010101011111100111000111001001111111111000011001001100100000100010110001011110110100111111000110011101010111000001011001011011011010111100000010011111101101101111111011;
#1 $display("%b", po);
# 1  pi=207'b111101100110000010111101011101010010010011001101100000110000001000010110001000100010101100011100011010011110011101010010001000001101011001101000100110101101010010110101101010110111011101011010110101001101011;
#1 $display("%b", po);
# 1  pi=207'b011100100011000110010001111110100010110110011110011011110101010011101000101110101001111001101111110110010110100100100100000101010110101001111111010111110111101100010001010001001011111110011000000111110100100;
#1 $display("%b", po);
# 1  pi=207'b001101000101011011000101001011101001100111001110001110011101010100011101001000100010011010000001011111101101110001010010101011000110011100011101010010011001110111011011011101110111000100001010010100001111111;
#1 $display("%b", po);
# 1  pi=207'b110111100100101010001001011110101101011000010100100011111101011011110001001110011010111010101000101010000010011010111010101010011101111011010001010101010111010110101100110000001011111111110101000100001110100;
#1 $display("%b", po);
# 1  pi=207'b101010101101010101000000110110101100111001001110110110100010001111010000111111010010111101100011001000100011111101110111111011010000000110011001100100011110000101011011101000110110000011101100001010110001011;
#1 $display("%b", po);
# 1  pi=207'b001010111000110001010110000110010110100111001001011010101101111111111001100000011101001111001100100011100000011001001001011111100000100100100001011100001000011111001011001110010111000110111001000001110001011;
#1 $display("%b", po);
# 1  pi=207'b010000011001100111011001011101011101001000011010101001100100101001100111000011111110111111001101000110110111110000111010100001010001001011010110100110100100110001010111000011110001110001111001101101000000111;
#1 $display("%b", po);
# 1  pi=207'b011010000100010000010100110101110101111111101011111011110011001100010010110000110110111101010010110010001100100001001111100010100111010011000000011000001001010110111011011100110000001101101000101000000001101;
#1 $display("%b", po);
# 1  pi=207'b001101011100001010111111100101000001011100101000110000000111110111001100010110000001000000001110011101100111010110101101010011001110111111010100111100101000010110101100010001100111001111000100100101100100000;
#1 $display("%b", po);
# 1  pi=207'b101000000100111000010111100000001001111101010110011100111100101100010110111011100011001110110000000100100001001010011000110100101111000001110111110111100110101001100111010101100001010100111110100111001000010;
#1 $display("%b", po);
# 1  pi=207'b010001100011001010110100111110000110011001010110011110011101001111001110110110100000100100011100001100110010001010101011010011001101011001100101101101011110001001010011111110101101000110101101011001001100001;
#1 $display("%b", po);
# 1  pi=207'b000101100111100101000111111001010101011010110111000011110001100100000110001100110011000110000101000111111001111001000111110100101101000011101111100010111011111101001011001010000001000000111111011000001110100;
#1 $display("%b", po);
# 1  pi=207'b010010110001001110010010010010100011011010011100001011010110001011011111101000000010010100100001101000001100100100001011111011011000000010011000001100001010110011010110111111100110101010111000011110111011001;
#1 $display("%b", po);
# 1  pi=207'b001001011001011100101100010000010101111010100111111101111010000111111101110110100111011111111110011000101011100011010010001010110111001101101000110001111010111111000100001100001111111010100101111001000110100;
#1 $display("%b", po);
# 1  pi=207'b011000011100010000000111011000101110110100001010101000001001000001011111100110000101100101100100110010000101000001100000000100010110011101101111010110001010111010111100010000110010010111100001100101001001011;
#1 $display("%b", po);
# 1  pi=207'b101011000110101001001001000001010111100011011011011110001101010100011010100111001110000111100100001001101100001010110101100100011100011010111101001111110000001110110100011011111010011110110111001000010111001;
#1 $display("%b", po);
# 1  pi=207'b100000100000100010110000101100000111010110010001101010010100000000111000111000010010101011011100110101010101000010010111110100101011011111000010101010110010000011010011101001001110110111001010100110000100000;
#1 $display("%b", po);
# 1  pi=207'b101111001010110001011011110111110100001101010001001001010110010001111000111011011111000100100110010011000111011111111101110110001111011110001010001100110000110010111111111101000000010001110011010111101011100;
#1 $display("%b", po);
# 1  pi=207'b001000111110111100000010011110111111101101110110100000001110001111011110100001011100011000100111000101010100100000111011110110100001111000101100101111000111010111111110010110111101100101001010011010101011001;
#1 $display("%b", po);
# 1  pi=207'b010011101010101111101011100101101101000001110011010100011101110010110100001100100010110111101000010011010011010001100000101011110111110001001100110110110111100110110010101000101100000111000110001010001010011;
#1 $display("%b", po);
# 1  pi=207'b001010001000010100010000101011101101010101100011001011111101001101000100010011101111111111000011110000111010110110001101000001010111000101110011110101011100001111100000010011011000110100110111000111010011111;
#1 $display("%b", po);
# 1  pi=207'b111000111010110010110010100000001000101011101101110011001000011111010101010011001011000101011101010011111000010101001010000111001100000011000011100100110000010011000100101101001101110101001000100010111010111;
#1 $display("%b", po);
# 1  pi=207'b000100111100101000000111110000101101101111100010100011110111101011001000000001000100000010000001010110101010001000011101011100000101111101110110110011100100101000100000101111111100111001101001010010111100010;
#1 $display("%b", po);
# 1  pi=207'b010011100101101001000111101011010100001110010010001110000110011000011110111110110011101000011101010001110000001001111111101010001001010000010111100111111001010110100111011000111001001011011111001111110001010;
#1 $display("%b", po);
# 1  pi=207'b001001010101110000111100101010100011010011001110101000000000101011111001110001011110011000111010011011001110000110101100100000001100001110011101000110111010111010101000111001001011101010100111011100010101000;
#1 $display("%b", po);
# 1  pi=207'b111010100001000000101000001111111100000101101110011000000011110111101011110100000010111110111000101001010100001110110101110001001111001110011010110101000101011010010000100111101110001011100111001001111101100;
#1 $display("%b", po);
# 1  pi=207'b000111110000110111000111000110001000000011010100101001010011010000010010101000001001001011001111100110010000001101010011100101100001000100001000010000111100001010010100111001001010010101100011001000100101111;
#1 $display("%b", po);
# 1  pi=207'b101010100000111011000010010110100010001101011100111011110111101101100100000001001111110111010100111000010000010010101011011000101100010000101111011111111000111101111101101010111011101001010111000001101110011;
#1 $display("%b", po);
# 1  pi=207'b111101101100100101110110111101101000000110001100010001001110011001100110011101001110110100110011101011101100010010011101011110110100011010011010000011010101000011001000011100000111011001110100101000110110101;
#1 $display("%b", po);
# 1  pi=207'b000001011010000110111010011011110110000000101010101011100001110101110010001001110111000101011010000110101000110110001110011000100010111010011111000110010001101011110101111111110000100010011001001111100001101;
#1 $display("%b", po);
# 1  pi=207'b011111000101011110001111100001110011001101111100011111101110100010101101001000110100010011000011100111110100001111010001010111110111111000101101110011100001000110110011000011111101101111101001011000110010101;
#1 $display("%b", po);
# 1  pi=207'b000000010011010100101101101111000000000100011010011001001000101001010110101001101010011000000111011001011001101001110101111100101110011111101100100001001110010010110010111111100011000110011000000001111010001;
#1 $display("%b", po);
# 1  pi=207'b000101000000111001110111110000110010000010110111001011010110011110100001010010001101101011111111000011001000110110100010010001111010001011000111100011001010001101100010000101000100000110010101000011001001100;
#1 $display("%b", po);
# 1  pi=207'b110001111011000010100001110011000001010110011111000000010010001100110111101000011110100011001100011010101110111010110000000111110000111000111010010111101101101100010111010100010001000010001100110011011010000;
#1 $display("%b", po);
# 1  pi=207'b001100010111001011011100110001001001010011001010111001011100010100001100001111010101110001100000100011010011011101111101101000001101011000101110010100110111101100110101010010100110010101011000100001010101100;
#1 $display("%b", po);
# 1  pi=207'b101111101110101011011111101010110110010010010100110110111011001011001011011000111000000010011010110001001101100110000110110111000000000011100111101010011010011011010110001110011000111001011011101011001000110;
#1 $display("%b", po);
# 1  pi=207'b010110110011101100010000011011100011101000011111010010111011111110011110011111011000011100010001010100110101101010100111111010100000001111011100000110010110110011000101101110011101011101011110010001000101010;
#1 $display("%b", po);
# 1  pi=207'b100010111010000111111010110101110011110100111010010001000000111000101001100111111111111111110001011011010001010000111101001101111101011000100100000101111011010111110010000000100100110100111111100101011001010;
#1 $display("%b", po);
# 1  pi=207'b001101001111000100010001100001101010100101000101010000110010001010110000010101000101101101011111110010011111111100001010001110111101000011111111000101101100010001100100011000011101011011111101100111010010100;
#1 $display("%b", po);
# 1  pi=207'b001011111001001110000001100011110001011001001110111000000110000011000101001000001010111001011010100010000011100001111000010111101010000011011100000110001010110100101010110110011011011101100011001110110100110;
#1 $display("%b", po);
# 1  pi=207'b101110100000000001101100010110001110111110000100011001010011110011100110011011010110010100001101110011101100011000011100010000101011100111110100000000110010010101001011000000001001100010110000011010101011000;
#1 $display("%b", po);
# 1  pi=207'b100101000101101010111101111010110100010111110111111000011100100100110110010010100001111111000010010011100001001100000100000100010100001011010111100011101001010101111101000100010010110101010101010100000101101;
#1 $display("%b", po);
# 1  pi=207'b110101011110010011011110001111101010100000100101011110000110000110111110010010001010101110111110100100110000010100000111100010100000110101100001110000001100110111010100100101011011101101101100000111010100010;
#1 $display("%b", po);
# 1  pi=207'b101111001001110011100100001000100011100001110110000101100010100110101001000000001101001010101001010000111010000011010100010001001001001110111001011100100111010000000110010001010011001011101110000000001110010;
#1 $display("%b", po);
# 1  pi=207'b010111111011011001011101111110100010011010011001111011010111000010111101110101101001101101101001010000101100111111000000001011101111010110111011111011111000100111110011011000001000010110110100011111011100011;
#1 $display("%b", po);
# 1  pi=207'b001101101000101011011101101001110000000101000111011001000010101000000011011000110111110110010100101101111100111110011010110011011001100010101101100111001011101111101111101111100001010101101000011110001011001;
#1 $display("%b", po);
# 1  pi=207'b101110011011100100101100110100100010101011100011101010101100110001000100101001001110111000111101000101111000101000001000010101110111001000001001100100101011110101111111111011001100111101010101100000110101101;
#1 $display("%b", po);
# 1  pi=207'b001011111101100011001110000100101111001100101100011101000100100110001000111110010011110111110000110111001101100010011110110111010011010100010000101110100010011110110011101001001010010010111011100011001110001;
#1 $display("%b", po);
# 1  pi=207'b010110000011010110011101011010010010001100010011001100100000100100000011011110101000100100100001110010001001001000100010111001100100011101110101000110011010011101001100111011100000110000001011000000000110010;
#1 $display("%b", po);
# 1  pi=207'b011110100000101010011110000001101100100011000000111011101110100100010000111110011000000111011100000110001101001100100101111101111000100001000110001110001000100011000110110010010101100010111000010101110101011;
#1 $display("%b", po);
# 1  pi=207'b110110010110011101110110101101111110001010011001100001011000101011100001011100011111110011110010010000011000001110011011010000101101111010001101000001101000100111111011010100001101000011010011101000100001100;
#1 $display("%b", po);
# 1  pi=207'b011101001110110111101111011000101011011000110110110110000100111001100111011001011000101011001101100110111101110000110011001001110111010000001011111100001101100100010000000000010000010111011000101110001111011;
#1 $display("%b", po);
# 1  pi=207'b110001111111111110010100010101101000000110111011011101100100000101110010100110001101110011100011110101010100010101101010001110101110101110000100010100010101000000010001011110110011111011101101000101011001100;
#1 $display("%b", po);
# 1  pi=207'b111111010101011110101010001010010011101110100011111011010011010100110111001010000010110010001000110110000000001011010010101110001101000111011001000000001010110001111010010001011101101010011000000011101010010;
#1 $display("%b", po);
# 1  pi=207'b011101110001011011000100111110100100100011001000111010110100100000001110110010000111000011011001011111001111100001111101011011111110111000000000011001111111101101100001011011101101101101010101010011101101100;
#1 $display("%b", po);
# 1  pi=207'b101100001010011101000000000000000011010110011000100001010110111111100111011000000110100000011011010101010011111111101001101001111101001100001110111000100100111010001111101110100000010111000001010010010101111;
#1 $display("%b", po);
# 1  pi=207'b011100000111101010000000010011001011001010101100010010001010101001001110010000000111110100001010001001001111010010010011100101100100111111100110010000011110001100101111101111011100100101111011011110100111101;
#1 $display("%b", po);
# 1  pi=207'b101011011111010101001001101101001011010011110110010010000000011000001011001101111100110101011010101010111011011010111001001110001111111110111101001011110110000100000110111110000111111110100000011100110011111;
#1 $display("%b", po);
# 1  pi=207'b110110001111101111100101010011110111110101011000011111011111101110101011100011001110000100000000111101001000010011000101111111110000011101000111111011000111101000000110001111001101001001100100100000100010100;
#1 $display("%b", po);
# 1  pi=207'b010101111011111111001111001100110100101000001011111101011111101111110101110000010000110110000100001000010111001001011100001101111010101101001000100001100100010010100001001000110000010100001000001100001101011;
#1 $display("%b", po);
# 1  pi=207'b111010000000010101111000000110001100111001100101001101010101110010011101001010101011010101010100110000011010100100001001111001011100000001100000001100100011110110100101000100001010001110100000110100100111010;
#1 $display("%b", po);
# 1  pi=207'b000111011001111010000111001011010101011101110011110011001111011000110100010100101110010001011000101001100001011110001000001101111001011001000001111110001111010101101100101001100110101100010101001001011011011;
#1 $display("%b", po);
# 1  pi=207'b011101110001011010110000000111010100111111011001101001110110101000001111101100100000000001010011111000100001110001110111101110101100111010001111111100110111111100101011001110000111010111101010000111100101001;
#1 $display("%b", po);
# 1  pi=207'b110111010101100010001000001100101010011011110111100111110010100001111111111101110000001000010111001010010000011010111000011010100100110010111010000000000110010100010001001001001001001100111010110000110000000;
#1 $display("%b", po);
# 1  pi=207'b010000000000110011111011011111000011001010111110001101111101100001110100010100010000010101010110100111110110000111001111100100110101111100101101101100010111010001100001010110000100001101100000000110000111110;
#1 $display("%b", po);
# 1  pi=207'b100011000100011010000001110001000100011100001111011001100101001100011011101111010101010010101110101100001011111000100011100001110001101010111110001110011010001110111011110111000100010110101010100000110011011;
#1 $display("%b", po);
# 1  pi=207'b100001001010011000011010100011000111011111111100100100110010100000011000011000010100000111100110111110110110111001110101100000100101101000011111000110011101010000111101010001001111001111110100010111010100001;
#1 $display("%b", po);
# 1  pi=207'b011011011111011001000100010010111100010111001000110010010110110101111101001000111100011001111010010010001110010111100011000011100101101010110011101010111010001011011110010011100011111001001000101110110100110;
#1 $display("%b", po);
# 1  pi=207'b101011010010011100110110110111000101010100010100111110101110001011001001110010100000011010000100011110110110010110000101100111101001100010010101001110101000110110100001110011010000001110001100100111100110101;
#1 $display("%b", po);
# 1  pi=207'b101110110000101100001011001110000011001010101111100101110000000100011010110110101111100011010001000100110100101010111100001100111011011100011000000001011000000101010101100101111011011001000110101101110010011;
#1 $display("%b", po);
# 1  pi=207'b011000101000100010000101010110110111111000101010000101000111100110101101001001000100110001010011011011101000101011100100001001010101101110101101100101000010000111010111010010111000110001001010101100100101101;
#1 $display("%b", po);
# 1  pi=207'b001100100111011111101011100100111011001111101101011011110001111100111100101111011010000101111000001101010101000001110101010111010110010000000110000100100000011110000011000000000000111011101011101111100110110;
#1 $display("%b", po);
# 1  pi=207'b000000001101111011110011110111011001101001111001111100110110111001100110110001011000111110111000110010111010111101011011010000110001101100011101010000010001110101011011010011000011000011011110110000101110010;
#1 $display("%b", po);
# 1  pi=207'b010010111001110010110000110110000011100111101100101100111111110100010100110011000000000100111001010010101111010101010110001011101001000011011110001110001101001011000110000011010000011111110100110000010101101;
#1 $display("%b", po);
# 1  pi=207'b100101110100100111101101001100100001001100001100010010111011110010101001011011101010011001111001111100110100111000100001110001100111010110001101110100010001111001100110000100111001111111000100110100010001101;
#1 $display("%b", po);
# 1  pi=207'b000011110000010011100111100001011000100000101001000111100010001110010101001011011110011000111010100011110110100001000101101011101101100101010011001001011111001000100010010001101011100011100010011111000101100;
#1 $display("%b", po);
# 1  pi=207'b100101100111100110000011111000111000010111110111101001100010100001010101100000110101111111010011110001101111110011101110011101110111111010100110111101111010101011001101000100000111111111001110010010111101001;
#1 $display("%b", po);
# 1  pi=207'b100000011000101011100010011011000100001010100100010000000011011011001111110100000000000001101101100111010001101101011000000110011000100011100100001010011011111100011101101101000111110000100011100110101011011;
#1 $display("%b", po);
# 1  pi=207'b010101101001000110101001010010111000000001100000110010100010110101001001000101001001110110000110001100010101000000010011100110111110000110101100011000001101110100100101101010110011111111111001100100110010001;
#1 $display("%b", po);
# 1  pi=207'b010011000001011100001011011000100111010100000101001111001000111000111100101001100001001000101001001100011001000110011000110010010000010101011001010111011011110010101111011001101110001000111101110111111001001;
#1 $display("%b", po);
# 1  pi=207'b100001101111110110110111101100000011001011101000100101110011010000111001100101001101101100111100011011010001111010101000110100011001111011001010011100101101001001111000011001010110110110010010001001101000101;
#1 $display("%b", po);
# 1  pi=207'b101110011001111101110001100111010001000000101111000010101101010011001001101101111101100010011100001101001100001100001001001111111001010101011000000111000010000110111100110111110001110000001010101100000011110;
#1 $display("%b", po);
# 1  pi=207'b001100010101000001110001110111000110110001000010001010010001101011101010000000100000110100010100110110011010110101100001001000001000100000100111101010011101100001001101011000011101000001011111100110101010111;
#1 $display("%b", po);
# 1  pi=207'b011010101010110011101101010000101011010000011011111110000100100011011101110011011001000111111001010011110111100001001001001110110100101100011111000010111100111000101011101100000111101011011010110100001000000;
#1 $display("%b", po);
# 1  pi=207'b111100101001010011110110010111010010101110101011111000010100111101110000111111010011000010101000001110011100000001001100001001001110011111000100110111010100110110001111001011100000100100001101100001010100101;
#1 $display("%b", po);
# 1  pi=207'b010000111010111000011111001000000001101001110111111010101001010010001110100111111111000111001110101000010100100010110100011101001011110000011111001100111010100110001111001110100101011111100000110111000000101;
#1 $display("%b", po);
# 1  pi=207'b000111101011110001001010011110101111110100110110101010100110001010011000111001110100011111010111100100010101011001111111101110111110111001000111010110000100000111110011000111111110001011110001010111000111001;
#1 $display("%b", po);
# 1  pi=207'b000100010010100100100000110010000110101001001000010001100011101011010000100000001100000011111010100100000101000100010011001110000010000110010001110011100100111000101100110111000001100000111000101100100000000;
#1 $display("%b", po);
# 1  pi=207'b110000110100011101001101001100001111111001100011011010101000111011010111100010010111100111011000000001000111000101010110111011001111111110010100100001101000111011101110101101001000011110100001101101100000011;
#1 $display("%b", po);
# 1  pi=207'b101100000110111000101100001001000110010100001001011000110110111100000010000110010100001100010101001000011111001111101000000111011110101110010100101100001001101110010100011110000011000010101101111011100001110;
#1 $display("%b", po);
# 1  pi=207'b110111000111100000100001010000100011000000001001001010110011011101111111100101010111011110000101110000101010001111110011101010111110100101101011110000111110100011100100101101111110111101101100101011111111000;
#1 $display("%b", po);
# 1  pi=207'b011010101011111111011100010001110101000110101111000111001010011001101010010010110111010101010001010010001011000001001011010110001101010111110100111100011100111100000110010111101111011001111010011011100001010;
#1 $display("%b", po);
# 1  pi=207'b110101001110011100000100001000001111100101110111101101001101010110010001100010001010100101110001000011000011011011010101101000000000110100010110011111010010101111000100000010110111111000000010111111101110011;
#1 $display("%b", po);
# 1  pi=207'b011001001000101100000011111111000111000000110000101110101010110010111111010011010001000011010011100001010011100000000111001111101010001011001001001111011011100110000110100101110101111010101000010100101001100;
#1 $display("%b", po);
# 1  pi=207'b001100000100011001000001011010010111001110010011100111110000011001011000100010110010001000110100011101101000011000011001111010001101101001010100101110011001010110111111101110100100011011100000111110001100111;
#1 $display("%b", po);
# 1  pi=207'b111110011001001110111101101000001001011110111111010011101000000000000010000011001011001110100000000011110001011110110101101101110011111001110011001100110001111111101101100110101110111011001110111001011000010;
#1 $display("%b", po);
# 1  pi=207'b101001001111000001110010101100100100001110001101001000000101001110101111101010100101111110010010101000101101101010001000000000010110100000011011001000101110010110111011100010110001110110110110011011001011001;
#1 $display("%b", po);
# 1  pi=207'b100011011000001111001011001101010000110000000111010000100110111010100111111101100000011000101010011010100110011111101100100000111011010000001010100100001101111100001001111001001011011111101101001101011011010;
#1 $display("%b", po);
# 1  pi=207'b001100010010111000010010000111101001111110100110111001110010100010111101000111010001100101110110010011110011100101100011001110001001011010111000111011111101101110110101101100111111100000110011000101011000001;
#1 $display("%b", po);
# 1  pi=207'b011011100010000101001010001101110010100111110101010110001100011110101010000010011010000010111110101011000110111100101011000010011100101010010110010000000101011000011100100001001001011111011111010001010101010;
#1 $display("%b", po);
# 1  pi=207'b110000100011011001101100101010111010011101100011111011010011000000010111110101100010011101100111110000001010110010000000111101001010010100000000000101100100111100001010110000001110100111010111100000000000001;
#1 $display("%b", po);
# 1  pi=207'b001010100000100010001110000100010001001111110011011101111010000001011000010000111001100011000110110010101011111011101010010101001110001100101001110101101101010010110010110101011110001111110010001001011110011;
#1 $display("%b", po);
# 1  pi=207'b110010110000100001100010011000011001100011001101111001110110100101111111000111100011110110101011110111100111100101111110010010000111111000100110010110111010110001100101011000010101011110110100000111000101011;
#1 $display("%b", po);
# 1  pi=207'b000111110100111111000011000101101100001111001001111011011111110101001101110110000000110011011001010111001101000010011110000111101101011110101011100100110101000011100001101100101000001101011100100100111011111;
#1 $display("%b", po);
# 1  pi=207'b111001000100001011010100010111000000010100111110010010101101011010110010010001110011000011000101101101111101100101111101001010000000101011010110111010010000000111101001110101100111001111000000111110010100010;
#1 $display("%b", po);
# 1  pi=207'b111100000101011110111010001101111000010000100100111011100111101000110110001111100010001001011110001111100000011010001100101000110101010100000100000101000001101001111010100110111001100110100110001100001111010;
#1 $display("%b", po);
# 1  pi=207'b111000110100011011101110111011001100001000010001011001110011100000000111011111110110101100011111110110011001111101100001101111101010101110001101000010011110000111100000111001000100000000001010000001001111110;
#1 $display("%b", po);
# 1  pi=207'b110110000011111000110000101010001010100110111110000111111011101011010101111101111010110100011110101011011111011001111010111101100000110001011000000100100101110011101100000001101010111111001110100110001000000;
#1 $display("%b", po);
# 1  pi=207'b010111011110110011111100011010000011010100011001111100000100000100111111111010000011000011010100110100100100100010000101010011001001010001010010111100110101000101100100011111010000001001111110100010101000111;
#1 $display("%b", po);
# 1  pi=207'b010011101001000100101100110011101001111010011110101010010000011101000010011101101100101110001100100110101010100110110100011111001100000000101111111110001110101011011110011110001001010111010110111101000100111;
#1 $display("%b", po);
# 1  pi=207'b101100101001110110100010101111111110000001100111001010011111111000011110100100001111101111110111101000000100110001111010111110001100110011000100001110001101110111101100001111101001100111110110001101110100111;
#1 $display("%b", po);
# 1  pi=207'b100001011111010001101001001011010101001100111100101110110111000110110011100011101111110111111000000100110100011110101101000100100101011000001100010100101100111000110110111110110001000100000100000110110110101;
#1 $display("%b", po);
# 1  pi=207'b001111111100111011011001000010100101100011010111100111011101010001010010101001001011110110111011011101000011010111110110100000101100011101000000000011111011110100001100010110010101111110000101001010100100000;
#1 $display("%b", po);
# 1  pi=207'b111101111010001010011110110011100000111000111011011000110110101011011111111011110101000011011011111111000001011010000111100111010001101101101010010110100110111000100000000010000110000100001111111011010110011;
#1 $display("%b", po);
# 1  pi=207'b110111011110110101100010100111001111110010000001010000110100001110010001110100010011010011100110001110000000010101001001011011101110011110001110111000000101011101100111010000001010001110011001101001010000110;
#1 $display("%b", po);
# 1  pi=207'b110100010011111101001000000101100100011010000100110110011000111010011000010001111010110001001110010001010100101110100011001000010011000010001011101101100101011110101010111111001111011110010011111011101010100;
#1 $display("%b", po);
# 1  pi=207'b101101001101000100111101101001010001111100000100100011000100000101010100100111111000110110000111111011000111110000100000100111011000100001110011001011111010100100011100110110000010110011110110000100001100000;
#1 $display("%b", po);
# 1  pi=207'b110110101000111001111001110000010100110110011110101111100010000111100111011100001100101111100111100100010100100000110110101000001001011100110001111100001100011011001000110011110001100111101001000001000001101;
#1 $display("%b", po);
# 1  pi=207'b101101000111001001101011110010111001110010001110111010101000010100111111001110001001001101011011000110011011000111010110000011011110001110001101000011110101010001011010101000011111000110001110000000101010010;
#1 $display("%b", po);
# 1  pi=207'b100010010011000011111000010110111100111011111110010001101011100000111100100000111011110011000011011011011010111100110011011101101110000010011011101010101011010001100011001100010010010110011000001101111100011;
#1 $display("%b", po);
# 1  pi=207'b001000011000011111010001010011110000011101111101101111000000110100001110000100000010010101000111000111110111010101010011011010110011110000100101101111100111101010000110100000111101001001100011010110110100111;
#1 $display("%b", po);
# 1  pi=207'b100001101001011110100111000000000101100011110110010000110011101110101001110101111100111011110111100100110010111111111001100010100010100010110010011101100111110100110110111011001100101110011110111111101101011;
#1 $display("%b", po);
# 1  pi=207'b101111100001100000101010110000010110111110001000110010011011111100010000101101101001001010001100100101100101000011010000101101000101111111001001001100101100011111010000000010000110011100010010000011110111010;
#1 $display("%b", po);
# 1  pi=207'b000001010001111001001010110101111110010101000101111011110100110111101001111111001101010100010010011101001100000010111111011111101000110101101100100000001011111001001010010101010011011001101100010010000111011;
#1 $display("%b", po);
# 1  pi=207'b110101100000010110100100001100110111001001010100110110110001100010000001010010001001001111001100110101111111001011000110110001101101100001001100010000110010111010111010010111111010010010010000001100010011010;
#1 $display("%b", po);
# 1  pi=207'b011001000001110000100011011010000011101110111011111011110101000110111001001101001001111101110100011100100011100000110101111001011110100011011011001001011111100000111001001010000010010001011010111010100001011;
#1 $display("%b", po);
# 1  pi=207'b110011100000011011110110111101100101001000101110001010111111001111101100101100001111100000111111101110000111101110100011010100000001111010011111101111110111100111010111010111110110111000111111111111010111110;
#1 $display("%b", po);
# 1  pi=207'b000110100101011101000101000100010101110010001011011010011101101010011100011000000111000001110010111010110100010101101010010101000000101011110101011101000000000011000001010010100001100011101010111010111100101;
#1 $display("%b", po);
# 1  pi=207'b101000100100011111011111011100100110001101101000110000010100111101000101000011011000110000001000001100111100010011110111001111010010011100010010001110011101111100000101100101110010010100100110000100111111010;
#1 $display("%b", po);
# 1  pi=207'b111100111011010010110000100100100010000100111111110010010100101100110101101110111110000000010100011001000101101101110100110010001110010000011110011011000100010000001010011011111010111000100110011110100011111;
#1 $display("%b", po);
# 1  pi=207'b100001011111011110010101010110000110000111100011011111010111000011111001011001100001110000110101101110001000001111011010101111011001111011111111100001011000111100000000011000100100110001111100000100101110110;
#1 $display("%b", po);
# 1  pi=207'b000100010100110111000000010101010101000010000101011111100000011010111110011100111100011101000001011100110101101100111011110001011010111011000111011100101100000011111000110111000111101110001100100011001011011;
#1 $display("%b", po);
# 1  pi=207'b011101111010111010010011010000010011010010100011010110011011100000010011110111001100010000000110000111010011110110001010110010100011110000010101110101001111111101110011011000100101001000110000111001110001011;
#1 $display("%b", po);
# 1  pi=207'b011000111101100101100110001111000111111001010100000111100010001100101110011110000110001001010111010111000000000001100111001111101110110100001110011001110101010101111011011011110101011000100111100111011111001;
#1 $display("%b", po);
# 1  pi=207'b000101010110010110111111100100001001101000100011010100101111100001000101011000111010110111010100000001110111010111011111110101010101111111100111010101000000110000100010001011110001011000110010000111001001000;
#1 $display("%b", po);
# 1  pi=207'b100100101101111100101110011100111100101001100010000100010100000000101101111110000100010001000100001010111110100111101100001000111110110100110110011011000010010001111101010100101001000010000000110001101000101;
#1 $display("%b", po);
# 1  pi=207'b101101001110100011111100011000001101101010011100101111110110000010010111101000010010000100110111111001101000011100110110111100011100110111010010110010101001011010000101011110010010100100000011100011000100001;
#1 $display("%b", po);
# 1  pi=207'b000011101001111011101011101001000011001101110110001001110001001000111001001100000101010001111101110100110001000000111111000110000011000101101101101111001010111110010101000010110011001010011001000111110111000;
#1 $display("%b", po);
# 1  pi=207'b010001000101000101000011010111101000110010010011010101110001110001010011101110010111100111001100111001110001101111100001000001101101010101000010010000101000000110111110000100111111110100011110111011100011000;
#1 $display("%b", po);
# 1  pi=207'b000000000101000100100100101001111110110110111101110001111000110101111000110100000111101011101110011111101101110111100110001101000000010111010111000010100100010100111100000010101000011101101100101011010000101;
#1 $display("%b", po);
# 1  pi=207'b011101001111111001000110101001001011011000110000000011111101000100101101101101011001101000110000110101100100101101111101100101111011100001000011111011001001011000010001010110001101100111110011111100001001011;
#1 $display("%b", po);
# 1  pi=207'b111100101010000100111111001101110001100011101110001110100101100001101100011001111000101111100110010011000110100111110010001001010000010111001011001010001010001110111000111101011100000110101010001010011100100;
#1 $display("%b", po);
# 1  pi=207'b000101000101100000100011100001011101010010000001110101000000111100110111101001111010000100010110010110101000100001110010000101111100010110101111011000111000000110111100101000001001111101010101100111101100001;
#1 $display("%b", po);
# 1  pi=207'b100111101100100001001100111110111100101110111100111010010001010101111001010111110001110011101101101101011101101011000100000111110010010010010011111110100100001000101111010011111110100110100010001010111110100;
#1 $display("%b", po);
# 1  pi=207'b011111010001000010000110000111000110000110100011111101101100111000110100101011111010111011001011110000010001101011101000101101111100010111100111110100000011000111100001110101010001110000111110100100101111100;
#1 $display("%b", po);
# 1  pi=207'b010000110001110101100111110100100001001010111110010101101001110100110011000010110010001100111110110001110001001011100010111101001111010011101010010010110001101001111011011010000100010111001001110100100001001;
#1 $display("%b", po);
# 1  pi=207'b110000011100101011110110010100111000100110101010100101010010101001011001010000010100010010000011100101001111010101100011111111000100101100011100011111011011111110101110110101101001111010011011110101000000111;
#1 $display("%b", po);
# 1  pi=207'b000010101110000011000001111000001000100110010101110010111011100010100001110100111100110010111010000101100001100010011010011100000000010000110111011101001111111011110000110111001000001111110011100101011001100;
#1 $display("%b", po);
# 1  pi=207'b110001000110010110101001100100100100101101110100010110000010000001010100011011001110100110001110101100010101010101001101101111001100010110000101110001111000000001111011010000100110010111101011010101110010010;
#1 $display("%b", po);
# 1  pi=207'b010110110001010100110000010111111010011100111001101000101100011111111000110001100000110010100110000000011101001110100100001110000110011000010101101111110000000001001001001010001111101100100010001100111001100;
#1 $display("%b", po);
# 1  pi=207'b101001101100011100001010001000011111001011101110100111111001011100101001110010000100011111001101100011110000010000000110001010000111010111011101010110110101011111101011101011001001110110011000001010001101010;
#1 $display("%b", po);
# 1  pi=207'b001101111101011101101101110100001111010100001100110001111000111100101101101001101100100101011100010001100110010000100110101111101011101000110011010101100010001001111000001100011011010010110010110000100111111;
#1 $display("%b", po);
# 1  pi=207'b110101101110100000000001100111000001110110111101111000111011101010101100100010001101110100110001110000101101010011001110110010001011001100100100000111000011100110011010110111100100111000010000110001010100101;
#1 $display("%b", po);
# 1  pi=207'b010110011011100110110011001000000110000000100101011010100001110010000110100110110111001001001010001110100010011010001011110010100110101100010110110011001110101001011000100111101001001011010111101101000110101;
#1 $display("%b", po);
# 1  pi=207'b111100000010100011001000100010011110001011111000110001111010010001001010000111111111111111001101000101010100100000010000110010111100010111100011011010000110001100001000001001110111100011100101111101110110101;
#1 $display("%b", po);
# 1  pi=207'b110110111111101010000000110110011111001101010011111010011101101101001110010001011110000101011101000100010001101001011111101010101011111011000001000010101111111011010010111011100000010010011011000010101100010;
#1 $display("%b", po);
# 1  pi=207'b011100011000111010101110000001010101100111110000001100001101001111010110010100110111101110110001111011110001110101000000101100110001111110010000110101110011000010001111111000011111001111101110110100111100001;
#1 $display("%b", po);
# 1  pi=207'b001000010110111000011010100010011101100101011000011101011100010101011001011111011110011010000010110000011101010110100011000000111011010010000100111001010011001101100111110101111011110011000000101000010110101;
#1 $display("%b", po);
# 1  pi=207'b100011001101000011010111001100010110100111101000111011011010010110100001010101111001110000100000101010000000100011000111011100000001100001101101100011001110000011011001010000000000010110110111001101101101010;
#1 $display("%b", po);
# 1  pi=207'b110101011101000111001010001100010101110101001100001001111100011111101001010100001100010101111100101100101001111101001000001101010010000101100100011110111010011111100011101001010010100100100010001110101100101;
#1 $display("%b", po);
# 1  pi=207'b000000101010101101111111000000110000100101000100011101001110000110011001000001101011111111010001100001001011000000110111010010101010111111000100110010011010100001110111010000111100100110011100001001100001001;
#1 $display("%b", po);
# 1  pi=207'b100000011000011100010110000101001100100001010101000100001000000111101011001001011110000011010101101110101110110111011010110010001001001100110101110111010100000110111001100001010111110110001111011111100100010;
#1 $display("%b", po);
# 1  pi=207'b100111100110101010100111101000100011001000010000110111111100111101001101101111010111001100010010111001001011001011000001100100111000000011010001111000010111110111100010000111111000111011111000000110011011010;
#1 $display("%b", po);
# 1  pi=207'b010111110111011110101011011111001100010011000111011110011000000000111100101011011100101100101010000111111110010110100100101110100000101011001000110110110001100001111001100010001100001010010000100000111110100;
#1 $display("%b", po);
# 1  pi=207'b001111110100100011010100001100000011001010110110111110010110111110001001111110100110100111100101101011000101011001100010110001100011011000110000100000000110001111110001110101100110011010111000100001111010011;
#1 $display("%b", po);
# 1  pi=207'b001000111010101100110101000001010001111011111111010111100000011100001100110110000010010111010000001110100000101101111101100000000001010010000111011101100000010000001110010010111011000010011110101111010011111;
#1 $display("%b", po);
# 1  pi=207'b100001000010001010000110010011011010100001010100000110110100100001010110000010110010110110111011010001011110101001100101001110011001001101110101010111100001101101001001001000010000111100000010111111110101000;
#1 $display("%b", po);
# 1  pi=207'b110010100011101001010110111010111110110001000001111100000111110110111101101011110001010111101011010111001111000001101110010010011010101111111010100101101011000001111011011010010100111101101110111011110101110;
#1 $display("%b", po);
# 1  pi=207'b101101111010010001101010011011100010110001001111011010011110011010000111110100111011110111101101110110100001010100011010001100100011000000110100101011011001100011001010110010000000101001100111101010001001000;
#1 $display("%b", po);
# 1  pi=207'b101000011100111100000101010000001001100110100011101000101011110100110111011110011110001000100011100111010111110110001100010011101011000101101010100101111010001000001011010111101111001010010100001111000100110;
#1 $display("%b", po);
# 1  pi=207'b001101110111110111100001110000010100101011111011111011001001111010111101110101000001111000111111111001111101110010101010011001000110110010001110111100010000101001111001100100010110001110100000010000011111100;
#1 $display("%b", po);
# 1  pi=207'b010010110100100010001110110110110001000001100101110100100010110100111101011010010110000001110001010110010111011110111100000111000010000111001111010111101001110100110110000001100011011011010000100100001001111;
#1 $display("%b", po);
# 1  pi=207'b101001001101010111001010001101011101000110000111100010010010010001101100010011101010011001101110000111111001011010001101001110001110100110000111101011001010001100010111100100110001011011010110101111100000001;
#1 $display("%b", po);
# 1  pi=207'b100011100001010010100000110101111111010101110111110101100101111011110011000110011011110011001000011010111110100111101010110010001001110001110001100100001000011100111001010010110011110110010011010100010010110;
#1 $display("%b", po);
# 1  pi=207'b001111000011001010010000101011101110100010011100000101111100101111010100011111111000011001010000111110010100110100000001001010011101001010010000010010100111010111010010010111000011000001100001010010001111001;
#1 $display("%b", po);
# 1  pi=207'b111101000001100101111100011101110100111110011011011100001000001110110010000110111000000100001011000001101100010010000101000100010001001001001000100101011110011000100110011101010000100011100111011110111001101;
#1 $display("%b", po);
# 1  pi=207'b010110101110110110111111010111011111110010101100011011111001010000001100111101001110110101011010011001010011101000010010110100000011110100001100011000010011011000000000101100000011000110000011101000110101011;
#1 $display("%b", po);
# 1  pi=207'b010000011100001011110001100011010000010101101010001001101011100001100111011010011100100111100001100100010010011001101001111111001101011011011001000110101111011011001011101110110011111011100111001110000110000;
#1 $display("%b", po);
# 1  pi=207'b101001001010000001001101100101101110110100010110110011111000011010010000111010001100110011001100001110001111010101010101110110100100010100011011011011010011100010000000110010101101000101010001100111011100110;
#1 $display("%b", po);
# 1  pi=207'b111001000111000010111000000111111001000011000001001101100111110101101110001100010100100110100001001011001011001100100011000110100110010010001001101101011100001000001111000011011111000000011011010011110111100;
#1 $display("%b", po);
# 1  pi=207'b101010101100111000000110100101101110010001101111100010101101000101110101010000100111011100000100100101000010101011100011010100111001010101111000010011100010010011111011111100000111000011110110000000000101100;
#1 $display("%b", po);
# 1  pi=207'b101111101011111100011101110010110100011011110111001010100110000101100111000011111101111000111010011101110100011011011111111110111001100011110011110001111001111001101011100001011011010100011000000111100011110;
#1 $display("%b", po);
# 1  pi=207'b011010110111000001100101000000100101101100010000101100000111100001011000100010101010101010011011111111000000000111000011100110001110000011010000110110111010011110111010011010100000110000000101111101011000110;
#1 $display("%b", po);
# 1  pi=207'b101011111100101001100001000110010101010101111111100110000111001100000001101010100110111011011101010111111011000110110110010010101111010001111000101000001011000001101100010101000110110111010001011111010101000;
#1 $display("%b", po);
# 1  pi=207'b011010011011101000111101001000001001101011000100001100111101101101101100001000001010010100110011010110000010100111101010100100010001011110101110111111001000000000001100101010110110000010110100001010010111001;
#1 $display("%b", po);
# 1  pi=207'b001101100111000001110101001111011011101001000010101000011011010111101111100101001001101001010101100011111011101001111001110011111011111000001000101010100011010001011011101011001010011100101111001000010000101;
#1 $display("%b", po);
# 1  pi=207'b111101000101010010001110101111111011111100001101101110101101111110101010010111111010100010011000110101000111111111001011001011111001101110000011101101101111100111011110010011001101100001111100010011101001110;
#1 $display("%b", po);
# 1  pi=207'b001101000010000100111110100100110001110010000000110000101000100010101111000000100011100100100011011011011111001100100111001100111111011010001010011000101111101101000101001011100010101111000110111010011101100;
#1 $display("%b", po);
# 1  pi=207'b100000101111001011010011100000110101001101111000001101101000110010011010110000000101110111110001011000001110001011010000001001111001001001001010011110101001000001011001001011101110110100010010011100010001010;
#1 $display("%b", po);
# 1  pi=207'b010001101011010100110011011101100010100111001011101111110110000010111111001101110010101100011011100011011011001100111010000100011100000010100101001001011100111000001010001111000001110000010101010010010111010;
#1 $display("%b", po);
# 1  pi=207'b011011101110101010001000101100100000011111100101000011110011000011000011111001111111101100001100010101000100101001001100100101000110101001011011100010001110111110010011001100001100010001110010101000110011111;
#1 $display("%b", po);
# 1  pi=207'b100001011011100110101010010111010110111010010111000100110001111011100011111010011110010010101010011100101011110111000011010110001010111101101100011110101011011011011100010100011001101010111001010010000001010;
#1 $display("%b", po);
# 1  pi=207'b110000100100011011101010100110110100001110010000011000111111010101101010010010100000101011010100111111010000010110010111110111001100101010100111101101101011100010110101101010010100011000101011001010000101111;
#1 $display("%b", po);
# 1  pi=207'b010110011110111001010100011110111111101110101111010100010110110001001110000010011000000100010011100100101101101101100010010010000000101100111100000111010000000001011001100010001001001111111101110110000111111;
#1 $display("%b", po);
# 1  pi=207'b001001100000110100111001100100011000111001011100100010111110111100100000101101010001011011001001011000110011011001001111100000111001111001000010100110100011100111010000000001001100101101100000100101011111101;
#1 $display("%b", po);
# 1  pi=207'b110011111010110100010110101111100010111110110011011111100001000111100010100110101111000100110111100010000100101000001000110100111011110110001100010001100100011110110111110110010110100101110010110011111100000;
#1 $display("%b", po);
# 1  pi=207'b110110100010001011110001010001111111111111000111010101111011001011100100010011001110111111101100000000000010111000100011001011110011011000110000110101101101100111111101101001001010110010100001111101001110100;
#1 $display("%b", po);
# 1  pi=207'b111100111101001101010101010100100110100101111111101001011001011110111010100001010100000100010010100110000100010101000100101101100101110011011001101000010101110110011011101111101101001101110010111101100111001;
#1 $display("%b", po);
# 1  pi=207'b011101011110110010111000010000101111000110011001011101010001010010111101111101000110111111000000101000110011100111001101111110011001101000001011000111111010000110110001110110001111000001101100000101000101000;
#1 $display("%b", po);
# 1  pi=207'b111100011100110111010000001110111110110001010011001110000010111111011000110011101000111110100111101111101000011001010110001101001010000111001010001100100110010011100101000011000011101000001000000010100010100;
#1 $display("%b", po);
# 1  pi=207'b110101101100001001000100111101111000111100000100000010011001001010000011100000001010001101110101000101111000111010111101110101101011010001101010100001111011001100111010100010100101111110111100011011001010111;
#1 $display("%b", po);
# 1  pi=207'b100001100011010111100111010100010110010110110101101111101001110001100111111111001001000111000011010000011000110111001010001011001011000110110111010111100011100011101110011100010100011001010100010000001111000;
#1 $display("%b", po);
# 1  pi=207'b011000001101001111010010001110000101011100100010001011000011111001011000000001011011110011110111010001100000110111000010111101101000100011110111100010101000010010011101000110001010110010001001011101110000001;
#1 $display("%b", po);
# 1  pi=207'b001001000011011000011101011011101100111010110010001011000111101101100101000011010011011100101010100101010000111001111111000010100000010000111110110100111001111101100110000001000010110011101010110110010110001;
#1 $display("%b", po);
# 1  pi=207'b001000111001000011000011100100101101111111101101001111010111000100111011001010111110111101110100001110100100000000011101100001010100101101000110011110101011100110100000011000000101110000010011010011110011011;
#1 $display("%b", po);
# 1  pi=207'b011101111011101111101011110110001010100110011101111111000110000110111111101010100110011011000101100000011001111111110011110010010101101111110001110011000011111101110100101010000000110100010111111101100101110;
#1 $display("%b", po);
# 1  pi=207'b111101100001110001100010110001010010100100110011111101000000010000011011010101111000100111100100000000001001001110001110000000010000101111000011100011010100010001110001010011111101001101001011001010101100101;
#1 $display("%b", po);
# 1  pi=207'b010011001111110000111011000111001100100111101111111000010000010101110100101110001010110101111100000011010010101111110010001001011011110010100000000100111000101101110000100101010101000111111010110101011001010;
#1 $display("%b", po);
# 1  pi=207'b111000100111110101110101111000101100111000101010010001001110011101110010110011111010001101010100001101100101000011101011010000100000111111100111111000000000010101010000010001010011111100100110111010111011110;
#1 $display("%b", po);
# 1  pi=207'b110001110011110000101010010010101100010101110001110011011000010101011011000100010011100000010100000111101000001010011111011110011011010000001010010001001010101110111100011000001000011111110011001100101001000;
#1 $display("%b", po);
# 1  pi=207'b011001011000110111101011010000000000100011110000111100110110110011011011111000001100100000001110010100011101111101101100110011010100101100010010100011011111101110110000000011110001001001110111001001101011001;
#1 $display("%b", po);
# 1  pi=207'b111011110000001111010011000011000111110101101000101100001010010001011011011010110000110010100001001000010100000000111011011111100010101001010001000001010101111010100000110110110000111111011000000000110110000;
#1 $display("%b", po);
# 1  pi=207'b111111010100000001010000010010101111110111001011011111111011011111011010011110010000010010010000100011001001110100011110111010101011100010110110011100011100001111111101110001100010101001000000010101100000011;
#1 $display("%b", po);
# 1  pi=207'b100100010011000001011011001111101110111110110111110000101010111101000011111010011001010110111001101000000000000010111001101001011001000101001101110000000000000110001001011100001100110011101001011010101011011;
#1 $display("%b", po);
# 1  pi=207'b100111010000011111000100011011110011100110010011100000111010010000010011111000000010010011010101010111000011101000001101110100000010010010011101001111101011011000101011100010111110101001011100100101001110110;
#1 $display("%b", po);
# 1  pi=207'b011111100001000110011100110111101101111000110101111000110000001111001100110000000110010101111110111001011100000000000001010111101100111001010111000011011110110010111010011100000101011111001011001001001101111;
#1 $display("%b", po);
# 1  pi=207'b100010111101001000011001011111110110100101011000000011100010000111110010101100010001000110000010011001111101000101111010010011110110100000011011011101111000000110010010001011000001101001001100011110111101101;
#1 $display("%b", po);
# 1  pi=207'b110000001010010010100011000110011001011001111001010110101001011011001011111010000010101000000011001110010000111001100110011110110111101010100000000100000111011111101110011010111100110110100001100001010110000;
#1 $display("%b", po);
# 1  pi=207'b010001000000110111110010101001110000011000110001111101001100101000101111000100001001010010001100010100010011010111011110001000111010111010001101110011110110010010011100101000010011010100101100011110111010000;
#1 $display("%b", po);
# 1  pi=207'b001101001010000111101101101000111001010111110001111101111110100010010000110100100010001110001011000101110010111001100001001100010101111000110000011011000110010110100111001000111111101100010111101110010110000;
#1 $display("%b", po);
# 1  pi=207'b100111110001001100100011011010110111101000111010111010001110111001111000111001100011011001011110010110010000110010000010110100101001010110010010100000010010011001000111010010100111001011011011111101000100101;
#1 $display("%b", po);
# 1  pi=207'b110111111001101100001000101101010111001111100001001001001101101101001011111011110001110110100111001001011101111010100110110100010001101001010000001100110100110011001101110011100000110110011010011100000101101;
#1 $display("%b", po);
# 1  pi=207'b000111111111010010000010001110011010100001111101011010100011001111010000010000110001101101110111010111100110011111001001001001110010101100101110100101000100000111111010111101000110111101010110000111000110001;
#1 $display("%b", po);
# 1  pi=207'b111010110101100001111011101100001100000111000011000000001001010110001000011100110110111100111101001011001111001111111100111100011100100100010100000000000010110001111010110100010101000010001011010111110000111;
#1 $display("%b", po);
# 1  pi=207'b001001100001000011110110101110111100010000111101011100001010000100111101110001000011101011101101000110111000101101101011000111110000000001111101000010001001100100110010111111010000110000011110111110001111011;
#1 $display("%b", po);
# 1  pi=207'b101101101110101001011101100010010000111110001111000011000110000010010100011000000110001011000010010111010001010111011000011001100101010100111011001100010111100100010111100110011110111101110111100110110010100;
#1 $display("%b", po);
# 1  pi=207'b100100001010100101101111110000001011000010000101001010100111011101011011101001011011001011001111011101011100010010000101110011000111010100110101100101001001100111101011110101010110000000000101010101111111000;
#1 $display("%b", po);
# 1  pi=207'b111101110010010101010101111001010100000100000001010111001111101000100000000001001000001001001010001110100111100001100011001101110011101101100111010011101111000011110011111011111110111110010001111010000000110;
#1 $display("%b", po);
# 1  pi=207'b001010000010000101010011110100010111110010101100101010101010100000111101011011011000001111000001101101100111010110100111101011111101000000011110110101000110001100100110000101100010111101011010100010010101110;
#1 $display("%b", po);
# 1  pi=207'b010110101101010110110010100010001001111110001011100100010100101011011001101011110110110011100100111011000101110110011000101110011111000000010111111101000000001000001100111000101000110011000001110101111010111;
#1 $display("%b", po);
# 1  pi=207'b110011101000001000101111101000011010101101011111111010110001101011010110000101110111110100010110101011111001101001010001011101111010101000111011101100000101010110010010010110010011001111001110010001100111110;
#1 $display("%b", po);
# 1  pi=207'b110110101111111010010010011110110111010110100110011011000000110110000011010000001110010110110101001101111001000000100110110101010101011001111110001010111111100010010111110111000101101010100001101111101101001;
#1 $display("%b", po);
# 1  pi=207'b001111011001000011011101111100010001101111101111011001100100011111010100100011100000001001111110001100101010100110111001001100100100101111100010010110011101111111001001001100101011010000000111100100001100110;
#1 $display("%b", po);
# 1  pi=207'b011110011001001100110011110011000010000100110110100010100000000100001001100110000011100100000100001101011101010011100001010010101010011100100101100000011000110011011110010000001000111110000010010001011010000;
#1 $display("%b", po);
# 1  pi=207'b110001110101100011110010011011110111000110000011011101111111000011001000110111000100001111101101011010110100111010010010001011111110110100110000000101101100101000111111011001101110001011100010000101100011101;
#1 $display("%b", po);
# 1  pi=207'b110001010001110000010010001100101110111110011011010011001111111111010100000110001000010101000010101010110000011011001001110001101101010010111000101001000110100001100110111000011000110010010010000010111010001;
#1 $display("%b", po);
# 1  pi=207'b110011100111100100010001111110111000001100010000100111011010000000011111100100111001100111111000101111001000000000001001110100111000101110010110011100110100010111001100001110100011111101000000111101000111110;
#1 $display("%b", po);
# 1  pi=207'b011011101000000000111101111000111110001000101011100010110111110110111101101000000101000111100000001010000110001110001100110011010010000001111110101000101000100001100001100110000001010000011110101100100011010;
#1 $display("%b", po);
# 1  pi=207'b100000111111110001011000101110011101100100111001011101110010111001000111110110111010001100010011000001010100001110011110011001000100111100111110010111010101111010001001011011101001000001110100101010011000000;
#1 $display("%b", po);
# 1  pi=207'b011000111000010000001001110101110111001011011101001111110110010001001010010001001001001100000101100111010100111111100000111010110111010010000011100011011101100111000110110010101000111111000001000001101011001;
#1 $display("%b", po);
# 1  pi=207'b100100111111000100010101110111101110001111010001111011100111101111000001001100001001110101100111100000000010110101110011110100010011101011000010011001100000010110101001001001100110111110000101100011001110101;
#1 $display("%b", po);
# 1  pi=207'b011100110110011101101111000010011110101111010110100100011001000001111101110011101100111000110100010111001101110001100101011101101101010000110010100110110111001100010101001101100111011011010110111110100010101;
#1 $display("%b", po);
# 1  pi=207'b100001000100100110110110001110011011110000101011000001000110010100100011000010100101100101011101010111001101001010010011010110000010100010100111110110010001101001001110000011011011111000101111101000001010101;
#1 $display("%b", po);
# 1  pi=207'b000111101101111001101010100011110011101110000111010001110100110101110010111011110001101000010010010010100110001011100110110101110110011000101111101100101010000000001001001001111010010100101111011110110110100;
#1 $display("%b", po);
# 1  pi=207'b010011010010110110001011001100100000101101011000000100010101000010111001001101101000111000011110011001100001110110101001000111011011001000100100010110110111110110000001101000100100010111000111010011110011000;
#1 $display("%b", po);
# 1  pi=207'b001101001111011100111100101011001110111100011011000001110010001000000110111110111110001011111000100010011000111110110110010110000010110011110000110010010011111011001011110111010111100100001110000110101001110;
#1 $display("%b", po);
# 1  pi=207'b100010111101001100100011111010110100001000100110101000001101110000100110100101011110000101110110000100011101011010110000110011001111100110100001111110001011001111010011011110010001011010111111010011010010100;
#1 $display("%b", po);
# 1  pi=207'b001000010000100010001001011011000010110000011000010011101100010100110010010111110111010001010101101011010111010000010110110100010011110111011010100100010011010111001001001010101101111100110000001111010000111;
#1 $display("%b", po);
# 1  pi=207'b100000010110110110101110111011010011001110100010001000111000000010111110111101010010010100110011000010101111000100110000001111011101110101010010001111010000100111001110001011010010110001110111001101110011010;
#1 $display("%b", po);
# 1  pi=207'b110000101010100100010010001110100110000000000001110101001011100000001011111110100110100110100010001101111000100001001110111101100101111111100011001010100011100011101110111111010000001111000000001000111011000;
#1 $display("%b", po);
# 1  pi=207'b100011011111000010110111111010110110010000001100010110010101001101001100001111111111011101101111100011101110101110010010111011001110111100010000010101000010110100010001110110011110001000001001000000001011110;
#1 $display("%b", po);
# 1  pi=207'b101000110111011001111001010001000011101110101011011111101101101101100000000110011000101011001010100010001001110001110111100000111111011111001001011010100000100101100000111110000010000000010110100010110100001;
#1 $display("%b", po);
# 1  pi=207'b111111000100000111100011010110000100101011101000110100001011110110000110011001000101010010110111100111110000000010000000011110101000101100100000100110110100110010101111001001100101010010011101111100101011010;
#1 $display("%b", po);
# 1  pi=207'b000010001111101101001110110101111101100010111111001100100000001001011010111111110110011001100000110110111110110101111001010100111011101101001100110110111101100111000110110011101100000101011011001111001001111;
#1 $display("%b", po);
# 1  pi=207'b010010010101010110011010110010011110100010111000000001111110100100010100110100011110100010100010100110111010101101011001110111101001011000010000000011010111001110000001100010001010001001100111100111101101001;
#1 $display("%b", po);
# 1  pi=207'b001011111101001110011010000100001100001011111001111101101010000010001011111000010100011100011101010101100100011101101011111000110111100010011100101110011000100100110001000010001111000000000001111010000001110;
#1 $display("%b", po);
# 1  pi=207'b000101011110011011000110001001110101111101110100101110010000001010111000011010111100011100011111100000000010111011110111100101100101100011110001001010101110111110110101000100100011101001000001000100101010011;
#1 $display("%b", po);
# 1  pi=207'b111100111011110011001000011111110101100000110111111111011001011001111011100001101101111110011011010111011110001101011111100110010100110101110110100100001101000010110101100101110011110000001100010101111011001;
#1 $display("%b", po);
# 1  pi=207'b010101110100101101001110001111110101110001100001100100111000101001100000101010001101001110010011110111000001111001110010001000111010010011100110100000101110111010101101110100000011011100101010010000111111000;
#1 $display("%b", po);
# 1  pi=207'b011111101010010101100010001011101100101110010111001100011101011000101111011110111101111110101110101010100000100110100100110101101111000011111101110011011110100010110101100001010100010110010010011100010100101;
#1 $display("%b", po);
# 1  pi=207'b111100001100100001111010010110111110101011001110100100111111011111000001001111011100011111100110110111111111111001001000100000100111101111100101011100001010100110110111111101110101110011011100100100110101100;
#1 $display("%b", po);
# 1  pi=207'b000111111100111111011001001100110011110101111010111000000000100010000101101111101110011110101111110001000010010001010000100110111100010100011000100001001101101100110101000101100010001001001010010100000011101;
#1 $display("%b", po);
# 1  pi=207'b010101111110001101101111111111100110000000111010111100010111111111110101000111100000000101111101100011001111110011010101011000101001101101001001011101100011111100101101100111001000110000101100000100101011111;
#1 $display("%b", po);
# 1  pi=207'b100111100100100000010110010001001111111111001110111000100100000110001010000100010100110101101101111001101101111101110111101110111010000100010100001111100101101110000000000110100101000110101011010110001001101;
#1 $display("%b", po);
# 1  pi=207'b001101000011100110001111111101111100010101001011010000101011001011001100111000110111101001110111001000010100010100111101000011001011001001000001110010001110110000001001111001110001101010001001011110101000001;
#1 $display("%b", po);
# 1  pi=207'b110111111111011011111010000110101001010000101010101101110010110100100100001011011101111010111100101100110111001001000101100010001111011011100000011110101100010010100100110001101010110001101110100111101101000;
#1 $display("%b", po);
# 1  pi=207'b101110010111000000100010110100001000101001110111000010110001100001010011111111000100101110000111001000111110101001111010101111001010010001110100000001101101111010000100100101100110111000000001000000000010101;
#1 $display("%b", po);
# 1  pi=207'b101011011110000100010111011110111000101110011000001010111010001101010111000111000110111000100101010000010101001011010111000010010111111111000011111010101010010011011101011110110011110001110110101110110100101;
#1 $display("%b", po);
# 1  pi=207'b000010101110010101110100011100011111110101101001101100110100001110010010100110101111001000111100001001001011110100001100001011101110001001011001100110010001111110011011110000111100111101111100011000100000111;
#1 $display("%b", po);
# 1  pi=207'b000111101100010001000010000011111100000001100010110111110111001001101010101111101111100111110101110101101001111110011101011100101100010010000111100100000101110100010101100010000000011010111110100011000000100;
#1 $display("%b", po);
# 1  pi=207'b110011000111101011101011011100100101110010100000101000100010011110011100101000111101000010111000011010110101011001111010000101011110001111000101100111111000001011111100111100001101100111110000110000011101111;
#1 $display("%b", po);
# 1  pi=207'b100000011100010101111000010110001000111100100100110100110000010101000101100110101111110011100001111000100110100110001111010000111100100100111100111100010110110101010110110000110100011110110011111111000001000;
#1 $display("%b", po);
# 1  pi=207'b101010000100111111010110001111110101010111010100101111110101100011110010010101000111110000111001100100001101110001110001110101111000110011011111011111001111111111111011110000101000110001011110100000010000110;
#1 $display("%b", po);
# 1  pi=207'b001110110111011101110100010010110011001011010111010000000011011111100010111011100010100111001001000110111001000111111101000010010101110011110011101010110000100111010001000101110100101101110111000100101110110;
#1 $display("%b", po);
# 1  pi=207'b100101000000001110001001000010111101010001011111001100011101001100000101101101011000001100011101011001001010111011110110111110100000010111101010110010110001010001011000101111100000110100110001001011100000010;
#1 $display("%b", po);
# 1  pi=207'b011111000111110110110011010110110001111100110101110111010101000010101100101011110110110000110010100011110000110011010111000111111111001110101000001111111011011000100100011111110101010010010001001010100001001;
#1 $display("%b", po);
# 1  pi=207'b000010110110110011010110011000011110001101000011010110010100010111111110110000000011101111111011100101110001001001000110011110001100001000111101001011011101001010111101011001001101001011100000101001001010111;
#1 $display("%b", po);
# 1  pi=207'b011011000001001001001010000000100000010100011001010100011001111100111011110101010100001011101010001100101100110111101100001000000000000011110000101110100101010011111110110101111001011111001100101000000101000;
#1 $display("%b", po);
# 1  pi=207'b000000011000101101111110111011111010101110110010100100010001110011011011011101101101111100000000110111110101001111011001000001001011001001010011000001001000010000110101111100001010110010000111001101001010000;
#1 $display("%b", po);
# 1  pi=207'b111001110010000111100100000111101111000100010110111110010111011110111001001000010010111101010001111100010000001101000001010111101100000010100000010000100001110111011000001101111110101101111010001111000001101;
#1 $display("%b", po);
# 1  pi=207'b011100010001101011001100100010110001010101100000101010011000000100011010010001111011100101001001101111111010010001111001101011001100111000010101011100101101000101110000110100010010001101010001110100001011000;
#1 $display("%b", po);
# 1  pi=207'b110001000100011110100111011110101101110100010111111010001000001110111000100100000001100111100000101101111101111010111101100101110001000010100100001010010011011111111000101110101110101111100101100111111101010;
#1 $display("%b", po);
# 1  pi=207'b100100001111010110111111101000101110101110101000100011000001111100010000011111111011110011111011001100011100000110111111110010100110110000001100100110110001111111110110101010100101101001010111000111110101101;
#1 $display("%b", po);
# 1  pi=207'b101110111000100011000100010001111111010000100011101011110111100001000110111101111000101000000101111101001010101110111001000100111110100000100111100100011001111010010110111100101000001001000110010100001001011;
#1 $display("%b", po);
# 1  pi=207'b001001100000011010011001100101010100011000111111101011011110001011111100100001101000001010100010100111011000011101011000110000101111011100100011101000011101000101110100000101110000100100111100110101000001100;
#1 $display("%b", po);
# 1  pi=207'b100011111100100111010011110011001010001010011110101110000110110001111000100010001101001011110011111011011010111011101110101110011011010110110110100110110110100111111001111011101110001111100011111100110001011;
#1 $display("%b", po);
# 1  pi=207'b010011100110101010001101000100100001110101000111100101010010010110011101110111000001101010110000100010111000001101111011111101000011011010111000111101001000010000100011010100100100101101001100010101111000110;
#1 $display("%b", po);
# 1  pi=207'b101000111110100011001100100111010001011111011010001111001000100000111100000001010111111001101011101010010011010111011011001110101010011100100110001011001110000011100010110000000010000000111111010100000000011;
#1 $display("%b", po);
# 1  pi=207'b001100110011101010110011100110100000000010111001001001011000100101011111100101010001000101010100001110100000101011011101101000111110000001011110111111110000111100111111110001100111001000010111110100000101010;
#1 $display("%b", po);
# 1  pi=207'b011010111000011010001010101011110101001010000111101000100100011011011100111011000011110111101000100001100111000101001010100100000100000110011000110010001010111000100100101111100110000010100011010010101000100;
#1 $display("%b", po);
# 1  pi=207'b101101011010000011111111001101001011011100100111011000011101001010101011010011100001110101100110101110101010101101000110001110010100110111011110010000011110111000011011001000110101111100001111100110111010100;
#1 $display("%b", po);
# 1  pi=207'b111010011010010001011100010101111000111101000000111101111011110010010100000100100011011101011110010100111111110000110111111101011000011000010111100011010000000011110110001001000100001100001110001110011111111;
#1 $display("%b", po);
# 1  pi=207'b100101011110110011111010010001101001111000001000111000011011110111110111100011110111011001001010101101100111100101100111110001101110100100111001000011101010111000011010010011011110101110010110100000000001010;
#1 $display("%b", po);
# 1  pi=207'b111000000100011110010010111101001110111011000011100101000001000111100111010001111101000011101010001001101011111110001011111000110101100110110110000001011000000100111001111011010111011011000111000100010011001;
#1 $display("%b", po);
# 1  pi=207'b000110010010000100100000100010110100101000000111110011001111100000001101010101011010111100011000111000101111001001111111011010010001000100000001101010000010100111010000000100101110011010101001000100101110001;
#1 $display("%b", po);
# 1  pi=207'b111111011110000000100101010000100110001111110101001101001101010110111110010110110001001001010011111000100101011000101010111111001101010001100001010110010100110100000001101111000001010000011011111010100010000;
#1 $display("%b", po);
# 1  pi=207'b101011111000011111100011110101110011101001010111101011001010000100000010001011111111101100010000011100100110111100011100100101100010111011101001101101100000101101110010011100110101110011111011111001100000111;
#1 $display("%b", po);
# 1  pi=207'b001110011101010111101110111011011000101101000001011111010000111111001000000000010111011101100100010001111000110101110100000011001000110000101011011100000010000011100000001001011111000100000101001001101010110;
#1 $display("%b", po);
# 1  pi=207'b001001100101000011010111011010101000100100111011111011111110011101100110111110010011000011000010011011010111101101011000011110101000100110101110100111010111010111000101011011111001101010111010001111010000011;
#1 $display("%b", po);
# 1  pi=207'b010011110010111100000001000000001101011011111010110110000001011001100000111110010101001001100011101011000100101011000101101000000010101011101111100000111011001110111010101111111000001010010110110100011101100;
#1 $display("%b", po);
# 1  pi=207'b010101001111100010101100001001011100100100111110100001011010001000000100010010110101100011011011111010010100001110111101101111000111010010100111010101101001010111111001011110110001101110111111110000111010111;
#1 $display("%b", po);
# 1  pi=207'b010101000110101000001001100001010011100001111000111011010101001110011110110110001001100101010111011101011010011000101011111100000001101110100111001001001111101101101110001000101110000011011110000001100110111;
#1 $display("%b", po);
# 1  pi=207'b111110111100110110010110101111100110100100111100001101000100000110101101111100100110101110011011110101000111101010000001111111110100010101001001000000100101100010011101001111111100110110100101110100001101101;
#1 $display("%b", po);
# 1  pi=207'b001101001100011011100110110000011001001100110010000111011000110110010001110100101111110100111111101100111100111001001111000011011011011101011111001000010100001100111101101111111010010101001001010000000100111;
#1 $display("%b", po);
# 1  pi=207'b111000110100110010000110110000001110100100100110010110001000111110010000101101110001001010010001011100000011100001010011100111101010001101111010010101010010101100111000000100000010111101100101011110011000001;
#1 $display("%b", po);
# 1  pi=207'b110000011011101011100001101011011011111100101100110011110100100010010000011000000101111111001001100100100010010110111001001011010111101111000110110000101110011010011010011110001100100001100100000110100001100;
#1 $display("%b", po);
# 1  pi=207'b100000110111010111001011000000110110001010101000011110001001110110111100101011101101000011101010000101111101100000110000011000001010001001101001100000001010011100111001011011001110011101110011100100001010110;
#1 $display("%b", po);
# 1  pi=207'b110001001010000111010100100011111101011101001111101010011110100111000100111010101101011101110110010011101001100001110011110101110101011111001011110111010011101100011111100000101111010000111010010101010111111;
#1 $display("%b", po);
# 1  pi=207'b011001010001011000010111101111101000100101001010001101000010001101011010000110011111110000010111110111010101001001101010101000011100100010010010110111000111000010100011011010101100000100001000110000111010011;
#1 $display("%b", po);
# 1  pi=207'b011111110100010111011000101010111010011001110100000100000010100100001111111010010101111010000111001110011001000100001001110111111100000011010000011101110000011010110010001110100001010110100101101101011010001;
#1 $display("%b", po);
# 1  pi=207'b101001000011000111000001001001110101011010001100000000000101111110110101000000101001100010001001010101101101010111011111001100000111011011000011001011000110101010100101100010011000111101010101011100011100011;
#1 $display("%b", po);
# 1  pi=207'b001000100010011101010000110001001101101100000000010110111111010111100110110000110101000001111001000100000000101110111010101010000000111000110100001011010100000101011110000010000110001110110110010110111110011;
#1 $display("%b", po);
# 1  pi=207'b110101001101100010010100101000010111110100001101000001000011001010110011010000110010110001010001111000110110100101110110010010101011101101010001101010001010000111100011000100010101001000111100101001000100001;
#1 $display("%b", po);
# 1  pi=207'b001110001100010011010001001010011000001100001100000111111011100000001100111000111000111101010111101100011100111011000111100010110110010010001110010111111111000011100001011110111001101111101110011010110110010;
#1 $display("%b", po);
# 1  pi=207'b111101101010001110111101011000111001111100101000111010001010100000100010101011010110110000001011010011100101010110000100010110110111000011001111111010000110011100100101100010111010011010110111011011111000000;
#1 $display("%b", po);
# 1  pi=207'b000101110010101000010011010000111110011010110100101110011000100001100011011001011001110101011001001111110111001100010111100001010111100000011110110101000011101100100000010100101110110000101110000011100010010;
#1 $display("%b", po);
# 1  pi=207'b000011101110001101101011000100111110100010100000010001011100010111000110111011011100110010100111111000011111110010111011110110101100110101100100001111001101001110010011000010101011001011101100110010100001010;
#1 $display("%b", po);
# 1  pi=207'b011010001101001011011111101011010110110110101001100000001111110001010111001110110100000000111111111110100010011000111111101000001000110101101010111111001101100101010100000111110011101111000001101100000000001;
#1 $display("%b", po);
# 1  pi=207'b010000011111011111110011100110101010001100010001011001011001001000100000101001111001001101000101001100110110000010000010100101110011011100011111111111101100010100100101100011000111010100101110100110000111001;
#1 $display("%b", po);
# 1  pi=207'b011110111101001001101101011001111101110110100101100010111110101011111010100001110010000001011001000011000100101111110000011100111111001001100010000001111101101000100001100111000111101111111101011011111000110;
#1 $display("%b", po);
# 1  pi=207'b011010101101111111011001000101011100111010011111100100101100110101000000100100111101010011111011101001011101111101000010001100110110101101110110000010000100110000100110010111100000011001101001011010110001001;
#1 $display("%b", po);
# 1  pi=207'b111000001000100100000011110011011011110001000100001000100001010001111111010001001011110111100001010101000110111110111110100011101001011011101101110101101000101111010100100101011001000011110011000110100110100;
#1 $display("%b", po);
# 1  pi=207'b010110000011010111101100011110001001010001001010010001011110001111011000110011111001010011000111111010110100110110000111101101011010110001101110011000001001010100000100001000100100011001001010010110100011111;
#1 $display("%b", po);
# 1  pi=207'b111000101111010100010011011011001011111101010100000011100101001110011100011001001001011100010110010001001010010111000101011010110110100110101101000001100011111001010001110101011000111110111011010001001101110;
#1 $display("%b", po);
# 1  pi=207'b110111000111011000111110000010010000111010111000101110111010111101111111000110100010000100111100000000011110111001111011001010101111011110001111011101111000110011101011011001100110001011011110111011111010111;
#1 $display("%b", po);
# 1  pi=207'b101111110011010101010001010111001010111011100011001010100011110010111101001000110010000000110000111010111100001100101001110101011100110100000111110111001010101101100011100000000001100111100111010101011010111;
#1 $display("%b", po);
# 1  pi=207'b111100111110110111001010011111010010010111101100111010011100111100000011001111011100101110010111000111001111001101011010011110001001011111010110101000000101001000010100010000001011101101001111100000101101110;
#1 $display("%b", po);
# 1  pi=207'b101100110100011010010001001010000001110100011110100111011000101101001011100110101010100010010001110110011110010000101110111100001010001111001111110100101100111111101101000000001011010001010000110101111100110;
#1 $display("%b", po);
# 1  pi=207'b011001010011011001010011110010100111001101001010111000100100000010101001111001110001000010100001011110000001111001010011101011010110000111000110010110111011100101100100001001111101110111011111110011000011001;
#1 $display("%b", po);
# 1  pi=207'b101001111101010001010111010001001011011110001110011011111101011011100111100101101100011010101101100000000111000010111101000000011001001001010010011001101101111011000110111000111011000110010010010010001100000;
#1 $display("%b", po);
# 1  pi=207'b111111010011100010111100111011101110011001000011000111011001100111101000101011101100100001010000101010101001100001110010110011100100011110000001000010000011101001000011100001111010101010100111101100100110001;
#1 $display("%b", po);
# 1  pi=207'b000000001101100000101110000111101110010101011100110011001010110011110110111101010101111110100010011000000011110110000010111111000000000010101110101111011101011101100001100010001011001100001110000011101000001;
#1 $display("%b", po);
# 1  pi=207'b011000100100111011001011000110011000001010011000101000000000101100111100000000010000100101111010100100010010000011011010111101100110010100011010110100010110000001111001010011000010101100111000010011011110010;
#1 $display("%b", po);
# 1  pi=207'b001100100010111000010011110000111110110100111011111011010001111010001100000000100101011100110000001101011001101111111110100011101111001011001011010111000010110010110010001010101001101010101010001101101000100;
#1 $display("%b", po);
# 1  pi=207'b010100011111110101111011110111010100101011010110110100001001110000100010011010110111011001110111110001000001101000101111110010100101110110010110101101110011011001111101000100101011000101001011000000000001110;
#1 $display("%b", po);
# 1  pi=207'b100011011011010000110110010110000111011111011011100010111100000101101011011101100100001101111010001001001000111010011010100101000011111011011010111111100011001000100000000101111011111110001010100100010010011;
#1 $display("%b", po);
# 1  pi=207'b111011001110010100110100111110011000001001101111000110100110101100011000011110100100100000001011000111000111110101011100001110010110001110011001010111000001010010101000011000000110011110110001000011110000010;
#1 $display("%b", po);
# 1  pi=207'b101010111000011001000100010001111111011110100100000011010101010100010001010000001010110111111001000100111110011010110110000011100001010110111101011010000010010111101011000011000000011000111110010111111111100;
#1 $display("%b", po);
# 1  pi=207'b001001111101110001001110011101010110011101010100100101100100001101010110111010100011100111001110010001001100001001111111101000001010111100001101101100001000101111100110001101110101011110111001001001101000001;
#1 $display("%b", po);
# 1  pi=207'b101010000110010000100110001111110010111110011100010001011000110100110001100111111000011100010001110001001101101000000101011111000110010010100111101110001100001001000001110100001000010000000011110100110100110;
#1 $display("%b", po);
# 1  pi=207'b101110000100101110101110110110010001011000000101001100110010001010110011011001000011110001111011110001001010110101110010111101100011011111001100111100001011100001111110101111010000100101000101111111101111011;
#1 $display("%b", po);
# 1  pi=207'b111000010000111000011101100001011111101001000101110001110001101101101001101001011100100010101001101011101111100001100100100001011000101011110010010000000100101100111110010111010101011001100001111000000111010;
#1 $display("%b", po);
# 1  pi=207'b100110100110010001110101001100010000111101100011111000101101001011100010110100001100000010011010100100101011101100111011111101010010101110101100101101011011101010011101001000111010001000100011001110011001000;
#1 $display("%b", po);
# 1  pi=207'b001110010101001001111101110100101110111100111001001100001110011111100000010001101110001010111011001110001010101100011101110011010001010001011101111010110010010101100100001110101001010101011000011011100011110;
#1 $display("%b", po);
# 1  pi=207'b100000010111101110011110110101000010111011111111000110101010000011111110010001000100011111111001001000001101001010010010011011001001110001100000101001001110101111010110011000001110100101101001000001100110100;
#1 $display("%b", po);
# 1  pi=207'b100101111100111000010001000101110010100000001010010110101111110001010100000110000101010011000010000111100101001001111000110111111011000010100101010000110111101111111110000010101000010100110010111011101110101;
#1 $display("%b", po);
# 1  pi=207'b000111101111101100111101101001101011101000010011000100101111000111010101101111101000000001100111001111111101110111100110111101110110111001010111011011110101010000100100000111111110011001011000100011000000011;
#1 $display("%b", po);
# 1  pi=207'b011111001110010011010111010010011010011111101100001100011110110101011000000010011100100010100000101110101011000100111011000101000101110101110101000001111011100001111011011111001111110000011010111001001010011;
#1 $display("%b", po);
# 1  pi=207'b100100011111001011011011011111111010110000100001001110010000000110101001000100100100101111101010011010001000111001111101010010001101111010000000000110100001000000101101100000010011110111010110111001100010101;
#1 $display("%b", po);
# 1  pi=207'b111001111110101011011111100001010000100011010111011111111001100101111111110100011110111001010010001101000101001101011010001001100000011010110111010101011000101011000110110001101000000010100100001001001011001;
#1 $display("%b", po);
# 1  pi=207'b111000001101010110001101001101010100111000101100010110100101010111100101000100010000001011101101001001000000101110000101011110000110001101100011010100000011011000100010000001000011110001110010111111100001100;
#1 $display("%b", po);
# 1  pi=207'b010001110010100010101100001010111110100010111100000111111111110100111000101010101011000110101000010111001010111100111101101110010010001000001111000110010111000110010110101000011010110101000001001011101010000;
#1 $display("%b", po);
# 1  pi=207'b010101100111000000111010000100111111100011001001000110010111110011001000010010111100011000010011000000100001110101010111110001010001001001110111100011111010100011001111000101111001111111011010101011110110001;
#1 $display("%b", po);
# 1  pi=207'b110000100110101011101011101110100010011000011000001010010110011101011000110100110010010011101000001101011101011000000101001111111110101111001001000100000011011000100011010111000001100011011000000000000011010;
#1 $display("%b", po);
# 1  pi=207'b110111010110000011010110110011110010000101000111100110010111011001011010110111011111011010011111000011011000011010101001010110011111010010101111111011001011101000000100000101011101111001111010100110100101100;
#1 $display("%b", po);
# 1  pi=207'b100110101010101100000000111011001010101011111110101001001101001000000110001001000011010110110010111011110010111111000011011011010010011010011111011110010000001101100100010011101111000100010100100110001010111;
#1 $display("%b", po);
# 1  pi=207'b111100010100110010101011011011001000010111100010010101110100000000010111011110110001000101011101101101001110011011010101111001100010110010111101001001110010000101110001011011110011101111101111000100000100001;
#1 $display("%b", po);
# 1  pi=207'b110000110010100010101010101011110100010011000000001111000011100011111100100101011010010101010010001100110010111001010011100101000100100001011110000100111100000000101110111011011101111110110111001100100110110;
#1 $display("%b", po);
# 1  pi=207'b100101000110010000100110111100111011000010000001001110010100110101011000001010010010111110000010111100101001011001101110100101010111001111100010111110010111000101110001111111010110000111111100100101110101011;
#1 $display("%b", po);
# 1  pi=207'b110000100111001011111011111111001010010011011100010001110100111000111011101101000000100011010101100110000011100010101111101110101001101011010101011111101011010101011111100000011111011111101101000010000100000;
#1 $display("%b", po);
# 1  pi=207'b000100111111000010111010011001100101110101000100001110111100011110101110111101010110010110011100010101001001010001000010010010000011000011011111110010010111101110000001110100110000010110011010101000000000011;
#1 $display("%b", po);
# 1  pi=207'b010011011011101011110001010001110110001100001011010001011001001100000011100100111011011000000001111011111011001011100110010000111000110011100110100000000001010010100010100010100010100100010101001110011001001;
#1 $display("%b", po);
# 1  pi=207'b001001111011100010110110001010011001100010001111010001100111110110100011110001110100101111101101010011100000011111001101101100111100111111110110101001011001101110100111100100110110110100100101010111010101110;
#1 $display("%b", po);
# 1  pi=207'b010101111011100101010110011011000011001111001110001111110011001101010010101101000010000110111001000100001111110100101100101110110011011101011000010011001101011100110110011001110011000100000111011110100110010;
#1 $display("%b", po);
# 1  pi=207'b111010011111011011100111000000101001001010011111010010111110110001001011011001111000100011011111001010011101000110110100000010111101010011111000111100010100011111111101111100010000001000011111010000100010100;
#1 $display("%b", po);
# 1  pi=207'b011000101101010001101010110111101011100100100001010010111101101001010010000100111100001101100100110011111001000111000001100011111010110011011101011000100000110010001101110011001100110011110011000001111010110;
#1 $display("%b", po);
# 1  pi=207'b111111100001001011010001010000010011000101011010010110010110001111110101110101010001011101111100001110001101101000111110100011010111100100000111000100010010110011100100110010101000001000001110111101110100011;
#1 $display("%b", po);
# 1  pi=207'b101010001001011000110110110011111100000011110000011010010000101001101000111110001100011111001011010110101100100011101101110100011101110111101001101110111001010100100001000001111111111100011011110011011000001;
#1 $display("%b", po);
# 1  pi=207'b000101001111010110111100111010010010010001010101101110011010110100000000100100001010000100001111011000000010000011010101110010100000100010011111100111111010000111110011101001010111111111110110011000101001011;
#1 $display("%b", po);
# 1  pi=207'b101011011111101000011100111101001110011010100100111011101110101111101100110011001000011101010111001101000100100101001100100011001011001100010110011111010011100011010010101001111111111101110001011110101010000;
#1 $display("%b", po);
# 1  pi=207'b000100000101010010101001100100010000111001000110010111000000111101011100011111110011011110111101011100010110001110010000100101110011011001000111011100111101110010101001001000001011110000011111010010011011000;
#1 $display("%b", po);
# 1  pi=207'b000111001000001001011000001101001111111001011000111001100110101101110100100111000101001100011100110110011111001011010010110011001001100110110111111101111110110111010100011010100011000010100001100011000001011;
#1 $display("%b", po);
# 1  pi=207'b110010001010000101111101001001100101001000001110110111110000111101000101100111000010100010000010101111110001101010011000000100000100101101100010000011100001110111000000101101111011001000111011101110111010111;
#1 $display("%b", po);
# 1  pi=207'b001000000010111000100000000111011110100100001110101111011110000110100011010100100111000101001111011001100101101011001111010010110000001100101011011001000000000010011011000100111101111111110101010101111111011;
#1 $display("%b", po);
# 1  pi=207'b101011011110011000011100011101011111001110110010111111011001000011111100111111101110101000010101010111110011000001010111100101111011000001101100010111010010101111001000000001001011010110001111011100101010001;
#1 $display("%b", po);
# 1  pi=207'b011110111100011011111001010110110011101010111110100101001001010011010010100110111101011111111011011100001110100010100011111100010010110010000001110000101011111111110111101000000100100110000111100000100011010;
#1 $display("%b", po);
# 1  pi=207'b111011001011101000000110000000111001111000000101110001011101011001010000010010001010100100000000000111101101101011001000100110010000100001010111001000110100000010010011010000100001000100001111100100100111001;
#1 $display("%b", po);
# 1  pi=207'b110011101001001110110100101001101000101011100011011101101111001000010110000100000011001011001011000011000010010001111101011001100111000010100101101000000110010111011111110110110011110011010010111010110010110;
#1 $display("%b", po);
# 1  pi=207'b001011010100011011111110000101111011011011001110010100010001011100001010001111000001111010110000010101011100000010111001001010100001010111000110110010001110100011001000011101111100110101001101111110000000010;
#1 $display("%b", po);
# 1  pi=207'b111010111010111010001000101110010110100011011111101011011001111001000010001011000101100011111111100011000101011100001101001010010101001011100000010110111010110001001010011000000110100000110110111010010000000;
#1 $display("%b", po);
# 1  pi=207'b100001001110000111100100000101000111111110001101011110010101010000100100010011111111010011100000001101100000001010111001001101011001011111001000100111111001001000100100101000010100010000011111011000100001000;
#1 $display("%b", po);
# 1  pi=207'b011100101010111110001110101111011100100011010011011111111111000110101100010101011000000111011001101001011011001011111011101100010010001001000001000001001001110110010110110010000011110010011110101011111000000;
#1 $display("%b", po);
# 1  pi=207'b010110110100001101000101010111110010110000101101111110111110111011111010010001000100001110100110110101111110000011011100101000100010011101001101100011101000111101101010010100111010011100010001011111010111111;
#1 $display("%b", po);
# 1  pi=207'b001101110111001101001100100101001010010101000111001110110111010101001101111011011001001101011110001011111111001011000000110110010110100110011110001110011101001001111100100100110110101101100100111111010110001;
#1 $display("%b", po);
# 1  pi=207'b100001010001001000000110111000010110001110101101111011110001011110001111100110001101011101111001001000100001000101100111100100001111001000101011111011110110010000011100001100100010001010100001000000010010111;
#1 $display("%b", po);
# 1  pi=207'b010100011000100111001011111010000010000010000011100101110100100000011001010100010101100001110101101111000010101010000010101111101101000111101110001010100010111111111111100010111111001110000110111101001010100;
#1 $display("%b", po);
# 1  pi=207'b000000010111001000110010111011010101101111110111111101111010000111001101010111010000001000101110011000101011000110101010110000000111101001111110000011001000100101010111111001001111110000100111101010111101011;
#1 $display("%b", po);
# 1  pi=207'b111111100111110010111100000110001111111111010010000000101110010011100000110111110010110001011110101010111111010010010010111011100110001010111000001110001110010001110010100110011000110110111010100001101001110;
#1 $display("%b", po);
# 1  pi=207'b101110000010000010100101000100000110011101110100110111101001111000111011101001001000010101011111000111111000011101000110010010001100010010011010001110010011001100011110110100101110001011100010100101011110100;
#1 $display("%b", po);
# 1  pi=207'b100111010100110101001111110011101000110111101000100000101100000101100101000010111011011110110001010001000110101110111001110111000101001001110101001101011110011010000110101000010011001111011010111101000101100;
#1 $display("%b", po);
# 1  pi=207'b111100011101100100111011100110010000011111010011000110101000010001101001001010000110110100111000010010010001101010101110001010000110101010001011001110001101100011100001000100100001101000011000000100111000101;
#1 $display("%b", po);
# 1  pi=207'b001111111100110111100101011111000110101101110101110001111101010000011010010001010100111000100101111011001100001100111110110111100100100110011010101011110110110111110111101111010111101010010000010100101101010;
#1 $display("%b", po);
# 1  pi=207'b100000100010110010111011101011100100110101011101110101000001101001011000001000111110111101101110010001110111000010111111101110010001001110111110100110001000110111110001001100010100011100110111011111111101110;
#1 $display("%b", po);
# 1  pi=207'b000101111001000110100011110010000110011000111010010111010110110001111000001100101001001101101010001000010110110110101001010100001000001011001111000101001000000110001000000010110010110110100001101111101001010;
#1 $display("%b", po);
# 1  pi=207'b010110101101111111100011001000001100001110100010001001100000001100000010011000111101001100001001100111001101100111111000010010010001001000011010101011011100100111001010011000010101010000101111010000000011101;
#1 $display("%b", po);
# 1  pi=207'b011011011010000000001110001001101011010101011000111101101000011101111110011010110101100000010100010001110000001011010010111101011110011010101000001011011001100000111101011101110101001111100011100100100100011;
#1 $display("%b", po);
# 1  pi=207'b100111011011111100001110011001000100111100111000111100011111001100011010101110100101010000100111011110010010110110001011100001010111111111100000110011111100011110000011011010011011000111110000010000111111010;
#1 $display("%b", po);
# 1  pi=207'b100100101111100010001100010111110111111000001001100000011001101010000100110010110000101010101000001000101000110010010101000101010010111000101100001110011010010101101101100000000000000111011101001010111000010;
#1 $display("%b", po);
# 1  pi=207'b101010101111111110100101000100010001001111100011000011010001011011001110110011000100000110101101111010111011101110001101010100001100011110101011011010111010000000111110010101101010100110000101110010101101111;
#1 $display("%b", po);
# 1  pi=207'b001000100010011100110000110110100001010111111010100000011000001001010110001100101011100000010110110110111001000111100101110011001010001111111111011000011001110000001101110110100100001100100000000101110110001;
#1 $display("%b", po);
# 1  pi=207'b100001000011010110010101001001111100101110000000010000110011011100110010100110001010100010001011100101010101101100011100101101111000101010100100010100110110110010101001110001010111110011101000100000101110101;
#1 $display("%b", po);
# 1  pi=207'b110010001100001110011000100111100000110100111101111011100110100010011010000100101010110100010100000100101000000101111011001110111110011001001011010110011100000111100100001101011111101100011100110011111100111;
#1 $display("%b", po);
# 1  pi=207'b010100001001011001110110101111110110101110000110000000011001101111011100101111100001011000110001101110011000010001111010101101000010011010111000010000000000111001001100001110110110100011100011110000101110000;
#1 $display("%b", po);
# 1  pi=207'b011011000000010011111010011110110110111010100001110011011010101001001010101101010000011001101011000000101101111010100011110111101001111101011000011111010011010000011110010001010101011011000010000011100110101;
#1 $display("%b", po);
# 1  pi=207'b110000000100111110011110010110000001011111000001100011010000100101100000000001000110101000000111101100110100001000001110101111000011010111100101101100110010111011000101110110001110111101111111000000001111111;
#1 $display("%b", po);
# 1  pi=207'b101101001111011100000110100110001011101111101111111001101010000111010111001010110011100110111110011001011010100111110110010001010010000101011010110010111101010110100100110000011111110010110101011111110111010;
#1 $display("%b", po);
# 1  pi=207'b101110010010101100111010100010011010100111000101000100000100001111110111010110011111001100111111101110010111000100000101001010110100000110010101000110010010101111101100100001110010111111101001100100011010110;
#1 $display("%b", po);
# 1  pi=207'b010000110101010000000010110011011001111110010011111010001011000101110110001001001110001100111000010110100001101110011101010011000101011000101110101000100100010111101101010100111101100101110011010101100101111;
#1 $display("%b", po);
# 1  pi=207'b111111010110000111000101110001100001110111001111001011000011001000011111001101110101110001100000011010111001001001001011001111011100101010111111101100000011101110110010110011101101111011101001100110101110001;
#1 $display("%b", po);
# 1  pi=207'b111101110011011110000010110111001110001011000110000100101110110000011010000111111011110110101101000100101011100000101000011101100111100001001110100100001111100110111011101111001011101110001110110000010000100;
#1 $display("%b", po);
# 1  pi=207'b111101101111110001010001011111011001111000110001010001111000100100100101011110100101010101011010100111111100111100110011001110010101001110101110001101001011001000001001001101011101011000110101110010110101110;
#1 $display("%b", po);
# 1  pi=207'b000011100101100011110010101000010111010000010100010011000011101101110010010111000101110110100010011110110101011100101101011010111111001100010101010100001110010011001010011010010011011000011100001001100001000;
#1 $display("%b", po);
# 1  pi=207'b100000001010111111000110111011001110100001111010011010001100111010100010111011110101101100101111111101000101000000101111100101101001010011101111000011001100001010000100110110011101111011000100110101001110101;
#1 $display("%b", po);
# 1  pi=207'b010001010100100101100011000101000001000100011010010010110011101001001000010110001001010010010100001110000101010011100001100110111111001011001011011011011100100111111011010010001110001110101100101000110100111;
#1 $display("%b", po);
# 1  pi=207'b011001110011011101110010101101100110111010110000001100001111100110101110110010111000001000100010111110001000010011001001100101101000111101110010011011101101100000110100010001101100010110100101100010000110100;
#1 $display("%b", po);
# 1  pi=207'b100011011000101101011101100000010101101110001100100101011010010111011000101011111011101000001100001000000101101011100010101000010010001110001000110101100100100011011101111111011010000110010000100110111010010;
#1 $display("%b", po);
# 1  pi=207'b001101111000111001000011011111100111000111100110100011010010011001101011100010011110001010010001111110010011010101001100111111001010101010100000010000111111011110110011111010000101100110110010111000000100001;
#1 $display("%b", po);
# 1  pi=207'b011001000101010101100011101101001101011001101000110000000010000001110001000101111101101011010111000111100010000100101001001111100010011001101001001111111101110010011111100100100110001000010100111000000010111;
#1 $display("%b", po);
# 1  pi=207'b010111010011011010111001110011001001010011011110010110000000100001111001011010011101100101001001111010010111111101011010010100110101011000010000100101100010011010011011010100111100010111011100011010111100111;
#1 $display("%b", po);
# 1  pi=207'b101001010100101010010111101100001000011111011001101000100100101101011100011000001101101000110100010101010011010010101010101100011000011111111101100010010111110000110101011100101011011011110011010111001011001;
#1 $display("%b", po);
# 1  pi=207'b100101111101010000001011101001110100001111000101100000000110100010000110001111100101111101100000001100010101001010110111000111011001010000110100001000110110100111100000100111010011000101100000010000100000001;
#1 $display("%b", po);
# 1  pi=207'b101111010101001100111110011101011010010001110111110000110110101011011001101011101011111000100010100110001101000011001000011100000010110111011010001111110111000101110101101000110010011111101010111100101001110;
#1 $display("%b", po);
# 1  pi=207'b001100000000110101010110111100101011010010101100010010111100000010001000100001001101000110110000111011010001110000010110011011011000010111111010100001100110110101001111000100001110110001000101001011111011111;
#1 $display("%b", po);
# 1  pi=207'b000011000111110101011011111111101101111011001000110000010010000001010110011111011000010011100111011001001011101101011000011100110100101001010000000101101001011101010001001011110011100100000011111110111101001;
#1 $display("%b", po);
# 1  pi=207'b000001011100101011110001010001001011000001010000100111110001111011100110101100100110110010011000001000010010000011100110100001010111110110000001001101111100011110010110001011101100110101010110100100001001000;
#1 $display("%b", po);
# 1  pi=207'b110001100101101001100010000000000110011000111001110000101011001111010100001100100101111101101010111111110001000010010000110001100010001010101110001101110100111100000111000000111000001101010000011111111100110;
#1 $display("%b", po);
# 1  pi=207'b111001001010000011100011001111001010011110100011000111001010011101110111110101101111111101100011100000010001100101001010110001110111101001001100000001111011110101101000010110011100001101110011111101110100001;
#1 $display("%b", po);
# 1  pi=207'b100101100101000000111000111100101101000110100110011001110011010010001011000011001010001110000010011110111110100001110011010101111000001000011100100011110010101001110110011000001101000010101101100010110010011;
#1 $display("%b", po);
# 1  pi=207'b011111100100100010001001001101001100111010001000010000101101111001000010110111000010110110001011110100110000100100000100010011010111110010111010010011000011010000000011011101011100001001011111001010000001011;
#1 $display("%b", po);
# 1  pi=207'b011010110111100101110110111110011101010010100101011101001011110110100110111101111100001110010011000010000010110011010011100001011110001111001000100011010010101010101011001111011000001110111110110001000101010;
#1 $display("%b", po);
# 1  pi=207'b100010100001101110111011111110111110101110111110111001010011010001001010101101100001001010011111110001100011100111101000111010000001110101011011011110101100110001000010000010101111000100110101100000010010101;
#1 $display("%b", po);
# 1  pi=207'b111001000100011110010100100111001110101001011011101001101010001100010011100010000001111011100100000101110111011010000000010111101110001000000001010100001100111100010101100111011100101000001011101111010000001;
#1 $display("%b", po);
# 1  pi=207'b010100001101011000011011111100000000001010011010111111100011101000101101110001001111111011110001000010100111110001001110100101100011111011001001110101001111001101110100001111001100110001100110100011101001011;
#1 $display("%b", po);
# 1  pi=207'b100000010011000100111011011111101110011011000001000010100001101011000111101110011101000100110000000100111111111100101011011010101001001111101111010000101100011100001110001011110101101011001100001011100101110;
#1 $display("%b", po);
# 1  pi=207'b001111011100110111000111011111000101010001001100001110100101001010101001010010110001101011101010101010110100111110101110001001000000110111001111011110001100100100111010000101000101001101111100000110001100011;
#1 $display("%b", po);
# 1  pi=207'b011011001011010111011110011100100000111101011011100101100001100011001010100101001110111001011000010100100100101000000011100011110100111111100101011111111111011101011100000110110010010101000010111100101110101;
#1 $display("%b", po);
# 1  pi=207'b010101000110111100100000101000111010010100100101000011100000111110000101110110111000010111110010010111010101100000111001001100001011101000111010111001110111001101110101000010111010011101000000010011001000000;
#1 $display("%b", po);
# 1  pi=207'b010101011010001100011010011111101111111010000010110001111011101010110010010011111011000111000111101110101010010110000100001011101001010010000111011010010110110011111001011000010010010101001110110010010110110;
#1 $display("%b", po);
# 1  pi=207'b111011111110001010111000000010101110100010100011011001010100011101010100100000100101110011001000011100010100100110000001001000001101011111000101011010111000000010011001000110010111110001011111011101110000111;
#1 $display("%b", po);
# 1  pi=207'b000101001100000111100011000110010000101001100111010000011000001100110011001001101011011100001010100001111110010001000011101101000111000010010001011101010001110011010101111001011011000001111110010010111110110;
#1 $display("%b", po);
# 1  pi=207'b111101001011001001111101011011001100100101010010000010010110100011001111010110101000011100110100101000010110010000101000111110011110110001011110100011110111010011101110010110010111111010101110001110100001011;
#1 $display("%b", po);
# 1  pi=207'b011111100110011000001100000001110110111000000110110101110010001111100101111011001111110001000101101000000001000011111011101001001001010010011000100110110111101110110000010111010000100110110100100011010101101;
#1 $display("%b", po);
# 1  pi=207'b101101011101011010111100100100101111001100110011111000110011001111100011110010101000011011001111011001111100001000010000011101001101000010011001011001001100110010101000011010001110000000010101011001010100111;
#1 $display("%b", po);
# 1  pi=207'b011111000100100001100110011111010110011000001000100100011011000101110010111110001010011110101011001111111001011101011110000000111101100101001111111000101100111100010011101100001011111001000001011001101101101;
#1 $display("%b", po);
# 1  pi=207'b000011010010001011100000101011011010011101010011011010000101110100001101100011011011111011100110001101000111011101000011011010101001011101010110000010001110111100001010011001010100000111010001010000101111001;
#1 $display("%b", po);
# 1  pi=207'b100101001000001110011000110100001010101110011010111110101000011100111111111000111111111110111000010111100110100011100000000010010111100011110101001100010111000101011110000101110111010011001101000000001000110;
#1 $display("%b", po);
# 1  pi=207'b010011001100101101110101001111000100110100101000000100111001001010110011000000010100111100001110000000001010110111010000100111001000000001001100100011011000110000101011011011111101000100100001100011111001010;
#1 $display("%b", po);
# 1  pi=207'b001101111001001001001100000100001010100000101011101001011110101110001001110001101011001100011101110111000100101100100100111110000100101011111111011100110101011110010000001101100000111101011001110001000000011;
#1 $display("%b", po);
# 1  pi=207'b100110100110101011110100110011000001001000111010000000010101101101011011111100100010100101010000100100001010100110110100101100110111111011001010001110111100111000001011011010110010000010000100111000101111000;
#1 $display("%b", po);
# 1  pi=207'b000111100100011100000000100110110000011101100111111101111001111101111011000101100111010001111100000001000111000110111100000000110010011001100101111110110010110010100101101001011111101000110011011010010101110;
#1 $display("%b", po);
# 1  pi=207'b011100010001000000011000101010110110110010001000110111011110100001110000111100001010011000110100010011011001111100111101010010000011011000000010111010110100001101001010011010000101101010111100110011110010101;
#1 $display("%b", po);
# 1  pi=207'b010111010110111100111101010110001111111100110010100111101000001011100111010010110001100011111111011100011100100111000101001010110110111111110101000000010000000101011011001100101110100000011001101110001001111;
#1 $display("%b", po);
# 1  pi=207'b110100010110010100011110011010010010101001101010101110000100000010111000111110101111001011110010101111111010100011111100000100010000010101111010010010001010011010010001100001101011001110010011000000001010101;
#1 $display("%b", po);
# 1  pi=207'b110000110000010101001000001100111010000011000110011010011100000011001111110110111010100010001010001100111011100110010010001001110010010001101011110100110110000101100111101100101010000011110110010111010110100;
#1 $display("%b", po);
# 1  pi=207'b100000100100000101101011100000011011110100011110100001101001000011011011010000000111010100011110011111100001100111001011010110001110111110000000111100011000000110011011100111101100001101001011111110000001011;
#1 $display("%b", po);
# 1  pi=207'b101011000010111111011001100111101100001010111110110111110010000001000001011100100100111000111011011100010000001101100000101101000000000011000001000000001100011000100100100010000011010100100101100010011000001;
#1 $display("%b", po);
# 1  pi=207'b001010101001000110100101011010100010000011101011011001001010000001010110101111111100001011000000111100100110110111000011111010000110110000101000000110111111111000001110111101011101000000011010001000111101001;
#1 $display("%b", po);
# 1  pi=207'b111001100111100111011010011010001010001101110101101111100101001010100001000110101000101000010011001000110111001100001111100110010000111100110111010011101100110101000101001010110000100011100100001101010010011;
#1 $display("%b", po);
# 1  pi=207'b101001001010000010100101000001111101000000111001110000001100010011011001011011111011110111001111110010111100111101110110101010011010001011000111011010011011000110001101000010101010010001110110110010010101101;
#1 $display("%b", po);
# 1  pi=207'b100111101111101100101011101100110101101011001110111100000010001110111011000010111110101110100000011101100011111001010100100010101110111111011000101000111011101111010011001110011001111101010001010111000001111;
#1 $display("%b", po);
# 1  pi=207'b101111001001011101000111101100011100111011110010101000100101011111101110011001010111100000111111101110001100000011101000010110011001000111100100110110000011000001111000010000100001000011111010101010010000011;
#1 $display("%b", po);
# 1  pi=207'b110111100001101010100010001101100110000111100001111000111110000101000111101101101000001001110010001100101101001011010011010101100110001101111110010001101111110100100010111011011011110111011011001001111100001;
#1 $display("%b", po);
# 1  pi=207'b101101101011001000100010110011010011111001100000011100011101101010100100100000111110100110100010111001110001001000000001010011111101001010100100100110100110010110110110001000010011001010011000101100010000001;
#1 $display("%b", po);
# 1  pi=207'b110000100100101001110010100010100110011000111100111111011100100010101010110111101110011000011001101001010010100011001010000000111011000110110010100010100101111101101100010111000011011111000100001101100000001;
#1 $display("%b", po);
# 1  pi=207'b101000110111101010111010110000101010111110000010100100111111001010101001110010000100000010010010101001100100100110100011000100001011100011101011110001000011111000111111111001101011110000001010111000110000100;
#1 $display("%b", po);
# 1  pi=207'b011110010111100001111000001001110101111010001000100011011111110001111101100110001010110000110001100101011110101000000111101000001100010100110001000111001011011001100101001011010111001011000010011010100010011;
#1 $display("%b", po);
# 1  pi=207'b000101010110001110110010111101000001100101101110001011001111011110100011110000111101111111110011111111101010111011010111011000110010101100010000011110111001000100100001100010101101110001011110001110011000011;
#1 $display("%b", po);
# 1  pi=207'b000010100111011111111110011100011111010101110100001011101010010010000001101111101111001001111100000001011010010101111100111011101110110010001100010111101011000110100111110000110100010000001010010101001011110;
#1 $display("%b", po);
# 1  pi=207'b001000001110000100010000011011000001101001011110000110011000100000010101101000110001011010001000101010111000100111111011110000110010001111011100100100010110101110000000110000111110111000011000011010000000001;
#1 $display("%b", po);
# 1  pi=207'b111010010000000101110001000100111011111010001001010010111010001110110000111110111001010001011110000000101100110011111100100001001110100101000001101011111000000010101101111110100111111111101110100101010011011;
#1 $display("%b", po);
# 1  pi=207'b010001111100000110110100011010001000000010010101100011000010110001000000000100111100101110100101011011010011011011110011011000000001111110100101111101001111011000010101100011101101110100101011110001001101000;
#1 $display("%b", po);
# 1  pi=207'b100011010011101110101000010011111000011001111110111001011011110001100010001110000011011000101100111010110101110100001110001101000111110010001001101110010100001100110101011100100111100101011011011001100101100;
#1 $display("%b", po);
# 1  pi=207'b100011110101100110111101111100100011101010001000101001001010100010101110001000000000111110011100001101101000010000000101111110001000110011011111001110000000010001111010110000101000010001001111001010110010100;
#1 $display("%b", po);
# 1  pi=207'b110100101111101110110000000001000000101010100011111110011100011101100100110110010101001100001001101001111101111100111110110111100001111000001001000100011111001010111011001000011111111000111111010011001010111;
#1 $display("%b", po);
# 1  pi=207'b101011110111110001100100011111000001100011001111100001000101010001001100111010010110100011000100101110110101010100000010011100111100110011110110011000101101011110000111011010101011000100011001100110110111101;
#1 $display("%b", po);
# 1  pi=207'b001111000010110110000001100110011110111011000011111000101111101001001101111110111000010100001010110010111011001111011010000100100100111011000010100000101100111001011001101011011001110110100000111010110000011;
#1 $display("%b", po);
# 1  pi=207'b001101111011011010010111111100010000000000011001000101101100111001110100001110111010001100001111010000001111001110111100100110000011011100011100101110110100100001000100100001011110010001101010011110011100011;
#1 $display("%b", po);
# 1  pi=207'b110110100000110010001111010010010011000011111001100010000110011011101111100010111100010011100000011001001100111100010000110010011010110000110101000010111101011001001111100001101110011010001101110100100101101;
#1 $display("%b", po);
# 1  pi=207'b110111011000001110100010101011000000011111110111111110100110011111111011101110111111011110011001000010101101011100101000001110110011100100100111110110001000010101001100110001110110100101000010011100000011110;
#1 $display("%b", po);
# 1  pi=207'b000100110001000111100000110001110111100011111001000100111110011001000011101100110001001000111111000110101110111100111111001101111001011111111110010001101000011111011011101100111001001110000100011111111011011;
#1 $display("%b", po);
# 1  pi=207'b011011111000011111111001001100001010010011000100100010011011111010111010011111010111011111100110110111110010011100000101110100001000111101000011010110010101101011010001111101000010101100100111010100100000001;
#1 $display("%b", po);
# 1  pi=207'b001010001110101010111000001001101101110001011111111010111101100000010110011111000000100011111000011110010001111011011100010011001111000011000100001001001000011001100100101100011101111010011100101000010111000;
#1 $display("%b", po);
# 1  pi=207'b001010000111100111100011100110000110011111010110000111101101011100111011001000100000001001000101100100000001000011011101000010010110111000010101100011101101100101100100111000000010001011010110111101101001111;
#1 $display("%b", po);
# 1  pi=207'b110111100011111100000001101000101101010100011101100110001010001110100010011011111011011010011010010111011001110100100001010001001110100110010010110000110101000111100110111100010111000111010011001100000100110;
#1 $display("%b", po);
# 1  pi=207'b011101011101011001000101000000100001101001011010101000011110010011001001011111010010001110101000001000000110000000010001000001101001110110111000100011000011101110000010110100000010011110110000100111100111100;
#1 $display("%b", po);
# 1  pi=207'b100110110001100000101000111101101011001001100111001010001111100010010000101011111010010001000110010001000101101011110110001011111011001011001001001010101010100011100000111110010000010111000010000011100001010;
#1 $display("%b", po);
# 1  pi=207'b011001001010010110000110001001000000100110111101111001110010010000100100011010101110100010011100100100111001010101000111011110110010001011101000000110111010110110000100111101101001001011011110000011111101101;
#1 $display("%b", po);
# 1  pi=207'b011001001111010100011011110011011110011111000001011110110001101011110110101111010010101011110110010010001011010111100011011011111100101101001101101010110111010110111000110011111111000111000011111100010011000;
#1 $display("%b", po);
# 1  pi=207'b101010000010000101111110101110010010111101111000111110010111000111111010000000010011101011111100001000000111111101101011001010110100010000000000101000101101111000100001000001001110001101011000101111011000001;
#1 $display("%b", po);
# 1  pi=207'b110101111110101001010110001100001101111001001111110001011011111100010101110010000110111101001011010100010001001011100101010000111101001000000010111000010111101111010011001010101110010110000010111001011000000;
#1 $display("%b", po);
# 1  pi=207'b110111000010001110111100000011010010100010111110100001101101000111110000001011010001011000010101101110001001111100000010111100101010101001011101001101101100111111010011011101110010111100100100010110111101100;
#1 $display("%b", po);
# 1  pi=207'b010100101100010011000010000110110011010111100001110110000011000001110111111011100110100100111110000011110011110000010001110111101100010110101111101111010100101110110001000101000000011101101101101100111101101;
#1 $display("%b", po);
# 1  pi=207'b111000100100100111111010100001010010110110100011111111111101101001001110110101011000101100001011111001100001111111010001001010000100001010010010000111000011000001010100010100001101101010001100100101110111111;
#1 $display("%b", po);
# 1  pi=207'b001110100000110101111011000110000111010100000110011111101101011001110101100100111111000101010011000101101101000011111100101111110010001100101101100110000111001100101011001111010111000010100111101001001110111;
#1 $display("%b", po);
# 1  pi=207'b100000011111100111101000111110110100110001010010001111111001101100110001100110010100000110000010001111111010100111110110111111011111100000110000001000010011011000100111011000100000010100101111001010011111011;
#1 $display("%b", po);
# 1  pi=207'b010011111001100111010001000101101100111000000111111111111001000111010101100101100011101111110001110011110011010111100110010011101101110110001010111111100101111101100101000110110110011100111101011100111000101;
#1 $display("%b", po);
# 1  pi=207'b100001000000111100010101001101101010001101111000000101010010110101010011110110010111001001101000000100011111101110011101010010100001111110100001100000011010100101011011101100000010010001111100011111001111000;
#1 $display("%b", po);
# 1  pi=207'b100010000000011000101010001011110001011101110001111000010000100111111001101010011100111000110010101010101000100001111001100111010010001100011000010011111110100000111011001011110010111011011010001011011100010;
#1 $display("%b", po);
# 1  pi=207'b100010100100101101011101000001000011001101000111100100010011110001101100010000001001101010101111101001011100000110011101100011000100000110011110011010001011000010010010110000010111110100111000010101101110110;
#1 $display("%b", po);
# 1  pi=207'b111100011110010110101100101001100110010100011000110110110000000011110110001111011000110010100111011101101110101011011001000111110101001010001001110001110001000010001100000110111010110110101001010000111111110;
#1 $display("%b", po);
# 1  pi=207'b101000010000010110110000010000010000100001110101100010111010100111111000011110000111101000101001101000100010010101101011000000011110100000001101110000110101110001000110110111100111010011100011110101010001010;
#1 $display("%b", po);
# 1  pi=207'b110000111111010100110001111001000010111111111001110010000011011101110010001111000110100001000001101111000000000110110101101010011000001001111001001000101101110010110110111001100101001101100100101011011101101;
#1 $display("%b", po);
# 1  pi=207'b011011001110000110011000001010010001111010011110010000111101111001010011010010000001101010110001011010010010110111000011001100000101100110110010011111011000100000011101100110011011000111010000101110011110110;
#1 $display("%b", po);
# 1  pi=207'b000111010110100101001000001111011011101001010000001000001111001000000111010111001011100101011001010000010101111011000000110100001001000101000001001110100100000101000010110101011011000000110010101011010111010;
#1 $display("%b", po);
# 1  pi=207'b101000010011010001101010110001001110000011011110000010000000001111001000001110110001101100000001100110100110110001010100101101001100101011000000101011010000001001101001000100011001001010110010001111101000101;
#1 $display("%b", po);
# 1  pi=207'b011001101001111110001100111100001011010100001011101101010011100101011000000011010001110000100101110101000100000111101100001110100010100110111001110111011010101010001101101000111110011011101101101101010111000;
#1 $display("%b", po);
# 1  pi=207'b101010101111111100000101110111100101101001101110010000010001000001000100010110010011101110011011000001110010101100010111011001101110100111010000000000101001010000011111011000011001101101000010011101110011111;
#1 $display("%b", po);
# 1  pi=207'b010100110100000001011110000110001100101101111000111110001001011010011111101100110001110001100101101110011110001011110100010110000011101000110111010110110100100101000010000111011110010100110001111010010100101;
#1 $display("%b", po);
# 1  pi=207'b110110011000111001000110000001000100110011111110001100100100111010001101111010101111101100011101001011111001000010100001110111001111001110100111111111011000010110111101111101110001011101110101001011110010001;
#1 $display("%b", po);
# 1  pi=207'b011101101111111001010110101010010000011101101110001001011110101101110011010111101110101000010010100010010100000000001111001101000000011101001000100101111100101000101110111110011000001011100100110000101010000;
#1 $display("%b", po);
# 1  pi=207'b010100100011111110110110110111111110001010101100001110010000110110111101001101110101111001100011101110110010101101111011100010110110000001111110011101110111110100001100010100001101010101100111000001011100001;
#1 $display("%b", po);
# 1  pi=207'b000110101111100101011010011010100101110100011110001101111011111000011000100000111110001010101100000101000100101101001100011001100000100010010011100001011101110010000001100110110001110101110101111100010010010;
#1 $display("%b", po);
# 1  pi=207'b000001011001100101110010100111100001101000100111001001011010111001100011101111100110010100111000111100111010001101110011111110100000001010001100001110101000111111101100001010110010100110111000100100110010000;
#1 $display("%b", po);
# 1  pi=207'b010001000000011001110000101010101100110001011010000010011111011011000000111110001101100110001100011111001001011110111101010000010100101101000001011010101010110100010011011001110111011010100111100001110011001;
#1 $display("%b", po);
# 1  pi=207'b000010010100000001010000010001001010101111000110111110111010110010011001011010000010000000010001110000011110100000101010101011010101011010001000110110011011110011011110011100111000011110000110111001101000100;
#1 $display("%b", po);
# 1  pi=207'b011110100100010111010011001110011000110001011110101110011110000010011101001100111001001010000000100000100101100010000000110111011111101001101111010010110110110010101110010001001110101000110011000000101111010;
#1 $display("%b", po);
# 1  pi=207'b001100100100010111010000000011001001101000101101111011010100011000011010001110100010100011000000010010010101000110011111111111000000010011011100011010110001100111001001111100100111010110011101010011110000000;
#1 $display("%b", po);
# 1  pi=207'b011011100110110110000011111010011100110101100010001010000100110001000000010001001100011111110110100011100111000001010100001101101000000000000010011000101010100101111011101010001111011110100000111000001011010;
#1 $display("%b", po);
# 1  pi=207'b000010000001101100110010001111001001101000111110101100010111101101000101011100010010001010000000100100110010011010001110110101110101010011111000110110100010111101110101111010110101100000011000001011010100100;
#1 $display("%b", po);
# 1  pi=207'b000111000001101101000101000000111100101111110101011110111010011101001101011111110111000001001010000110100000000011010111010001101001111001111101111111111000001100111111010010101111100010100010101011011101011;
#1 $display("%b", po);
# 1  pi=207'b110110100101010101110000010010110101111000011111000001000010110110101000101001001000110110000101101001101110100000010011111000101011101000111110001100010100001011001110100010110110101010000110111110011010100;
#1 $display("%b", po);
# 1  pi=207'b000011100101001110011111100110000000000100000111011001111000101110110111000111110101101110110111111101001111010101010100111100011011110010010001001101001100000000101010101111000010001001011100011010100010101;
#1 $display("%b", po);
# 1  pi=207'b101010110011011010100101101000011011010001010001010000011001001110010000010010000010110111110101111110101101110011011100100100110110111101101101010000001010111011110000101011111111111101010100000100000001101;
#1 $display("%b", po);
# 1  pi=207'b001100010100010110101111111000001000111101101101110110100001011111001101011100111010010100010100110000101001010001001001001101101101000111010110011100100110001010010100101011001010110111001101101101101011000;
#1 $display("%b", po);
# 1  pi=207'b110101110111000110001000101010011010001110100110011000010010110011011010101100110110111101011001101101111101100100101111101010110011111101011000110111110010010000011001111110000011100011110101010011101111101;
#1 $display("%b", po);
# 1  pi=207'b001001001101011011100101001111011110011000010000010110010100100000110100010000001101000101011001110011010010100011010101100101001010011110110001011000111001011001101011010100100010100101110101110101110110001;
#1 $display("%b", po);
# 1  pi=207'b001110011001101100101001101111101100010111100011111001100100010100000100010010110011111001001110000000000111111001011100111001110010000010001110101011110001010100011001101110011010111101001110101110110001000;
#1 $display("%b", po);
# 1  pi=207'b011000100001101110100000100000111111011000100001001001011101011011111000100001001111110101011110000111100011111101111011001101010111111101110100011101100011111001010100000100111111100010100000110001010101011;
#1 $display("%b", po);
# 1  pi=207'b111011011011001110111010101000011101101110011110110111001111000001101000010011010001110011001000001001001000001011001010101010101011101111111111111111010100011101010011101110010010101011000100101110001111000;
#1 $display("%b", po);
# 1  pi=207'b010100010000110011111111111011010110000010111010000001000001111000101001110111111101000010101001110110110110010001101110100001101000010110010001111100010101001011010000001101001000100001110011010101000101011;
#1 $display("%b", po);
# 1  pi=207'b010101111001101010011100011100000111010110110100011010100101000110011110011100010100000010101000110001001011001000111011100100101110011101000011111000101110110000010100001010010101101010100001011001111100011;
#1 $display("%b", po);
# 1  pi=207'b111011010110110101110111110110110101010110111111100110011001010111110110101101111000000110111011001101110111101000010111001110101010001001100011000001110001100100101101000000000010001110000101001001011100000;
#1 $display("%b", po);
# 1  pi=207'b100101110011101000101001111110001011110001100001110110111000011100001000111000011011011110101010000001101010110010101000110100101111101101000000100000100000001110110010110001110000100101110110111001101000010;
#1 $display("%b", po);
# 1  pi=207'b100100001001100101110100000110101010101110001110010001110110110011100010000101100111110000010011001100010010011001011001111000100110101010100100011101101111110100111100010100001100100100000011100110011111100;
#1 $display("%b", po);
# 1  pi=207'b100011101100011011000110010111010000010110100010011000000001101011111010011100001111010001110001000111111010111100101011000111010101110100101000010111011101010010111110110000100001101011000100011010000100001;
#1 $display("%b", po);
# 1  pi=207'b110111110101011110011010111110101011111110100111110000000110101011001101000110110100100001100001110000101001100100111100000010101001001110101011010000111110110000011110011101011010101000110001001001111101100;
#1 $display("%b", po);
# 1  pi=207'b010000000000100101010001101111010000000110110010111110101011111011111110101110110100101000110000111001111011011110010110010010011011110011101100111110000110111101100101110101000000110010000110011101010010101;
#1 $display("%b", po);
# 1  pi=207'b001100001100101100110011100100000010110010100001111011111101001000111111110001100000001100110010000100110100110001011101100101110000000100101001110101110111010100000100001101000111110010110101101101101001010;
#1 $display("%b", po);
# 1  pi=207'b110011010110101101010110110010010010001000000000101111000100011110111101001111001100111111011000101000001000011001110100011010100001110010000000111101101110110000000000111001111001000001011101110011100111001;
#1 $display("%b", po);
# 1  pi=207'b101111100101000010110001100001010110111110011000111001110011010001110001110110110010000111011100100101101001111101100111011001001011000011000101100010000110110111111010110100000100111000100001001101101100111;
#1 $display("%b", po);
# 1  pi=207'b010001010001001000111000110010000100001100100110010111100000100110000110010001111001110011100110010011011011111101011001000100001000011000001000110001101100100111001101010111000111000110010101111000111001101;
#1 $display("%b", po);
# 1  pi=207'b000011100101110010110010100111100001100001101010101010010100001101010001011010110101011100011110010101100001111110000100001001011000101010100101010111001101111011011101000110101110111110011100001101011100001;
#1 $display("%b", po);
# 1  pi=207'b010011100101111001110110010111100011101110110111011111110000100111110111101110100111011010110011111101100111000001111111100100010001011001011011101000010101100101101001011001000011100010111011000000000011000;
#1 $display("%b", po);
# 1  pi=207'b010011110100000111101111111000111011001000110010011010100001110111010110111011100110100111100111100010101101010010110111100101011100100001010011010100110011101000100111000001001000111101010100011101010001000;
#1 $display("%b", po);
# 1  pi=207'b000100001110110110011001100111100100100101100001000111001011100010110101000000010100111000100101000001001001111011010110011110000111110101010011100011110010001111110011111100011111111111100010011100000100111;
#1 $display("%b", po);
# 1  pi=207'b010111110100100110011101001101000000010001100011100111110110001011111011111011000100101000111110111100101100110011100010000110101000101000110010100000001111000011010010101110010101100011110100010010100000010;
#1 $display("%b", po);
# 1  pi=207'b000010101110000010101111101000101101100000101101001100001010010101001110100100000001011001101010010000111100010110010011000110010011001110011011011111100100101110101011111001110110010101101101001001001011110;
#1 $display("%b", po);
# 1  pi=207'b000010000110101000010100100010101011100001011011001110110011011110010001000100101010011000001101110011001010100101011110011001010110010011000001101100111010001000100011101101011001011110110001011101011000001;
#1 $display("%b", po);
# 1  pi=207'b001101010001000110110111110010010110110011000010010110011010110111010001111110100011000100011000111101000111110111001101011010100110101100001101110110111100001110111001100101010011011100000101111101101101101;
#1 $display("%b", po);
# 1  pi=207'b100010101110101100101111011100100001010100110010111001011011100001100000111011010000000011111100100001000111100111111011100100100001110000101110000110011010101011001101011100111001110001000110101110001111001;
#1 $display("%b", po);
# 1  pi=207'b001010001110011010100011110100101001011010010111011111110000111101101101111011100011001111111010000000011100101000101110001100010011010000000110010100010101110010100001101000011000010000110010100101010010010;
#1 $display("%b", po);
# 1  pi=207'b000011100100011111111101110001100101110011001001010010010011000000100010100000110011010110110100111011100011010000100110001001011000110101101100010101100110110001011110000001100101110011111001101111101001011;
#1 $display("%b", po);
# 1  pi=207'b011101010001011000110101001000011101110001011010100011110010110111100101000001101010101010000010101000100100101110001101100011010010001011010001101001111001001100111011101000010001011100001000011011001000101;
#1 $display("%b", po);
# 1  pi=207'b110101000011011011001101111010001100001101110011111110110001001111001100110001100011101011001101000010001111000000110110101000101000111000101010001010100011001011010011000000111100100011110011001000100100011;
#1 $display("%b", po);
# 1  pi=207'b001100101111111001101000100111110001000111011101101100100011110010100000001110100100100101010000010111001111001011110010110000111011001101010000100010011001110101000101100001111010000110101110111000010110101;
#1 $display("%b", po);
# 1  pi=207'b001000011101010010001111001110010000110000101111111101011000110100110101100010110111110110011110000110101001010110110111010110000001111111111001001011110000101011001011111010111111100001010000111100101011110;
#1 $display("%b", po);
# 1  pi=207'b011100001001100101111001110011000000100001000001000100010010100000000001001111111110100111111011101001010111101000001100101111000101101111000101111010111110111111011011110001010101010101010001001110111100101;
#1 $display("%b", po);
# 1  pi=207'b111111010010110000100111101101101001010011110111000010000101010110001000110000101000111100001010010001100010010111001010100110101011100001000100000100001011111111010110111001010101001010110011000001011111110;
#1 $display("%b", po);
# 1  pi=207'b100001110110000000110011011110101010101010010100011000011101100001000100101010010011010110011100101100011110000010111110111010011100010101111010011100011101011100101010100011000111111010111011010001110011000;
#1 $display("%b", po);
# 1  pi=207'b011000111001010100110100110100011100111101010101001001001101011010010011000111000110110010001011000001010101110111001111000011010101011100100010010011001100101001000101001101001000001101000011010000011111010;
#1 $display("%b", po);
# 1  pi=207'b110111101010100101000100001110110100110010011110110011101110011000010011001111011111010101110110100111110101000111011101100011100000101011010011010110101001001001111101100010001011110010011111010000101000101;
#1 $display("%b", po);
# 1  pi=207'b000010000110000001000111100000111000001011110001110000001001101110011110100010110101011110110110111000001101100000110011010000101111100101111101111100111100000001011101111011100011111001111111001101101011000;
#1 $display("%b", po);
# 1  pi=207'b100010010100100001000111011100100001010001010100101011101001011100001011100001111100101010110100110011010011010011011100010101110100100100101101100011100011011101010000001111110101111111110110001000111010000;
#1 $display("%b", po);
# 1  pi=207'b101011100101011110011010110000110100011100100001101000100010010001001110100001110001101000011100111001110101010100011111010010101010010010010101001011010001111100000001000101110111100001011110101100110001010;
#1 $display("%b", po);
# 1  pi=207'b001001111111100011101100011110111101011001110111010100100111110001101111110011010001011000110100100011000110011001100000111111010001110001010000100011101100101000110001001111001000010101011101011001110111110;
#1 $display("%b", po);
# 1  pi=207'b000111010001000111110000101100110111011010100100011010111010010011110110110101011100100000001100111111010011000101110000001001100101001000101011111011011111110110110100010011101011100110110100001101010000000;
#1 $display("%b", po);
# 1  pi=207'b001001101110101011100100011010001010110011001000111110110001001110111011011010110011110100110010000000100111111000001110100000000011110010110101010011010110000011111001011001000011111000100101011101010001100;
#1 $display("%b", po);
# 1  pi=207'b110100110100011110000011110111100000101010110000010101001101011011101010000101010101010000001001000111111000100110111001100011111010100111010010100010000010111001011000111010100000110101001010110101100011000;
#1 $display("%b", po);
# 1  pi=207'b001101110011001000101111111010100110000101101111111111111110111100011111001001110100101000011000011101010100110001011000110101110001010110000001011100000110111010000001111010101011000001000101000110111000111;
#1 $display("%b", po);
# 1  pi=207'b011000101001001010010010001101001110100111011010011100101001000100111101001111111011010101100010010010100000111011111101011111011111011001010010011001110001101011110000011000111011101010010010011101100000011;
#1 $display("%b", po);
# 1  pi=207'b011011111001010011001100101010010101010001100111010101100101110001011001011100100100010011001010101000101111000000100101101000010010110111011100111010001101011100110011011111111111001001110111000110001101100;
#1 $display("%b", po);
# 1  pi=207'b110100000101100010011111100100110001100011010110111100001001010100011100011100100011111111110111101001011100010010001000010101101000001011010010110101100000101011010100011110100000110101011100000010110000010;
#1 $display("%b", po);
# 1  pi=207'b010111100110110110101010010010010111111100010010011101010001111001001000010000110000111001000111110001100101011110100101100001010100100100111101111011001101110101100100110001101110001110110000110001111101011;
#1 $display("%b", po);
# 1  pi=207'b100111011111011011101101110111111111111100010010011110111010110111011100000111110100111000100000100000101001010010111000110110011010100000000101101001111110001001101101100101111011101001101101011110110010001;
#1 $display("%b", po);
# 1  pi=207'b101010000001011111100000010001010111101110110001111011010010001110000111100010000110000011000100011000101101010000100010000001010001101100000000001101010101100100100100101001101011101001111011000000011011001;
#1 $display("%b", po);
# 1  pi=207'b010000111000100101101100100001111100000001011010111110111000011111010001000000001001010110000101001000010010111001100001001010001101111101101110110111010110101110100001100110010011010110010011101001101101000;
#1 $display("%b", po);
# 1  pi=207'b100100100001101010100010000011010110000011100110000011011110010100011001110101110001110011111101010101011101101101110001011111111100000100101111101100011111001001010011001000011100010110100010111011100110110;
#1 $display("%b", po);
# 1  pi=207'b110111001111010001110101111111110000101010000101111101110011010011111000010110000000100001001101011100111000101110111001111011111101001100011111111000101100010000001110100101101111011100100100100111000111000;
#1 $display("%b", po);
# 1  pi=207'b010011010010111010101000000100110100001101001111001000100101110110100011101000101101111010001000111011110100111000111101010000100000010111111000100001010101101000000011110011101101010011110110111001100000001;
#1 $display("%b", po);
# 1  pi=207'b101111101000001000001000011110110100110010111111001011101101011000001110000001011101110011011110011010101011100110010100000111000100111000101101101111101010000010010111000101011001100001100111000010101101010;
#1 $display("%b", po);
# 1  pi=207'b010010011000001010100000000010101001010011000100101101000001000010111111011010001010001111000110101111001101110100010001000000001111011110110001000000100000010000101010111111001101000100001111011100010010010;
#1 $display("%b", po);
# 1  pi=207'b110100010100000101100000110100100000000010110000110011000011100010011011110000110100101100011100110010010000001010000001000000111010000001100100001101111001110101101111001101000001100100001001111001101101111;
#1 $display("%b", po);
# 1  pi=207'b101110010111000110001001110110110110110100100100010010100010110010010011010100111001101010101001101011110001101011010010101011001000111010111010110001001010010101110101110100101011101001111001100110100010100;
#1 $display("%b", po);
# 1  pi=207'b000011001010111100000000000111010101101000111101000011100011100111000001111111000101101100001000110111111000110100100100100100010011100100100011001110001111100100001101001101000111011101011011011111100101000;
#1 $display("%b", po);
# 1  pi=207'b001001011000000101010000101000000100011010100101011111100010011101100000100110010000010100110011010101000100001011011000111110001101101101100100100001011100000000000111101000010000101111000001001001111111000;
#1 $display("%b", po);
# 1  pi=207'b101010100100101011101110110101100100011101111001000010100100101111101011111101101001010001011000100111111100111001100110010001100001101010111111100011010010101001101100100001110101111100000100001010110001101;
#1 $display("%b", po);
# 1  pi=207'b011101011000111100111101010100110010100111101011111000010001011010100100100101010111101000111000000101111111010100010000011011010111101110010111011100101010111111110010100010011111000000110000100010111010100;
#1 $display("%b", po);
# 1  pi=207'b111010010111101101010001010100011000111011010110011110011010101110100111111110000110101100011001101110001001111110110001000111101101001100011100111001100100101101001001000010001101000000010101011010001100100;
#1 $display("%b", po);
# 1  pi=207'b111010100001110011101010111011100101000111111001011100000110110110000100000100101111000000101110100010011010110001001111011101001001101100110101010100100010101101011111011000110000110010110011001010010010100;
#1 $display("%b", po);
# 1  pi=207'b011100100110100001001001011000000001111100100110101111011000010111110001101000011000100111100000100011001010001100001110001010101101001100111101000110100111000001111000010111100101111001100101000011100101000;
#1 $display("%b", po);
# 1  pi=207'b011101000110110010011110010110100111101100010110011000110110111101011001001100101010111000110010100011000000111001011101101111000001101000110011111101101010101100110101101000100110000110100100101111110110011;
#1 $display("%b", po);
# 1  pi=207'b000100100010001111001011001011001110000011000011000011100100001001010111000000101111000010101111011001001011011011100110001101110110110110000001010101100000010001111110101111000100110010101111000111100110110;
#1 $display("%b", po);
# 1  pi=207'b101010100010001001110001010111010101000111111011100010000101110101000100101110010101101101000001000100010111110001101111001100100000111111000000011000001001011001111101010010011110101100011010000111100010111;
#1 $display("%b", po);
# 1  pi=207'b011011001000111011111000000010110111000010000100110000011001001010110000000110010111001100100010011111100001110101000111100011000010100001110010011111110101100001111101100000000100010001101000000101110010101;
#1 $display("%b", po);
# 1  pi=207'b011100110011101010111110001011011110100010111110100010000001110000001110011101111001110000001111000111110001000110111010110111010000101010000001000100000000111011111110001111001000001110001010100010110111001;
#1 $display("%b", po);
# 1  pi=207'b000110110110110001111011101101111010010111010011100111010100100111011111011101001111000101100111100011100001101111011011001101010110110111101010010001001000111001101001010111000101111110000000110000001111101;
#1 $display("%b", po);
# 1  pi=207'b110001001101101011101111001001101000101000011010011100110110100011010101001010011100110110100010011000011101111010011000110000001010000011111110001100000100100001100110110011111101111001010010001001010010110;
#1 $display("%b", po);
# 1  pi=207'b100100001110110010100010011010100000011110001010111000110111110011011010111110100100010010001100111010001111000111010101100110011001000110111111111000001110011111001001110111110100101110101011011000110111010;
#1 $display("%b", po);
# 1  pi=207'b100110100101000111100011111010000110010101101101111000011001011110110101000100110010101011011100110101101111011011010011001111100110010111000010110010101111111111101101011010111000010111100110101100111010001;
#1 $display("%b", po);
# 1  pi=207'b010100011101110111100100101100100010111100011100100001101001110011011001010001001110111100111111101110001001011101101100101110011111111110100100110010010110101000001011011001011011010000011111011111010011100;
#1 $display("%b", po);
# 1  pi=207'b100111011111010111100011001110001010100111011000010000101011100001101111001011011111110100101100000100110111100000010011111111011000011110101011111110010000100111011001100111010011001110011111101111100000101;
#1 $display("%b", po);
# 1  pi=207'b011011010101001110110000111010001000111110101010000101000110000011010111110100111110111101111100110001110101010011111110101111111011011010101010110011011011111010110001110101011001011110001001110100101101001;
#1 $display("%b", po);
# 1  pi=207'b000001001011100000011001011100010011101000110001011010100110011001100110110010100111001011011000101101101110010110000101001110010101001000111110011100000100100100111001000001000111100001100110110001001000101;
#1 $display("%b", po);
# 1  pi=207'b000001110011110011101001100001100001001100100001100010110100110010010011100011000110110100001111010110000010110010111010110101110111101011001011011010011010011101101011110001101110001101111000010010110000101;
#1 $display("%b", po);
# 1  pi=207'b101110100011011010111000011101001110110010111110101010111110111110011100110100110000101110010001110011100110000001010100111001101110111001111110011001011010010110001111010100000010110110101001100010100000010;
#1 $display("%b", po);
# 1  pi=207'b110010101011101111001010010011001111001100101111011101001011001011011111001110000100000110111011111101100000010100110110100001000001001011100110010000010010010000111110000000001010110001111100101101111011101;
#1 $display("%b", po);
# 1  pi=207'b100010101100001101010101111000111101110001111010001110101000000100011001111110010110010011111011110001011110011101000010010101011111110100101001110011011011100100111011110101111001001010101011011101100110100;
#1 $display("%b", po);
# 1  pi=207'b001110000100000111001011100000100000100001011011110011000001010110100110100000100111100011111111010001011000000111000000111100111101011111010001111010010001001001101101011000111110001100100000100000010011010;
#1 $display("%b", po);
# 1  pi=207'b010011011110011110111101001000110101111100011011011100111010100101111001010001010010010100101010100101000100111000100010101011001111110111000011110101011001000010110001010100001101111100011111100011110110110;
#1 $display("%b", po);
# 1  pi=207'b011000110000000010011010000001011100000011001111001010001001100010110000011110100101111000111011110011011011101011011001111010111111011100001011001010011111001001100110101011010110011000101110011100100010011;
#1 $display("%b", po);
# 1  pi=207'b111011100010110000011100010011001100001010001110111101001010110001100000000101111010001011111000010010100011110000011100000101111110101010111010111111000101001000000010100111100000011110100001100100110001101;
#1 $display("%b", po);
# 1  pi=207'b011011000110101100111111111001001101011110111101011001110010001000111111100101000001000101011001011011011011011100011011111011010111110010011001101011011101100001011010011100000010110001001011100011000010111;
#1 $display("%b", po);
# 1  pi=207'b111010111100010100100111100110001001001001011010011100110100100100100101010100000100101110111111111011101001000011100110110101010100110001100100010001101000010011110001111011110111110000101000011000000010000;
#1 $display("%b", po);
# 1  pi=207'b110101101110011011010001001001011101010101110110110110101000010100011000001101111000110010010000100111111111111010111000110100011011000000100110111111101001110000000010100011111111100100100001100111000001000;
#1 $display("%b", po);
# 1  pi=207'b000111011100010000100010001110100101001011011001111101100010100110110001100101011011111000110000010101111001001111100010110000111101011101111101101101101101101101101000011101110001110101011000001111100010111;
#1 $display("%b", po);
# 1  pi=207'b001101110110100010010010000001011000110011110101010010001001001000000010100101110001111110110100001110011101000101001001001001001100111110000110111001000111010001100110100101000110111001101101011101111100011;
#1 $display("%b", po);
# 1  pi=207'b000010100010110101110001010001001100110100111111000001100010001100011100101011011010001101100001011000110000110101010000101010101100111000111000000010110011110110000111110100101010111000101000000000001100011;
#1 $display("%b", po);
# 1  pi=207'b011110000011011000101000111100110011001101110010011110010100010110011000101010100101101100001110101010101001110001010100100011110110000100111110111010001111001011111100100110101010110101011111110001001011111;
#1 $display("%b", po);
# 1  pi=207'b011011011100100100001110111110111001100000001100111100111101100010110010011101001101111010110011000111011001001110101010000010000001000000000111000110101101011010000001101011101100001100110011011111101101000;
#1 $display("%b", po);
# 1  pi=207'b000010110110010101111111001001101101011000101001011110101110010001110101001000100110011001010111010100111001010011110110011111000101100101100100100011100000011111111110010101011011010010100100100101010100000;
#1 $display("%b", po);
# 1  pi=207'b011011100010111010110111101000011000010001010001000111010101110100101001101000011100110100110110011101111011101011011101100101010010001110011011000100010010000001001110010010011011011010110101011010111110000;
#1 $display("%b", po);
# 1  pi=207'b001100010011011000101100011100010110111001001101100000000011011010101011110100101101000100010101000100011010010101011011111101000001000111110000111001010011000001010111111111110100000011011100110011110011111;
#1 $display("%b", po);
# 1  pi=207'b000010011100011010111011001110001000001000000000000011100101010011011001001101101110010011100110100111100110001001111100101111100100100000011001000101010110000111111101000110010010010001100101111010001111001;
#1 $display("%b", po);
# 1  pi=207'b010100001110000101011101011001101111101001000010100100011100101000100111000101111111000111110001010111100010110101100011100111010111011110000111001101011011101110111101000111011000111001110000001111110000011;
#1 $display("%b", po);
# 1  pi=207'b110001011010110000101101100100101001110011111001111100111110010011100100001001100100001010111100100001001101010100011100010010111100011011110011100000101110111110010101111111110100001011001011111111110100000;
#1 $display("%b", po);
# 1  pi=207'b011110111110111000000111101100110111010111001101000001111101011001001001001111010011011001111000111110110100000100111100010111000011100010110001000011101000111101001110010001011000000111100110010101011101000;
#1 $display("%b", po);
# 1  pi=207'b100111011011111011101100001010011101011110100101011100110111010110101010110000101011000000111000111010011011101010011000000011110000111001010110000011111000110000110011110011111010110110111101011000000001111;
#1 $display("%b", po);
# 1  pi=207'b010100001011111111110110011110101001000001101001000001000000000100001001001110111011100111111111111110010010101111001010111100100101101100110001100110100010000010101110111001000010101110001110100000101011100;
#1 $display("%b", po);
# 1  pi=207'b101010110101101101011011100000011101110010100011100000100011011110110101111100011100011010011110001100001111001000100110100000111011000110001011100011010011101000010000111111001010101111111110010001010111000;
#1 $display("%b", po);
# 1  pi=207'b011001101111101001001010101000010110001000110011100010111101001111100000111100000001111011111001001110010000101001010000100110010011111101111100010111010110000011101000111001001011101101111000101011100010101;
#1 $display("%b", po);
# 1  pi=207'b011100011101011010010011001010110100011110011110011101001100101111011110010000100001111011000100110110001111111100111000111001010110011011110110101000100011010011000111100100011011101111000111011111010100111;
#1 $display("%b", po);
# 1  pi=207'b110100000110000001000010111100100001110011100111010010010011011001000010001001001011000111010010110000110001010111111001011111001010111010001011011010000011101001110101011100000010011101011110001101000111101;
#1 $display("%b", po);
# 1  pi=207'b000100110111001101010011111001010111000011000011000001000000110111101101001001001000001010001111000101010010100100110100100110110000011101000101110100000011111111001010000000010110010000101010000110001100010;
#1 $display("%b", po);
# 1  pi=207'b001001000101010110100010010001101000111101111110011100100111000011011010101110111101100001111100111011010100101000011011110001101010011111011011110011101011111111101111011010000100100000110101110110001001110;
#1 $display("%b", po);
# 1  pi=207'b100110101110100111001110011101111101110101111010000010000001000100110001001101100000111000101110000000011100100011100110110011001101010010001011000101000010000010010100001110100100110001110001111100101011011;
#1 $display("%b", po);
# 1  pi=207'b001000110100101000101011010011011111111011010001100010011010001101101110001110111001000011000100010010101001011101000111101100010001001010001111010100000010001111011001100011010011110011110010111111011100000;
#1 $display("%b", po);
# 1  pi=207'b101010000101011010110111011110100101001010001101010000100011101111111101100100111010011111011100101111100111101010000001000100000001100101100111001100100011111110011111100010111111101101101101010110000011111;
#1 $display("%b", po);
# 1  pi=207'b001000111101110111100010111110110101000001010010111100101101101110111001010100000111110010010000101111011001111000110100111100010001100110001000001010011100001001001001110110001011101001001110101100100000000;
#1 $display("%b", po);
# 1  pi=207'b111010010110100101001110000010110111111001000010001000011111001111010100101011000111101110111111101001100001111010101111110010101111101101000000000001110001001011111110111100110100011111100010111101110110001;
#1 $display("%b", po);
# 1  pi=207'b000000110010100100001001101101010000101000010101100011110011001010110011001001001001111110110010000000101100100110101011111111100101100001010110101100101110000011111011111010101011101010011000000011110000101;
#1 $display("%b", po);
# 1  pi=207'b010011010000111110000011010011100111100101001110111111110011010111011110001000001101010101000110100110001010011010001111000011111110101001011100111110101111111110010010001001001010010101100101001011100011100;
#1 $display("%b", po);
# 1  pi=207'b101111111000011001110010110001111000110100101010101110110011000111100010111011000001100100010000001011111001011101011101000011111000001011000000000110011101001110101101100111001111101111111000100000100000010;
#1 $display("%b", po);
# 1  pi=207'b010000100110010100101011110110010010100110011110100110001011101010011100011001101001011010010100101010100100101100010100111110101000010111111101110000110001010111101001101101011001000010110001000101100011000;
#1 $display("%b", po);
# 1  pi=207'b000100000010100010111110010101111111011100100010100001110001011000111001010010100110010001000010011011101110111001001101101011110000010010110001111100101110001011100011011111010101000011000011000001110101100;
#1 $display("%b", po);
# 1  pi=207'b001000010101110100110101001011000100001111110010111011101010001010101001110001011111101111110111010011100101010000110110001100011111101000011001001110001100111010011000000000110100000101110001001010000011101;
#1 $display("%b", po);
# 1  pi=207'b010011011101001010011000001010100101101000011100100011111010000100000011111000001010010011111011111110000010010110010000011011001001000100101011101000001100101011000010001111100101110000110101001010010000110;
#1 $display("%b", po);
# 1  pi=207'b011110010010010000100100000110011010000111000010101110000010000001100001111011111100101110001110011100101001110100101110101010110101110111100111110000111011110101101111101100111101101101001100100111000000011;
#1 $display("%b", po);
# 1  pi=207'b110101110011111011110111101111000101100001000111101000110101001110000110000100011000111101000100100010001001100100111001110110101110001000101101101110010011110111000001001111000110111100110001011100110111000;
#1 $display("%b", po);
# 1  pi=207'b111000001111001000101110001110001111100001011101011011001001101111101111111111101111100111110111000100000110000010011001011001111110000100111111111110110101101110011011011000101100000010100101111101110010111;
#1 $display("%b", po);
# 1  pi=207'b001010111101101111111101111000111110101101001110000100100001110101110110010011111010001010000011010010111100011101000111010011000111111101100011110110101001111000101101100101011000111111111000100000111010100;
#1 $display("%b", po);
# 1  pi=207'b111000100011100111010100010010000111110100111000111010101001010001111001011011000010100010111111000000111001010010001011001101111000011110000000001111011110101100110011011000100111010111100010101000010100110;
#1 $display("%b", po);
# 1  pi=207'b010101011010000010101001101011100011000100001011001000111011101000010100001100110110000100101011101110001101011111001011000110011111011001000101100001000100100000011000110100110000001100001011000111001110101;
#1 $display("%b", po);
# 1  pi=207'b001000101101000011111000110101010101001110100111011110000110110101101101100110111100001010010011011001000011111101101111010010010001100010001001101011011101011001011111111110011000011000011111000000111001011;
#1 $display("%b", po);
# 1  pi=207'b011110110101110110010100000000101011001001000100010101110010100111001000000001001111011111001010110001011001011111000100001110110011000010111001010110000000001101110100010011011001001001000110001011110101100;
#1 $display("%b", po);
# 1  pi=207'b101110111110110011011101011000111010010100011011101110011000111000100100111001000000100100000101100000000000101000011011000001111111110101000111001000011000111010100011001111101000001100110100100100100001010;
#1 $display("%b", po);
# 1  pi=207'b010000010110110101001010101110101110111100011101011110011011100101010101000011111101001111110011100110010001001111000001000101001100001100110101000110011101111101010000101101110110111010100011011010001000011;
#1 $display("%b", po);
# 1  pi=207'b000000110000110001111101110001111110000100011100010101011011011101001000001010010000101011101110101000100010110000001011001101111011110110011110110011100100100101100010110001010001110000010111010000000001110;
#1 $display("%b", po);
# 1  pi=207'b101001000000100101110000001011001000100111100111011011100011000011110100001010110100011011101010011001111100101110111111001010000011000001111011011101000100011000010011011000010101100101010100011010001010000;
#1 $display("%b", po);
# 1  pi=207'b000011001110110110111000010100111001111001100100100101111010010010001010111101000101101011011100110001111110111001010001000111011000011010100001000000101111100011000111111010010001001010111001111001001010000;
#1 $display("%b", po);
# 1  pi=207'b101100001101111111101011011001011110001000001011011110011001011010110000111111110000101110010010011011100000001101011001000100000111101000001011000010111001101010111010011000110010101100000010001001011011010;
#1 $display("%b", po);
# 1  pi=207'b100010000010110110011000000100010001111001111000110000001011111111111110110011001111001110110101000001111111100001000110000101111110011101110010010010011110001111001111010001010100111000011100111101000011110;
#1 $display("%b", po);
# 1  pi=207'b100100110001001111111101100010101010110000100011111111100110001111010110001000101110001010101111000000000000111001011010011111100001001110111110001101000100101111011010010101001111011111110011001111001000111;
#1 $display("%b", po);
# 1  pi=207'b011000011010100010011101110011010111010110011011010001011000100011101011000101100110000100000000010101111110110111110111111010000110110100111101100000101110000101100111110100011101000101000100111101010010111;
#1 $display("%b", po);
# 1  pi=207'b100110010000000000101001101000111010001100000000110100000010001100110011010111110011101010011111100100110010110000000010101011010011110001110110110101101101011100010001100000010111101111110010000101011111010;
#1 $display("%b", po);
# 1  pi=207'b101100010100110000100010101000100100100001010010101111111110100101010110101111101101001000100011110100100010010011001100111000010110010010010100111011110010001100101111101011011000010110000101100011011011000;
#1 $display("%b", po);
# 1  pi=207'b001100110010000000000100000111010100110000010001000101111010111011001100001111011101110001000100001010111100111100001011011110000110110000111000101010110111100010001101000110010001011010111000011001110101000;
#1 $display("%b", po);
# 1  pi=207'b000011100110001111000010110110001011010001111011011000001011101011111110111000000010110011100100000110110100111001000101110100101011011110001100000000101110001010011111001101111010011111001001001001011011101;
#1 $display("%b", po);
# 1  pi=207'b000000110110011110111001111010010000011111110110110010011110011000000010100110010100011110101101111001000111111000101100010001110010111010001110101001010011111010001011110111111010100010101001110101000101101;
#1 $display("%b", po);
# 1  pi=207'b010111100000101110111110010110000111001010011001110011100011010111001111101111000001110001100001000011010100001000010010111001111010011011100011110110001010110010101111101100010011111000011111011100100010000;
#1 $display("%b", po);
# 1  pi=207'b111100100000111100110111110000011110100101110111010000101111100010001010101110010100110010001001011010000111100000001100010110010011101001111101000110011001111010111111000101011010011100010100011101000100010;
#1 $display("%b", po);
# 1  pi=207'b011101111010000000001110000010000000110111111111111110110110010110100110110011111100000001111000011100111110011011110100100010001001000001100010010101100100001010101001000100101110001101100110011110110001011;
#1 $display("%b", po);
# 1  pi=207'b011001010111000110011100011010000100110111001101011001001101010100110111110111011110001001101100011100110000101101001000100101011011010111000100101010111000101101001110001100001000010100100010111111111101101;
#1 $display("%b", po);
# 1  pi=207'b111110110101001111111000011100001101101001010100001010010011001010101011101101111001001111000001000000010111001110010110101010111000000100110001001101010101110010001001111110000111001101111000000111001111110;
#1 $display("%b", po);
# 1  pi=207'b110000111010100101101000101001101101110110011000000100010111100000011001101000010111100010100100010101010100010010010100011110000001111111111111011011011111101100110000110110010111111110000110111010010100011;
#1 $display("%b", po);
# 1  pi=207'b100000001011110010001111011000011111101101010011010001111101101011001000011111110110111010110001111001101111101110001000000001001111111000111111111000100010010101000111101010000000011110000011100000100110111;
#1 $display("%b", po);
# 1  pi=207'b000001011110010011010001010010101000010011100011000011011011110011010010110110011101101100011011011111000000010101110011110111100111110010110001000101011001101011100100101010111010111111111011111001100010110;
#1 $display("%b", po);
# 1  pi=207'b101010011101110100000100001100011111011000010111100010011000111001100100001000010000101100110100010111101010101111110111010001010010001001111111101011011101001000101100000111001010100000000101010010001100111;
#1 $display("%b", po);
# 1  pi=207'b111011101111000011100010010110010011000110100000000011110110011001110011000000111101100101010001111111111001000111001110110110010000000011001011101110100111111000111011001100010011011101110111011011010001110;
#1 $display("%b", po);
# 1  pi=207'b110110010100111010001011011100110010101111010111000101111001000000100111000101100000111001110101000000101110000000000011010111100101001111011110111110100111111110001101001010111000100101011100110111111110110;
#1 $display("%b", po);
# 1  pi=207'b101111001010101100011001111100111010001111010101111101011100010011111111000011010101110101001000001100010000110101101100010101110010111101100011111000101001011011001010001000001001010100111101010111010100011;
#1 $display("%b", po);
# 1  pi=207'b001001101110111010000101001111000011111100000000110000011100101100101110101100101101101111011000111000101111011011111111011011101000010001001001001010011100110111011100010110101101010011000001011110001100011;
#1 $display("%b", po);
# 1  pi=207'b011010110011001111100001001011110010010100100110001011101000110110110010000001001001100110000101001100110000100110011111100001101010000100100110100001000101100110111011001111011000010111011101101110100101000;
#1 $display("%b", po);
# 1  pi=207'b111101100010001100010101011111110111010011000011001000010111001001010010110000100010101101111000111110010101011001000001110011101000111001000011011011010100010000001100001111001001010000000111011111011001011;
#1 $display("%b", po);
# 1  pi=207'b010011101100111001011000100100100101111110101111100101000010011111010010011011110110110110010000000010010110111100000101101011101110111011100100010101011100110111110011111110110111100110110010111000000100001;
#1 $display("%b", po);
# 1  pi=207'b111101000011110001111110101000111100111101000101000100010100110001010011000001111000000101101010011110001101111110000001101100101011110111100101011000111101011111111000011000101000110000011101000100111100001;
#1 $display("%b", po);
# 1  pi=207'b000011110111001000110011011111001001000110010101010111111011011111010110011001001110101010100011111011111101100001001111101110000110001111111111111000110100100110101110000100010010111110000100111101000111001;
#1 $display("%b", po);
# 1  pi=207'b001010001000110010110011011111110100100100101110100000100111100111001001010111001000100101101000010001001111000011000011100111100011001110011001111011010000000011101110111001000100111011011101110010101110100;
#1 $display("%b", po);
# 1  pi=207'b111001011111001011010000100011000011110101110010000111101011101001000101111010000100000011010011000111101011101101100111110101011001100111011110101111100111000001011111111101010000001111111100101101000001101;
#1 $display("%b", po);
# 1  pi=207'b011101011101100101100010001001101001001000010010111111110110100100111111111011111000101111110011101000001011010000101101100101011110011100000000111110000011010000001111111011100000101001110100100100001001111;
#1 $display("%b", po);
# 1  pi=207'b101111111010000011010101101100110010100011101111011101100000000101011011000101100100110000011000010010000100011010111011100010100101111100011010101010101110011001001010111011011001001010011000100000110011100;
#1 $display("%b", po);
# 1  pi=207'b011110111101000110001010110100101011100100001111101001100010110011111100100110101101000100001001100010000100000000001100110011001011110000111110001100110000101001011000110000010111001011000111110111101111110;
#1 $display("%b", po);
# 1  pi=207'b011101101111000100010011000100011101100101001101011000000001110000101001100010100010001011110111101010000110100111101010101001011101010101000010100100010111111001100011010011111001001000001010100001010011011;
#1 $display("%b", po);
# 1  pi=207'b101100010011000111101110011111101110110100011000111110100100101000110111111001000110001101100110001011101000010101010110000101001100110110101111101110100001110101010010101011110111110011101101000010101111010;
#1 $display("%b", po);
# 1  pi=207'b001001110110101111000100100111000100011011000111000110100010100000010100110101110111010110110100101110000101001010011011010101011001000011110100101000001110110010110100111000111011001011010011000001011001011;
#1 $display("%b", po);
# 1  pi=207'b101011101111010111001000100100011101110100000101010010000111000001001000011110000000111010010111100100011101011100111110111000110000010011011101001110000011010001001000110000100110011101010110001110111110001;
#1 $display("%b", po);
# 1  pi=207'b110001000101000101011101110101001100110011011111100111010111010110011011100000100111000101001011110101011100010111100000110001110000011110101011110011101111001100100011001100100100000110000100000111000001111;
#1 $display("%b", po);
# 1  pi=207'b001001101111010001110111111010011011011101110100111101100111111111011010101111010000101010110101001110011000100001010000010011010101001001100001111111011111100001101011111010100011111011010101111101011001101;
#1 $display("%b", po);
# 1  pi=207'b000111100000010101011001101011010111110000010010011001010010110000010101111010110110011001100110010111001100010101001111101010100110010100011111101000111101011110111111001101011011101001001000111110100101100;
#1 $display("%b", po);
# 1  pi=207'b001110011111010001010001101111100100111000101000001110000010101101111101101100011110110111100111000111011100110011011101101010010010100100010000010010110110010101010000101100001110011011001001111111111101000;
#1 $display("%b", po);
# 1  pi=207'b000111011111101000001111110001011010010111011000110011101111101011011101110101001011100011110110110111000100010111010110111000010110001110001001001111110100011100000010000100101010000100110000111110010011011;
#1 $display("%b", po);
# 1  pi=207'b001000000100011010011101101111001000011101111110101101110010100011010100100001000101010101011010110100011100110100001100001001101101100101000001100111011011101100110000100000010100010110101000011101001010001;
#1 $display("%b", po);
# 1  pi=207'b110110101101011001111011011010111111000111111101101010000110111111111011101011111011100000011101001011000010001100111110101110001100000100010101111011110111100000001111000010111110101111001011000111001111110;
#1 $display("%b", po);
# 1  pi=207'b101110000101111011101010011010111101010011101010101101110110101000001010011001000111100000100101000001111111011001110101110001011111111001100101011001011101101000111010001000110010101111001010010001010110111;
#1 $display("%b", po);
# 1  pi=207'b000110110010101010100100101101010011011001100110100110111110011111011111011000010001111100000011010100111110110110110101001110101011111101001010111000100010101111111100110000110010101010011110001111111100001;
#1 $display("%b", po);
# 1  pi=207'b011110100001000011001101011111111101001101111100001100111000110011000110010111000110100000001110011011010100000000000110111101101001011100111110101101101011110100000001111011011100100011011001000010011100100;
#1 $display("%b", po);
# 1  pi=207'b111100000110010010001100001011011001110110101110011100110100111011101011110010011010000011110001101110000000101110010110111001110010110101111011010001010101101000101010001001100100101100101111010000111100110;
#1 $display("%b", po);
# 1  pi=207'b110010101000110000101101101110111110100111000100100000101011010011000000111101111101101011101011101010001100010111010110110111000000011111001101110000110011010011101101101001000101100110110111111001101101001;
#1 $display("%b", po);
# 1  pi=207'b111101111000001110000110100011110110111010101111011110110101101110100011101001000011101110110111001101010000010011001001100000010111100010011100011111010111101010101110000010000110000000100000000000101100011;
#1 $display("%b", po);
# 1  pi=207'b100110101010101110001011100110110001111010010010101000001000001010110111001001111101100111001001011111010101111101100110000101110111010010001001100100101110000101001011100100100010001100001000101011111110001;
#1 $display("%b", po);
# 1  pi=207'b111111110111100100100100000111101000110001011100010110101010101100101001011000100000000000110000100011101100011011011001100110100011101101110000000011110000111011011110100101011011100101101001101110101101101;
#1 $display("%b", po);
# 1  pi=207'b110111010101101101100010100010110100000111000010111000110011001101100001011000101000111011100110010111110101101010010001100010011111000000110101111000110100111000100000100100111100101111010001001011000100100;
#1 $display("%b", po);
# 1  pi=207'b010101111111010011001011011001100100110000111010011100111110101001111100110001100001011000111000010101001001101011010101011111001111110011111101000000110000000100011101011100111011011001011011100001001011001;
#1 $display("%b", po);
# 1  pi=207'b001110000001111000010111010110101010100010001001101101011001101111011111110110011110100011011011101001000010011110010011100001011000001111110101110011101010101110101101011101110101111111101101100101110110101;
#1 $display("%b", po);
# 1  pi=207'b000010010010111101100010010101001111001110000110101101010000101110010101000001001001111100010010000010011000101111010011000101110100101101010001011100000010011100110001100011100010000101100110100000001101110;
#1 $display("%b", po);
# 1  pi=207'b001111100101010110000010111001000110011100111111010101111001000111111110100011101110000011111111101000101001011111010110110110011101100110111000000000011110110011001110100111110001111111011001101101011100101;
#1 $display("%b", po);
# 1  pi=207'b010010101111010110001000110011011011110011000111110011000010010001010010111101101110011101010111001110011001001100111110110101101111110011000011100000110011000110100011100001010101000001111101001100111001101;
#1 $display("%b", po);
# 1  pi=207'b101011010100001110100010111110010110100001011111101000010111101110010011001101011111000100101101100011110001011100001010011101110000100101011000100010111011010010010000110111001111010000100000010100110110110;
#1 $display("%b", po);
# 1  pi=207'b011010001000000000001101100010000010000110101000001011010011100000100111000001101011110111111011101100100101010001101110100100100011011110101100101010111000111001111000101011000100110101101110001011010111011;
#1 $display("%b", po);
# 1  pi=207'b010010001101100010111000011011011100101111010001010100110011110001001001000010100101011011001001011010101100101111011000000100001101111000001011011100111100001000010101000111100001001100010001101011011000101;
#1 $display("%b", po);
# 1  pi=207'b110001101010100000001101011001010100001011010011100011010010110001101111100010100101101110110000111100111000111111101001010010000010011010001110110111111100001010011010111110101111100101111001111000010010101;
#1 $display("%b", po);
# 1  pi=207'b111000001000010101001001111111101000000001010111101101000000110110000111000010011010100101100001111111111110111100010100111100000010111010101001011000000111111101101010101110011110111100111101010111010011000;
#1 $display("%b", po);
# 1  pi=207'b001101011111110100011001111100001010011000001100100110000000100110101010100010101010110011100101011010010100010100010101011101000110011010011101001101110011010011100000001111010010001010100011010111011111010;
#1 $display("%b", po);
# 1  pi=207'b101000010001111011110110011000001010100110000100111110011011000011011110111001000001010110010111100000000010101000111001110011111011100111010000110111100001010010000011101111100101000011011100111101100011001;
#1 $display("%b", po);
# 1  pi=207'b010101111011100010011010011100011101111110100001100111011011100111010110001011101101110011110011000111111110000001101100001100110010010110110011000010000111000100001111101001110101111111101001101101001100110;
#1 $display("%b", po);
# 1  pi=207'b011010111110000001101111110100101010111111110111001101000000011110001110100010100010110101010111011000101000111011100110101000111001101110011111010111010010000110001011110011011100010111100010100111111001111;
#1 $display("%b", po);
# 1  pi=207'b000011101111111101101100110011011000110111100011011100111000011001110010111110101010110110100111011000110010100001000111011010111111011001000100111110010000111000111011011010011100000101110111110011010010001;
#1 $display("%b", po);
# 1  pi=207'b000110010101001000111111110110110100001100000111111100110001100000000000100000010011010001000011110011010101100001101101010011011111100100011101011001011110011000100111101111101010100011111000101111110011100;
#1 $display("%b", po);
# 1  pi=207'b000000110110110000001101100100001001000100101100011010101001101001101010010101111101010000101000110001111001101010100000010101011100110011001010010100001011100100101110001100011010110010001010011110010100111;
#1 $display("%b", po);
# 1  pi=207'b000010101001100000111101101011111110001100111000000011100001111011101100011000011010000100110001000100111100111101001101101100110000001100100100001010100101010100101001110111110111101100100100101100101010001;
#1 $display("%b", po);
# 1  pi=207'b001010100001000110110000001111010101110001100000011110010001010000110011001001000000111110111000001010001001111000100111110011011001100110010101011000001111101011011010101110100010111010010011111111010101110;
#1 $display("%b", po);
# 1  pi=207'b010111111001010010101100100110001111001101011100101000111110101001001110111011101100100011101100011011101011000101000011111001111001100010001111101010111100000011001000110100011010111111001011110100111110011;
#1 $display("%b", po);
# 1  pi=207'b001010000010101110000100101001010010101010000001011100011011100001000100111000111010101011000000000010011101111111001011000101001111101010001111110010101101011101010111110101101010110111111101001100101101001;
#1 $display("%b", po);
# 1  pi=207'b111000010011001000100111101010011000011010011100111100001100100000010001101010110010100001110110011001001011011010000110101111111110111011010101000011001101000011000011100000100011111101000100111101010000011;
#1 $display("%b", po);
# 1  pi=207'b110011001101010100111000001100111010111011100101000110101101010010011000100011110010100111010111110001011111101100111110001111001100110110010010110101010011100000100110111110011100100011000111110110010110101;
#1 $display("%b", po);
# 1  pi=207'b010100110110110001110011110011001111001011001100001110010100011010010010110100111110011000100010010110001010100100010100010111100110101101001011100001011010010100111010111111011111001101000010011101010110001;
#1 $display("%b", po);
# 1  pi=207'b011011001011010110010111100111001010101001111000110010011100110100011010001101001110101000111011001101100000100101010111110010000111001000010111100011110111110000100111101110101100011110001011010111001010011;
#1 $display("%b", po);
# 1  pi=207'b100010111000101010101000001111010110110110000001000010101011001111100000010100001011101011010010001100011101010010101000001010001000010011101110011000001001011101100100000001101011101101110000010011000011101;
#1 $display("%b", po);
# 1  pi=207'b110000111001100000111111100011000110100000111010010011011011000110000001001011110111110011101001001011001100000001101100110010000101111000001001011010111111011010111011010001001010101001110001101000101111001;
#1 $display("%b", po);
# 1  pi=207'b011111111111011110011010111011111010111000110011101111011011011110101001111111101111111111011101010110100001001000001100111100100010011110111101010111100001101001001110001100000100010010110101100110110010101;
#1 $display("%b", po);
# 1  pi=207'b001010011001101001100100110010000100101110110111111000110010011001011000111000011010011000000011111110001011100100100000110010111101110011101010000010010110101010001000010110100000011010011000101001001111100;
#1 $display("%b", po);
# 1  pi=207'b100101101100001100100011001110001010010001100101001100010110100011000100011100001001101110110101011110001100101011000100110010001111111011101011111101111111111011111010011001111011101010110011101000110010001;
#1 $display("%b", po);
# 1  pi=207'b101010001101010110111100001111000011011111000101001110001010000110011010011110001000100101011111100010011100101011100100100110011011011110110100000100101110001101101110011100111011100001000010011011100111001;
#1 $display("%b", po);
# 1  pi=207'b100101011101111011110101110101111010110001111100010011011000110010101100010110110101100000001110111010001001101001100100000010100011110110101000010101100101101011111010111101110011110100100001000101110101110;
#1 $display("%b", po);
# 1  pi=207'b001011110101110001101110100111100110100011010000101111000010110001010010111000000011011111000000100001010011101000101010001011011010110000101111000100101011011110111111110101000011101111010100101111000001001;
#1 $display("%b", po);
# 1  pi=207'b101001000001000110001100010100000101001010100000011010100100000101110000000101000101101000001010101011000100111010001100001000011111111101001001111100111001101100011100101110100101010100000100011010011000111;
#1 $display("%b", po);
# 1  pi=207'b101110011001010010000111111100001010000110101101001110001010011011010001110100000111010011100110100011110110110001100100100111001011000000000111000001101000011001101001001110001000001101001011000000001111001;
#1 $display("%b", po);
# 1  pi=207'b110110110101001010010111100110100000111010101111100010101001001100111001011111111110110001110110000101000101110110000111111110011100100001111010011101000100111111100100100001110100110001100011011000111010011;
#1 $display("%b", po);
# 1  pi=207'b011111110111000100001101111001111000001011010101001000101011101000110110111011101111111100111111001111111000001011111001001001010100001101101110100101010000011110110001101100001011011110000001101000010011010;
#1 $display("%b", po);
# 1  pi=207'b010111101001111011111000101001101110010101011111101101011110011100110100001110010001011100001110110011011111100000111110111110000111100010111110111010010010011011001111100011101100110110010110010010000001111;
#1 $display("%b", po);
# 1  pi=207'b011100100001001010110011111011101001011010110111011111011101101010101001110001111010100000011100111101110110001101111011100101000000010010101010010101001000100000010110001011101011000110001010011100110010001;
#1 $display("%b", po);
# 1  pi=207'b000101110100011110001000000000111011101100011001001111111001001101101111011111111111010010000010111101101001111111111110011010101001100110001110100100111011011110101000010001010111101111010001100100001111001;
#1 $display("%b", po);
# 1  pi=207'b010100101000110111000101010100011011011001000100111110110010100100101100000000010010001101011111001101010100110101110001100110011011110111010111110101100101100000101000101111000111001111001010011011101000111;
#1 $display("%b", po);
# 1  pi=207'b010011010000011101111101100001100000110000000100010001001111001110111111111111110110010101100101110010011101001100111010001100010000011110010001100101010000111001010101010011000011100101111111101101110101110;
#1 $display("%b", po);
# 1  pi=207'b011011001110100011110100011111000011111100011111101110001000100111001110110111110011010000111100001000110100001110100100111110111010011110011101101000011110010000100011011000100010110101001101110101001100000;
#1 $display("%b", po);
# 1  pi=207'b111010101010010111011001000100001101110010011010100101100010110011000010111111110101100001010100110010010001101100011001001001011101111011111010100101100010111111101000110001010011010100011010101011100000001;
#1 $display("%b", po);
# 1  pi=207'b110001000001011011101010000110001011100010000110101111011010001111100111110011011011010111110111001111111100011111110010001100001100001100010000010101111110100010100110000101100110010101101000001100010000011;
#1 $display("%b", po);
# 1  pi=207'b101000100001101100001110101111001111100011000001010000100010000110010110100010111010101101000011011100100110101001001111111011010011011101111100001011101100000010111101001000000011101010010101010011001001010;
#1 $display("%b", po);
# 1  pi=207'b111011000100111100010001110001001000001000101010001001110001111111101101100001000000011100100011111000000010001000000100101100011100110110101111001000000111110010010011001000100100111111110011110001001100000;
#1 $display("%b", po);
# 1  pi=207'b010101010001101100010000010110110010010001011110011100111000111010001011100101100111011101010111000011010011110101011000000011100111001100111010101010010110100010111100111100001101110001001110000001101100111;
#1 $display("%b", po);
# 1  pi=207'b110000001101001101010010010110001001001100100100010101011110110110100000110001101100011111011011010001110010000010000110001001000000001010101100011100110101110111010000000100111101101001010101001000100001000;
#1 $display("%b", po);
# 1  pi=207'b100011001010110011100001001100101111101110001110111000010101000100000000110111111010000110000001010111010000101100101101100000101111000110011001101011001100011111110110011001000110110000010011110000101111011;
#1 $display("%b", po);
# 1  pi=207'b000101001101100011001100101000001100000100110100010101000010001111111010101000101111010111010010000000010101101111011101111011010101011001111010100000001100000011110010000100111011100001101011010111011011111;
#1 $display("%b", po);
# 1  pi=207'b100001110111010010010100111100000010101011100000010100001101100011100000101000000111110001011111111000000001011110101001000001010111000010101001011011001000010101111010000100011110110110011111001111100110010;
#1 $display("%b", po);
# 1  pi=207'b011101001001110101111010110001111000001110001110010001001101010011110000110101110000110000011011100110010010000011100010101110100100011111001000100111111001001011010001010000100110101010110111111011111111010;
#1 $display("%b", po);
# 1  pi=207'b000100011000001010101001101001110011110100000000011111011101111000010111100001110010001111100000001100101110100111010000011110001011100000110110010111101111100010010100011100110101111110111111111111100100101;
#1 $display("%b", po);
# 1  pi=207'b001100011010111111101011111011101100011111100110011010001000111111000001010110110111000101000010001011110111011110011101100001100000100010011011000110111110010010110001011000100101011101101111001010110001010;
#1 $display("%b", po);
# 1  pi=207'b101000110010000111100011101010110100100011001011100001100010000010110111101101100011000100101000101011110011001110100011000101000011001011000110010010110100101111010110110111111001111111101011101101000001011;
#1 $display("%b", po);
# 1  pi=207'b011000111011000100110100011011001010110111011110000110111111000110100100100010100011010011010100010000010000110101100110101000110110100101100110000010100011000111000100011101101101101001001110011110100011001;
#1 $display("%b", po);
# 1  pi=207'b001110011100110011110110000100001011110111110101000011100101000000010011001100100111011100000100111011001111101011011111011110011001000110011010011111000011110100101110000111100010101111110011011101000010101;
#1 $display("%b", po);
# 1  pi=207'b110100111000000011111101101110011011100011110011100000110010111101010001001001101001100110100110001110110110011011000010100101001001100001100000110011101001111110010100110011110010010010000010011100100011010;
#1 $display("%b", po);
# 1  pi=207'b100011100110000010110111010101110001111011000010000111100110111100110011101000011011100101010110010001110010010001100000100110011010001001011111011010110110111000000110011001110111111110111010001000101001001;
#1 $display("%b", po);
# 1  pi=207'b011010001010000001110101000100110011111001110101110000001101011111111011100100000001001010000000110100011110100100110000110000111110101110101000000010110000010100111111001111100101010100001000110111110100101;
#1 $display("%b", po);
# 1  pi=207'b000001010001110011100000011010110110101011011001101100000111010000111111011001001100010100100000100100000010101001001001000110100100010110011101000000001000110011111110001011111111011111010111100001111000110;
#1 $display("%b", po);
# 1  pi=207'b101011011000000101011011011101011011101100110111000000000010100010011101011110000010111111111001001000011110011100110011011101110100011110111011000101010000111111110000010111100011111110001011111011101000100;
#1 $display("%b", po);
# 1  pi=207'b101011000000111110111010111100100001101001100010101010011101100101111100100101000100001001011001010001101101010011011001010100111011111100100111011111100101110011001001000001010110111100000001010110100011011;
#1 $display("%b", po);
# 1  pi=207'b110101100111110101000001110001000010010100010110011011010100010100010100010101100111000100010010010100000111111010110010101110110010111010000011011101001100001011100011011101000101010100001111011010000001001;
#1 $display("%b", po);
# 1  pi=207'b111111101101000100100001001010111101011011101011000101110111101100011100000010010111000010011001101000011001000110110111101011010100001111101000011111011000000100000011100010010110001010011101011111010011010;
#1 $display("%b", po);
# 1  pi=207'b011100010011010011011101101011010010111111011001000000000000101100000110000000100111110101111000011011011100011011001000001001000110011101000001000101011110110100111001111000110000101111001000000011101100000;
#1 $display("%b", po);
# 1  pi=207'b100001011000110100110000001101110001010110011001001011110100100111011100100111101100111111111111010101010111001011101111011101110111000111110100000011101011101100000000110010110111110010000010001110111011000;
#1 $display("%b", po);
# 1  pi=207'b001001000000001101011001110110000010110011000101111001001111000100100110101111001000010000100100101100111100101100100100011111101100011000011001000001010100011010101010110111010010110001100011000110000110100;
#1 $display("%b", po);
# 1  pi=207'b000101001100011001101000101110110011000100001101111001111000110110011100101100000101001110110011001101010010001001011111100011100100100000101011011000110101111100010111010101001010110000100101101011100000000;
#1 $display("%b", po);
# 1  pi=207'b011100010101000111010010101000011001000110001000010101001101011110011000010010101110000001111101111101111111111011111000110111110010101101001010001100010010101111100111111000001000001111100101011001010000011;
#1 $display("%b", po);
# 1  pi=207'b011010001101100100010010010011001011000010110010111111111010101100100110011010011001010111001010110111110110001100011111001100000001000100110010101000010010110101100011010000000000011111011010001100000011100;
#1 $display("%b", po);
# 1  pi=207'b000000000001100110101000111011111101111011101110011110101000010001010110101100100110001101111001011010010111110110111000111000100110011100110110101100101001010001100001100001110000011100011111100100100001001;
#1 $display("%b", po);
# 1  pi=207'b010010101100100101111000001000011000110010011001001011000111010100011001000010011001111111101111100000011000111100011111101011110111000001100001010001010010110011100101011001011110111001100010111010100010101;
#1 $display("%b", po);
# 1  pi=207'b110111101101010000111000011000110001111101101010101011010111001000111110100001101011001100001011000010000101111101101001110101101011011010101100110110010110001000100110000000000111110100000111000110101011111;
#1 $display("%b", po);
# 1  pi=207'b111010001000110011000111111100110100010001011011000011011101111010111101011101100000011000110000000001010001000010111000001100111110111111101010101001001111101111100111100111111111010101000110100101101110100;
#1 $display("%b", po);
# 1  pi=207'b101011011111011001101000101100111000011010001110011101111010001101010011110001110000011011110110010110001010010111011110000000011111010011101110101000111010001100100100011010111111100001111011000010010011111;
#1 $display("%b", po);
# 1  pi=207'b110010100000111001101010010000100010111111100111001011110111101011101001011101110010100101011101100111010001001000100010101100001110111101010000011111111110110100011001011000110100001001011110101101011011001;
#1 $display("%b", po);
# 1  pi=207'b101111000100100010000100010010110001000101011111010011011001010000100100110011001010010011011101000010010100101000111001000000000110111011110001010001001110011001011010101111101100010010000001100100111000110;
#1 $display("%b", po);
# 1  pi=207'b010100101101010100010011100010000111011001000110100011001001011101000011100001110010011010001111010101101011010000101110001111101111000011101101001010001111110010110000110000001110010101011101001110110100100;
#1 $display("%b", po);
# 1  pi=207'b011010110100010010010010000100010110101011001000011010110011010010111010000110010111100010111010101011100110101010101011001100111100010100000000101110110100010111001101111000000011111110101010001011110111000;
#1 $display("%b", po);
# 1  pi=207'b001101010010100110001001001011111001011100001001110110000010010101111111100001111001101110111110010110111101110010000010110110101111011010000110100111111010100100110000100000010000001000100101110110010101101;
#1 $display("%b", po);
# 1  pi=207'b010000011001110011000000011100101110011110100111001101101101011011011000010011110101111000101100101011010001000010110100000010101110101000101010111100110001010010100101111111000100111011000101110111010100100;
#1 $display("%b", po);
# 1  pi=207'b110011001010111111111011111100000101010111001100101000111001101101111101111001010010010110110011111111100001101111111011000110111101010000100100110010111111101001001100110011001001111110000011100100110010000;
#1 $display("%b", po);
# 1  pi=207'b111101010001010110001001000001000011011101100010011110000111001110100011011001101001110110101001111110010111001011110000001111111000011101011100110111101010000010010000001101111001111100100110001011011110010;
#1 $display("%b", po);
# 1  pi=207'b000111100110100111000000000010100000110110010010010101110100000011001010110111100000100110100101001001001111101111100010000000100110000011100001000001110001011111111100010100111110010010001011011001110111100;
#1 $display("%b", po);
# 1  pi=207'b011010010000010111100011111101110011011000100110100110110101000111000000010010000100011000011010000010010100110000010101100001100100010101111001111101110011100100000101001100000001010010011011101000011001110;
#1 $display("%b", po);
# 1  pi=207'b101101101110101000111111010001100110100100010111101111010101001100100111110011100111111000111110101011000011011110100110101100010111010000001100010010111101100001010100011111010110000011111001100100110010010;
#1 $display("%b", po);
# 1  pi=207'b011011111010101000001110000110110111100111100101101010100010000010011001000100010001101001001101000111011010110001001010000001111001101010100110001111011010011000101001111100010100100111110111111000100010001;
#1 $display("%b", po);
# 1  pi=207'b101001101010000100001000001100010011111101011001010101101010110001110101010110011000100111101011011111110111010111110100011001110001001101000101001001101111110101111111100010011011010100101110000111000000011;
#1 $display("%b", po);
# 1  pi=207'b111011101011100000001011111011111001101010001011101000011000010001001101001011011011111100111111001110010110111110010101100100010100010010110011010011110011101000000110011000011101000001100010111001101101001;
#1 $display("%b", po);
# 1  pi=207'b100001110101010000101110101001111011011001000000001001011101101011111011110000100101110100111101100101111101110000111000001001001000101100100110100110011110101111011000010110011000010001000100101011110011011;
#1 $display("%b", po);
# 1  pi=207'b110011000001110110110101110011100100100001010101001100100111101110010011110101111011110111111011000010111000001000011010100100100100010110001100000111010101000100111110101101001000000101000011001011101111101;
#1 $display("%b", po);
# 1  pi=207'b011000100001000010100110111000110001110101011000010110010000010100011010101111001111100110111010111010101000111001001011110001001101010011110000111010010110000110100010111101110011001010110010010111010100111;
#1 $display("%b", po);
# 1  pi=207'b011110001001101010001110111001110000100110010010000111110110010000000100101010000011001000001011111000101110011010000010111111110011110101000001111000011010000000100110010100111100100011100010101101110001100;
#1 $display("%b", po);
# 1  pi=207'b011000110001101001100110011001010011101101000101101001000000111100000100111000000000110010100101111010100111111001110101101000111111000101111001101111100110100001001101101101010100100101000010010010110101001;
#1 $display("%b", po);
# 1  pi=207'b101100001000100000100010110011000110101001010010000101110011001110100110111110001011100010101111111011101000111101100001010000000101001101010010001111100110110111010011101001110001010101111101101011110011000;
#1 $display("%b", po);
# 1  pi=207'b101100100011010000101011010001110011111011001111001011011000011111000101011100110110010111000011010000001001100000101011100111110001011111001110110000000101100001010100010100111010100101111110101000100100001;
#1 $display("%b", po);
# 1  pi=207'b010011001100010000011111101111101110111001100000101110101010010001100111101000111110001111101101101001011101101111010101101010011001010101000100011001110010101010000011000101101001000000000011101010010110011;
#1 $display("%b", po);
# 1  pi=207'b110101010000010111001100010111101111111000110100001110011111110010010011010110001000100010010111100010110010000111000001011000101111001000011010110111011011101110101010010111101101001110010110101000001100000;
#1 $display("%b", po);
# 1  pi=207'b101101110001011001011001000110110010101110100100010110111110000101101010001110001000011101111001011100011010101001001001101100110001011010001000100101010001010011100010110111010001000011111010001100010000010;
#1 $display("%b", po);
# 1  pi=207'b001010110001011110100111100111011111111011110101011110100011110111111100110100010111101101101100000000110100111100100111111101100111110101101010111101110110010011010100110100111011101100001000110110010011000;
#1 $display("%b", po);
# 1  pi=207'b011010011000011001110101000111010100010111100101110101101101110000001100000000111110000010010000110110001111101001100000111111101010010000000010100011010100100010111011000111110011110000100010000101000111001;
#1 $display("%b", po);
# 1  pi=207'b111011001100111100011100110100001000000101100110000000000110110000101010110001110101001111110000001011001100101110110000010111000011111100111110010111010110001101111000000110000110110101111011011011010100011;
#1 $display("%b", po);
# 1  pi=207'b110010100000100000001110000100101011011011100100001100100010001000101111000100000011000000110110101111010010010001101011011011111011110100001010100010100010011010010011000010011010111010000001101010111110111;
#1 $display("%b", po);
# 1  pi=207'b011110010010100001110100000111100010000111001110101011100010101100010101101110001011001010000101100000100111110101000000101000100100001110001010011100101100100110110101101100010011010101100011010100001110101;
#1 $display("%b", po);
# 1  pi=207'b000101110111000101011001001011100110011111010010100110000010011101101000101101100010011011101100111001100100110001010111000111010011001100010001111010001010011011011011110011011000110110101011111010000110101;
#1 $display("%b", po);
# 1  pi=207'b101111100011011001000101111101010001001000010100110111111110010111110110010110000000111011011111100110000000100010010000001001110011001000010100001010100101100010010101101110011010111101111110001101011000000;
#1 $display("%b", po);
# 1  pi=207'b000011110011000011110111111100110000010101010110100110000010010000111110000100001001000011000010010001110110110010011011101010110011101110001110010111001100100011010111000111000101111111001010110011111000001;
#1 $display("%b", po);
# 1  pi=207'b001000111010010110111000100111010000011010100100111100100100001100000011000111010100001001110001101011011101101010001101111101011001100000100010101010101101010101011110110100010110101011011000011110000111111;
#1 $display("%b", po);
# 1  pi=207'b110011000000001111010010010111010101001000011100110100110111100110000010010100000100111101110111110000101001001011000100110010100111101000100001111110101100000001111111001101110111100110110110011110111011110;
#1 $display("%b", po);
# 1  pi=207'b100110101100000101101011100010101011000001111111111001110001001010011110010101010110110110110100110001011110110000001011101011011001010000100000011010111011000110010001101101000000010111101011101111000011110;
#1 $display("%b", po);
# 1  pi=207'b000111011100110011100111110110111100111001111111100000010010101101111011011110100010000111011000010111010001001000101011110001010011000011100110001001101000010101011110011011101111111011100011111110010000011;
#1 $display("%b", po);
# 1  pi=207'b001101011000101111110100111000111110110110010110001100101011100100100001101110110010111101111100100101001101100110111101101011001111110000111000111111010101001011100001011110011000000000100011011010001110101;
#1 $display("%b", po);
# 1  pi=207'b100011010101011011110010001101001001010011111110000011001001010110101111001000001010101000001000111111011011101011000001101100010000001001011010010100110100011110001001101100000100111011011101101001100101101;
#1 $display("%b", po);
# 1  pi=207'b111100001101111111101110111100110100011001011000110110110111011010100111100011100101110001010101100100110101011010111000101111100010001001111111010001010101101110111110000101000110100101101110011100010100100;
#1 $display("%b", po);
# 1  pi=207'b010101000011011000011010101101011011100110100110111010001001101011000010110010010000010110000011011110001100111001111011000110110010100001101001010001010100110101101011000011111100110011001010010011100101001;
#1 $display("%b", po);
# 1  pi=207'b000010100101000111110101010000001011010000101111100011100010100001111011111101101010111011010000110101111001110111110011100111110011010010101001011110000000100100111011000100111100011111010001010010111000010;
#1 $display("%b", po);
# 1  pi=207'b111011111000001100100001111000000001010100000001100001000010000010101010110000000000011011011101001010010001010001001001011001010001110100100101011101011010011011001010010110010101100111011101000000001100010;
#1 $display("%b", po);
# 1  pi=207'b011101100001001110000000001110111000000101110000011000100110110110110111101101010110000111001101000000010101000001100010011101001000111011010010110110011000010110101111110100111111001111010011000111101110111;
#1 $display("%b", po);
# 1  pi=207'b100110011111011010011110111100010011000010001110110000010010101101010101010110000010010001111000100011101111011010001111101000001000000010111000110111110101111000011101111011101000000101111000001111010111111;
#1 $display("%b", po);
# 1  pi=207'b000011110000011000111010101000110001100101101100101101101100011101010010000010001000111111100011011001101010000100100101000110100101001101101110000101111010111011001000011010100001101000101101100110101101001;
#1 $display("%b", po);
# 1  pi=207'b010100110111011011111001101011010000001110110101110001101110100000100010000001011111000101001100101101000001001100011001001110001000000010011000001000110010101001000011011111111001111011000010010111001101101;
#1 $display("%b", po);
# 1  pi=207'b001010011111000010100011001011101101000011011101111111110010100111000101000001011100111010111110011001001110110001111100111110010110101000001111100011110111111011110101001110011111000011100110011101011111100;
#1 $display("%b", po);
# 1  pi=207'b001011100000111001111000101100011100111111100101011101011111010100101000110111010001110000111100010101110011010101010111000110010110011011000010001001011001110110010110101010101100010110111100000000111101010;
#1 $display("%b", po);
# 1  pi=207'b110000110011010001001000110001101011011011011110000011100101000011100100011011111011100101110000100011101010001100100001000100110110111010101110111010011011110110001011111110101110100100100111100111111000101;
#1 $display("%b", po);
# 1  pi=207'b111000010100011001101101001001000001100000100000011001110101001100000110111000100001101000101101011111011110100111010010011000011111010111001011100100010011011100111000000010111010010111000011101001011100001;
#1 $display("%b", po);
# 1  pi=207'b101110010011011001100010100101110011111110100001111000100011100100101100001110000000100000011100100101101101001011001101011111111010101100010000100001101001010110001001100101100010110101011110110010111111000;
#1 $display("%b", po);
# 1  pi=207'b000111100111101001110111101110111101110110111101100010101011101101101101110101010010000001101001101011100010001010000010100010000010101100011111001111111010111000000000000110111001010000000111100011111000011;
#1 $display("%b", po);
# 1  pi=207'b101001001111101101111011000100110111010010110000101111111100001110001011000101110110101010000110101010100100011011001000101100010001110010001011001101000000000010101010111001101101111011101111010101010100100;
#1 $display("%b", po);
# 1  pi=207'b001110100110110100101000010101001110001011101000000000011010111111001101111110011010110011011100110111110001101100101111000001111011110101000001010000101111100010110010100110111000000100110111100111100101000;
#1 $display("%b", po);
# 1  pi=207'b011111001111111000001000110001111110101010110000001100010110111000001000111100110100011111101100000100100000101001101000001101000000010110010111100100111101000011011001011100010000010000010011101110111010101;
#1 $display("%b", po);
# 1  pi=207'b111001100111100110111001011100001110000010100001001111011100001101110101101110111111111001111100100011111010101000010000111011110011110111000011011001001001101010010010011100101011001101001110110010100000101;
#1 $display("%b", po);
# 1  pi=207'b000111100000110100101110100100000011111011001011100001001011001111111101101000100100111101110111100110110001101010110011111111111001001011010000101110000100101000011000001000010011111010001010100110001001111;
#1 $display("%b", po);
# 1  pi=207'b001110111101001000010011000111010100110110001111110001100001000110000010101011000011100001100001111101110101100111010011010100101010100101101001010111001100000100010101000101011011000010011010101100001110011;
#1 $display("%b", po);
# 1  pi=207'b111000011101101100111001011110001001010001101100100110101011111110110001011111001010001100001010001111100001000111011100111000010110001001010010101000011111110110110010110110011110110101110100010001111100101;
#1 $display("%b", po);
# 1  pi=207'b010101001011100010011010101111111000110111001000000110010011100000100011010111001110110000010101001010011001011111111011010000110011001100100010100101011010111110010010111001101100001000010100011010010000010;
#1 $display("%b", po);
# 1  pi=207'b000011111110000100010010000111011010110100100111000101110010101000010011100100101011001110001110111010010110010101110101100111010001001101101001001111010111011110101101111110100111000100100011010001111011001;
#1 $display("%b", po);
# 1  pi=207'b110001000110000001010010000010010101001110010001100100101010100110000000000100011110100000011110100101110100110110000000010001100000110110010100111001001000100101011011101010101111111101011101110100110001110;
#1 $display("%b", po);
# 1  pi=207'b100100101001000100000100110010010111001110101000111110001001000101100111101101001010010001011011101001010011110111111110111000101100110000101111101101001001100111011001010000011100001000111111001100100011001;
#1 $display("%b", po);
# 1  pi=207'b011100111000100100011110001010101011001111100011101101010101011111101000011010011011101000001011010110101000001101101111110001011111101100110101111111111111001010101111010011101001000111110110000110100010001;
#1 $display("%b", po);
# 1  pi=207'b111110111001100111001001101010110111010000101011111000101000110001011011101100110111110101001100111101100010110010101001100000010100110000100000001000100101001001110101011010010001010010001011111010011101101;
#1 $display("%b", po);
# 1  pi=207'b011110001101110011111010100111101000000010000010110010101101111000110100100010010110000011100010011111010100110111010111011101111100000001101010011101010101111111011101010110100010010001011000001101001101000;
#1 $display("%b", po);
# 1  pi=207'b101011100011010010001100000000000010100110001111011010110011011000011100001010011010010111000010001001000000101101111111101100110000100011000110100111011011011000000000001010101001000100011000110100010000110;
#1 $display("%b", po);
# 1  pi=207'b101101001010011110100011010111000111110111100010000010110001101101011011110111110011111010101110001110111010011011100001011011101100100101110000000110001010110100100110011010010010111010011101000101100111101;
#1 $display("%b", po);
# 1  pi=207'b110111100100001111100011100110011110011110100011011100110111000010101110011110001110011110011001111100010111111000110001100110001010101011001010100010001000110111001111001010000111110100100100101000111000001;
#1 $display("%b", po);
# 1  pi=207'b001000110110010110001110110111010001010000101100000000011000010100001011101111000000010001011101111000000111100010011100011111101110101000110010001000110110111101011001111011010111001101000101010011111001101;
#1 $display("%b", po);
# 1  pi=207'b110001000101000101101101100101110101110111110000101100111010011010100111111101111000000000001000010010110110101111101110111011010011011001001111111000110010100011011000111100011001011011000011100100001100000;
#1 $display("%b", po);
# 1  pi=207'b000010111000001101001111010000001001100011001001001011011110000111010111100110010010100011010100001101100011110000001001110010011001011101011110011000000010011001000011011111011000101100111111111000110010010;
#1 $display("%b", po);
# 1  pi=207'b110001101000110110001110000100110001010011101100000011000101010010000100010010011101101101111011100001001000101111000011011110111111011100101101110010111111001001100001010011111011001001000100001101110101000;
#1 $display("%b", po);
# 1  pi=207'b010000011110011111100101001001000010100101111010100110001001001100111010001100110000001100010100100010001110000111000111010010100100001101000111111011111000110010101110000101000110010010111010010000001100111;
#1 $display("%b", po);
# 1  pi=207'b001010110100010111011110010011110011010010000011001101111001011110111010110111111110000101000011100100011101001001000101100011101110110001110111001101011100011000111000000110111010100010100110000000000100100;
#1 $display("%b", po);
# 1  pi=207'b101010111111101010110100101011110111110010011011101001100100100010111010111111010101100011010100101101010010110011010100010001100000100111100010101011101110111100101010000110011100001110100011110001011101100;
#1 $display("%b", po);
# 1  pi=207'b101100000000100011001100111101000111100000100001011001011101110101110101000010010100011111110010101101001101101111010011100001011011101100000001010100000100001111010110001000011000001111100111111111011001000;
#1 $display("%b", po);
# 1  pi=207'b111011001100100111000001000101011110010111110100010011000100011101111010111101011101100101101001111101011110010101000010001001111111111111011111010100111101111011100011101010000110100100001000111101111001010;
#1 $display("%b", po);
# 1  pi=207'b111000000001010001101110010011001001100000101010110100100010001100001001011001111000111010001011101000000111110110011101010111000010001101111010101011010101011010101101001110000101000100011000000000110001110;
#1 $display("%b", po);
# 1  pi=207'b011110110100011010100010100101110001000011100000001111110111101001101101100001011001000101100111111011010011110000001011100110010000101101011010101110111111110101010001101111101110101001001010111011000001101;
#1 $display("%b", po);
# 1  pi=207'b110101010100001110010011110010010101110011010110001110001000100111010011010001111001100111001011100000001101100111100111101010101100110011111011101001010010011000100011010100000100100101001100101100010000101;
#1 $display("%b", po);
# 1  pi=207'b001101111010111100000011010110110100101011101101000000100111010001111011100110111101100100010100001111101001111011010111110111001100101011000100011011100101011111100111110110000100110100100000011001001011001;
#1 $display("%b", po);
# 1  pi=207'b000100001011101001101101010000110000001111011100000011101110100101011000011110000011001111000110110000011001000110101101010010010100001111111100111010101011100001001000000010010100000001110001110000101000101;
#1 $display("%b", po);
# 1  pi=207'b110111010000111110111101011000110110111111100111000111100110111010001011010100100001010100110110101011111001001100010101011001101100001100011010110011110000110010000110100001010111110111000011111100100100101;
#1 $display("%b", po);
# 1  pi=207'b101110110100100001110001011110011100110010000000101100101001001111001110010101010110000010000011101001110000010100100011111011101110110001011100101010111010111001001100111101010001111011100111110111010000100;
#1 $display("%b", po);
# 1  pi=207'b110010111010011001001000111001110110110010001111101110010011010010010110001111011100010101101001001101110011101010100110010111011001110111001010000110100110110010110000100000000010001000011011111001010101000;
#1 $display("%b", po);
# 1  pi=207'b100100001111101011011010110101011110100100010011011101110101011010010101010110000111111010011010111111101100010101001100110010000100101010000101101011101010111101111001101000001110100101011110110100011010001;
#1 $display("%b", po);
# 1  pi=207'b010010010010110000010100110000010000100001011011011110111111101001110101010111101001011000001001000001001110010101100000010000000110000010101010111110110001101010100100100010010101111001011010101000011111010;
#1 $display("%b", po);
# 1  pi=207'b011001010110001010010001110101000010011010100001100010010100010011001111010010001000000111100001010110110000011011111100000001111011111000011000111111011110001100001110000001100111101000101101111010101010101;
#1 $display("%b", po);
# 1  pi=207'b001101010000100010110111110101101101111101001111000100111001011011011000001110111001111101101111110101010011011111000111101011011011010000001100010111110110101001111110101011110100110000101101100010111111010;
#1 $display("%b", po);
# 1  pi=207'b100101111001110110100010001000001110010100010001001101001010001100000101000110100011001001001011001010010001100000110010110010010000101011001010001010111010101100100000101111100011110100110111101100111010100;
#1 $display("%b", po);
# 1  pi=207'b001001101011101101100100101110111100101001000101110100111000110111001110000110110011111100011011001010100111111110010101110010110011010100111100010100100100010100101010100010111001001010001001101101011000001;
#1 $display("%b", po);
# 1  pi=207'b100001000111000110010001100000101111101001011110101001001010101000011100100001001101001010011101111111111001010011010100011110011111001001111011101011011001110010100011000011011100011101000000010111110010110;
#1 $display("%b", po);
# 1  pi=207'b110010111111100000000101011011101000110000101111010001011000100100000100110100111110011111111111000101100111001011011101111001000100101101000000101111010111100111000111010111010011101101101001111100010010011;
#1 $display("%b", po);
# 1  pi=207'b000001101000001101011000111111010100001101010111110111011111010000100111000110100001110101011010000001000111111111101000111101110110000110001111101001000110111011011001100110110001001001011011111110001101100;
#1 $display("%b", po);
# 1  pi=207'b101101001100001110001000101000101010110101000111101110111001000100010101100010100010001101101101110000110001111011001010100000100110010001101011110110100100101100011110000011101010101010011001100101011001010;
#1 $display("%b", po);
# 1  pi=207'b100100110110001100001101101000010101101000110100111111111110110010010000000110111101010110110110101011100111000001010111110100101111100111110000101100100100010011000110000000011000111011111111000001111010100;
#1 $display("%b", po);
# 1  pi=207'b010100010000000111001101000001100010100111111001010100111111100100000000110001001011010111110101001111011110111101010101000111001100010101101100110101001110111011110000101110001010111010100110110101100000011;
#1 $display("%b", po);
# 1  pi=207'b110010000011001110001001100110001000011000110010110000100000001011101010000101101111011001001011110110001011111100001011111101000010010110100100011001110011100101101001100101111010001010010100101000010011001;
#1 $display("%b", po);
# 1  pi=207'b011001011101001000000000111001110010110001010111111111100011011110000000101011111101111111101000111110001101111110101010011111000101101000111100111000000011111110001010000110001001000111010001101100010110110;
#1 $display("%b", po);
# 1  pi=207'b001010100000110001000001101110101101001100111100100110011100111111110111110011000111110011100101000101100010001110101010110110010010000111001101111010001001111011110001110111011001000011100100011110100110000;
#1 $display("%b", po);
# 1  pi=207'b101100101101100100111111111110010011001010110110000010110110101000100001111000110110011101000001111011011101111011010010000110000110001010110111111011110110000011100000010110001001111100111111101001010100111;
#1 $display("%b", po);
# 1  pi=207'b100101010110101010110100000101011101000100000011101111001010010001001000111011100000100111100001000111101110000101111101100001000110111110100111111000110101010110000011000000001000000111110101011110101100100;
#1 $display("%b", po);
# 1  pi=207'b101111011110110111011001100010100000011101100010111111100001001100100000101010000100000110000000111000011000011111110101100001110111001011011010010001010010000110011100001101000001100110000010100100010010001;
#1 $display("%b", po);
# 1  pi=207'b101001111101100010011101111101011010010001111000111111101010000010000110101111111110011110001000001010001111100010110111101111010110110010000001000011000010010011111010001111111100110010110010100110010100000;
#1 $display("%b", po);
# 1  pi=207'b100111101001110001000011111101000100011101000111111110011111011011100001000100000011110110100100100000011100000000110111000110111100111000110110111000110101100010111000111011001110101100101011000001011110010;
#1 $display("%b", po);
# 1  pi=207'b101001000010010001000000001000101001101001101100010011011011011000101101111000011011011100000011001011100110100110000010010011100100101000000110101101100010100011011111010000001111101001100011101001110110110;
#1 $display("%b", po);
# 1  pi=207'b011110101100010100010101100000101010101010100010100110111000000101101011001111101000111000100111110001011011011101000000000010110110101010111101111011001100001011111111000000010111111001010110000101000111111;
#1 $display("%b", po);
# 1  pi=207'b100000011111010011011101111100010000111101011111000011000101110010101011110011111111110011000010011100101110100100100001111001001010111111101111010101011100101110011111101001101111111001001100001011010001000;
#1 $display("%b", po);
# 1  pi=207'b101110100101110001000111100000001011111111111001100001111011111100101101110100100110010001011101000110100100110100001011101010101011111110011100001000000001001100100111001110000110100111110001110110100000111;
#1 $display("%b", po);
# 1  pi=207'b000101101100111110101111000000001101001011001110101111011111101011101100000100010100000001010010011000011011100101100110001101110000011010111001001111000000001101110001110110100010101011110000010100011001110;
#1 $display("%b", po);
# 1  pi=207'b000010011001010000110000100111101010100000111101111100110010100000101100110111010110010000001000111001010010010001000100100110100011001110111001001111010101110000111111011011111100100011010001100101111001100;
#1 $display("%b", po);
# 1  pi=207'b110100001010001001100001011110010101010010011000111011110000000100000000011001001111001010000100000011110000000111001111100011001010111000011110011100000110011010100101101010010111000111011110010111001011011;
#1 $display("%b", po);
# 1  pi=207'b110101100000100001111000000100000101101000100110010100000111001110010000000101000110101000000110001011001010000011011111101000111111011000111000001010100011001010000101110000001101011100001111011111010000010;
#1 $display("%b", po);
# 1  pi=207'b000111000000111101001100100011000101001101110101011110001111110111110100001101111100001100001001111000001111110011100001001110111111111101001011010111010010101100010101011010111001101110011110100000000010000;
#1 $display("%b", po);
# 1  pi=207'b111011110001001110010000000100100010100010001100101001000101100001101100010001101100010010100010110010100000110001010110101100100001000110110110100000101110111010111110000100010000010111010111011011101100001;
#1 $display("%b", po);
# 1  pi=207'b001000100100101011101000111100110011010100000010101101001011001011110010000010101111010001001111111101111111100011000100100101100111101100011001000111001011000000111000110001000001100111111110010000011111110;
#1 $display("%b", po);
# 1  pi=207'b100101111000110100110010000111111001101001110111010101001000001000110111110111011000000101010100011101100010010010001010000101110100100100111010011011100010010101110011011101111111010011011001001010111010100;
#1 $display("%b", po);
# 1  pi=207'b100011100110010101001011000111100101011111110111010000101011111010100110100011110100100001011000001110000000001101001111010001111011010001001001100001010001111100010010111101110010111100100011101011011010101;
#1 $display("%b", po);
# 1  pi=207'b101111101010001111011011110111010010000100010011001001010110111101110010001001100010001110011111011000010000101010000111111001111000110010100101011011010010010011000100010011110100000001011101110010110111111;
#1 $display("%b", po);
# 1  pi=207'b000011011010000000010000001010001000111101000111010100010100000001100000101000110001011100100001001010000001101101111111111101111100010011011101101010010010100111100101011000111000110101101111010010110001101;
#1 $display("%b", po);
# 1  pi=207'b010110010011010001100011011110010100010101001110110010100100101001100001000111111100011010010111001000000101000100011000110100101111101001010000101011100110101111000000010000001000111111110100111011011001110;
#1 $display("%b", po);
# 1  pi=207'b101101100101111101011111110000100110101111111111101010100001001101000100100010001111111001001011101001010000110011000001001001001011000010101010101111011111001011001000001000110101110111010100010101011000100;
#1 $display("%b", po);
# 1  pi=207'b001010011101011011100010010101100011100110110010001110111101010000011111001101101111110011001111010011110011001110010100010010010111100011010111001010011001010101110000110010100011100111001010001001010110110;
#1 $display("%b", po);
# 1  pi=207'b001101010011010111110011010000101011101000001111100101000110011000010011111001000111101101000111110110111001111000011010101011011001100111100011010101101111010011010101001000111010000100010100110100001000001;
#1 $display("%b", po);
# 1  pi=207'b010011011000000011010011111101001010110011110111000001101100000010000101110001101011011000101100101011110111001101000111100110111000111001110000100101111100100010001001010110010011001101000110001101010111011;
#1 $display("%b", po);
# 1  pi=207'b101001001011100001011100011100110110101110110010010000101100010011000000010001001000110011110001000110101111101111110110101100110100100110010001100000010110011000000010000101111110111100101000000010111001000;
#1 $display("%b", po);
# 1  pi=207'b000100101101100000100011011111101000001100001011001001111011010011000010101110101000111010000110000100111000100000010100101111100010001110001101010000001011101001110001111001110111011011100000110100101101101;
#1 $display("%b", po);
# 1  pi=207'b100000101010101111001101101110100100110000111111101011100100000000101100111000001000010100001001111001100101111010000110000101111110110001010000001100111101001000110101110100000000010101000111111010010101001;
#1 $display("%b", po);
# 1  pi=207'b001000110110111011011100010101011111010101111011101011110001000110111100011101001111010101110111100001110101100100101100000100111010111011101111110100100010000101000110110111101110110000000001011001001100001;
#1 $display("%b", po);
# 1  pi=207'b001100110000101011011111100101000011111011011101000001111100010111001101110010111111110101100010010101001101110010000000001101100101011010010101101111111100111011000111010111101000011010100110110000111111111;
#1 $display("%b", po);
# 1  pi=207'b010000011110011000110110100110011100101010001010100001001110111100000010100100110101010010101111000111100110111011000011000010101010111110011110101110111010000011101100001011110011010110000100001111011100001;
#1 $display("%b", po);
# 1  pi=207'b010110101111110011011000100001100111000001101011100101100100101101100000011011011101100001100100011111101100110010101000010000101001001100100011100010101000101101000111011001000100001010101011100000001000101;
#1 $display("%b", po);
# 1  pi=207'b011000000001101000010100111110000100001100001110100010011100000110111100100111110011101011011001010100110000011111010101100000000000101010101101110100000011100010101111101000001100100110111110100111000011010;
#1 $display("%b", po);
# 1  pi=207'b101001000011111101110111110011010111001111101010101011000101001111010110101101100101011101001101011110000101111111000100111001111000111011001110011101110001101101100011001100111011001111000011111100011101110;
#1 $display("%b", po);
# 1  pi=207'b010011101000100100111101100111011001000001100010110100101100101100011101000111100000011000110010010010111010011000011111010110001001110001010001010010101011100101110001100010001111000100010111110001101010010;
#1 $display("%b", po);
# 1  pi=207'b100111110000110000001001100100011000000001011100001111110000010101111001011000001110111001110110111010111100001101110011011100011000110000101000111100000000011100000010000111001101101011001010010110010101101;
#1 $display("%b", po);
# 1  pi=207'b011100010010111010001000000000000111100000010111000100011111110110011011000011101110011111110010000111011010010101100010101010101100110011001110110111001111010000101011101111011100110000000110001101111101110;
#1 $display("%b", po);
# 1  pi=207'b110000100100110110101110000111110001011100111101111010000011010010010000111011001100101000001110111101111000000110011101000111000101011000011001001000000000001010001011101011111010111101000000011101111010010;
#1 $display("%b", po);
# 1  pi=207'b010010100001001111101001100110110010010010111000101001001000110100111100110111001111010110100011001001011111110011010010001101000111111000110110101000011010010100100010001111010110010010000010101011001111101;
#1 $display("%b", po);
# 1  pi=207'b010110110011101100001100110101101001110101101000111001100000110100000011100100111101001011111011010001111000101101100110110101111100111011101011111111010101110001101010000111011001010000111010100010101010100;
#1 $display("%b", po);
# 1  pi=207'b011001011000110001011000011000111110000100010010011000100111111000001000110101110111111111001001001001010001111111101110010001001010000101011010101110100000001000000000000111100110110101001000110111110011100;
#1 $display("%b", po);
# 1  pi=207'b010111110100101011110000111111100011110001010111000011110110001101101011010000010100111011001101001011100101100101000001111100101111110010000100010011011101100001000101101100001010000100000111111001001111110;
#1 $display("%b", po);
# 1  pi=207'b001100100111000011101101100011000110110010001001101111001001110011000011110101100111111111000000111100101111001111000001010110011001011100001111000110010010011110010001011010011000111011101011110011111011110;
#1 $display("%b", po);
# 1  pi=207'b011100101000010111011100010110111101101001111001001000011110000001100010000100001000000100011001010010011110111011000111011100001000111100110101111010001011010101011100000010100001111010001000101100101110100;
#1 $display("%b", po);
# 1  pi=207'b101110000110111100100011011000110011110110100100111011110010111100101000100001111000011101000111111001011010001010110111000001010000101111101000101001110111101010010101001000000111010010010000001011000011111;
#1 $display("%b", po);
# 1  pi=207'b010100110100110011001101111010010110110100001001000100011010010001001010011010000001011110100011111000110000001011100000101100110100000100010111101110001010100101101000101101011110010111001110101111110010110;
#1 $display("%b", po);
# 1  pi=207'b110100111110100100110010101010100010110011101010100001000010010011110101011100110000100010101010000010111111100001011100000111101011001010100100011110010101001011100011111001010011001001000010110100000111010;
#1 $display("%b", po);
# 1  pi=207'b101001000110000011000000101110011001101001000011110011100010101000010101101111010010111010111100011111001111110001101000000001011111101100001101011100010001011001011000100101100100110110000000010001110110111;
#1 $display("%b", po);
# 1  pi=207'b001000110011011100100011101010101001011011010101100111001100111110011111010001110011100010010001000001011010010100100001101010001100001011011100111111100010110011110100011101000101011101011110001111101110110;
#1 $display("%b", po);
# 1  pi=207'b011000100010000110110001100100111100010010001111101001100111100110100101011101100011011110011101111001001110111001000100110110010000101101011101011010010110010010011100101010100111000011010100110100001111010;
#1 $display("%b", po);
# 1  pi=207'b010011101101110011001111110001110001110000001000010100111110011011100101000001111100111101001000100100111001101111101111110001111111000000111001010011000000111001010111001101101000110101111110110011011111101;
#1 $display("%b", po);
# 1  pi=207'b111110001111010100110100011000111010000101011001101001101010111100111110011101110111011110000110101111111001000100101000110001101001010110000100110110110101000110010000001000100110111011110001000110111010011;
#1 $display("%b", po);
# 1  pi=207'b010100101111111110001000011100011101001110011000111101010011010111011011010100111000100111101110110100110010111011111101101010001000111110100010101110010110110000100000111110001010010101100110110100000000011;
#1 $display("%b", po);
# 1  pi=207'b100101111111101001001101111010100101100111100100110110001100010000011001001101110000100001101111110001110001011001011010011100100010110110111010100100010000001110001110001100110100110110100110001111001011010;
#1 $display("%b", po);
# 1  pi=207'b101001111000110110110001100110111110100001110110110001010101101000111110101100111111111011111001011001110001010000000001111010010001110011011010000101100010000011100001001010000011100101101001010000110011110;
#1 $display("%b", po);
# 1  pi=207'b101100011111011111100100100011101101011000010101011011011011111000000111000011000101110100011010111110100101000010011000000100010011100110010001010110100000001000101001000100100101011000110010101111010000110;
#1 $display("%b", po);
# 1  pi=207'b011010010111010001011001110101011010011100001000101001011000101100110101000010110111100010010011111000001101011010001011000110111000111101011101101000111001101101010011000000011011001110101000011010000100001;
#1 $display("%b", po);
# 1  pi=207'b100110010010100001111000001101011000111000000100101011001000010001000001010000010010100001010000000011100010111111010000110001101110100100100010000100001101000011110111110010100110011010001101001000000101111;
#1 $display("%b", po);
# 1  pi=207'b001111111011001101001101010000001000010011110001001101010010010110010110111101011110101001000100101010000000101000100010110010101011110110100011011011100110001010000100010101101001010110111000110011111101111;
#1 $display("%b", po);
# 1  pi=207'b110101101000101101010100111001100100000100101100010011100010011000101110111000100100100100000010110111001100010000100010010000011001001001011010101111101000010100100100110111100111111101000101010001011100100;
#1 $display("%b", po);
# 1  pi=207'b000110001001000011011111011110100110010000000100001001111110100100101101101010000111111010100100111101111110001100111100101110110011011000111001010000011010000110100010001001111001110001010001110101001110000;
#1 $display("%b", po);
# 1  pi=207'b001100100110111101001110101001011000001001111001010011010000001101110001100110001111110100011010011101000011010001101010000101100111011111001000001010111000100000010000110010011100010011100111110101100100100;
#1 $display("%b", po);
# 1  pi=207'b011000010101100101111101001011100100001011000111100010100100111010100110010110110100101011101101000111100000001001011010001011100011101000010110010000100111001110001100011010110011110010101001010110010010000;
#1 $display("%b", po);
# 1  pi=207'b010110011000101110110011000010011100111011010000110011001110101111100001110000110000101110100101010110110011111110100010001011011001011100110010110110000110000010110100100100101011010000100101001001101101111;
#1 $display("%b", po);
# 1  pi=207'b111110110101110001001001100100001101000000110110111111011100010000000010000101110101100000110100101110111100011010010111001000011001111011011001000001101100001100101100000011100000110111111011110100001100010;
#1 $display("%b", po);
# 1  pi=207'b010001000101110101010101010111111010000101101100001000011000011100110010010001110111001001000100101011101110101001110101111001001001010110001100100101011111001001101001010000110111001101001101001110110000101;
#1 $display("%b", po);
# 1  pi=207'b000000000001110011000010010110000011111010000110001111010100010011101011110100101101001010010101010001111101101101101001101010000101110111100001111110101100001101000110110010001000010001100110011111001001110;
#1 $display("%b", po);
# 1  pi=207'b011101100110010010101101110000010101111100100000101001110000100010110110000100001111010011000000100011000111111110001011101111111110101101111001101110000111010010011001101011111000000000001000100110100010010;
#1 $display("%b", po);
# 1  pi=207'b101000010010110001101110101001101000000101100001010100010011100101110101110100111000111011111010000100011110101110101010101100110110010100100101001000010001011011110100111111010111011100001010100000110000000;
#1 $display("%b", po);
# 1  pi=207'b111111010011000101000000111011001110100011001101001001111010010110000110010001000001010011011000011000101111011010011010010001001010010000110111110010000001100110101100100000001010100101001110101010110000111;
#1 $display("%b", po);
# 1  pi=207'b011110100010101110110110111011001111001010000000011101111011010100010010001110000111011001101001010111110010101100101111011111101100100111110010111000111010010110110111100000101000101111110010101110000100010;
#1 $display("%b", po);
# 1  pi=207'b111011001101001110100100100010001010111010101110001010110010001000110111110111001001101110000000011111100100010111010101100011001010100000001100000110101010011111101010100010110010101111110001001010001110000;
#1 $display("%b", po);
# 1  pi=207'b111001111010100100001011111111010111001010001010101100100111001101001001111011111111100011111111000010101001111001011010110010000010011001001110000100110000010001110010011010100111111010010011101000000010100;
#1 $display("%b", po);
# 1  pi=207'b011010110010010010000111000110111010010111000001001000011111101000011110000101101111011111110000110100000011111110001100001001000110101010110100001111100010011010001000001111000011111010000010111010110000000;
#1 $display("%b", po);
# 1  pi=207'b111111110110110111010001111111011000101001101111000100111110110110110100111100001011110001110010101010111101001010000000000110010010011110101010100000110011110100100101000000011011011000001011000001010010010;
#1 $display("%b", po);
# 1  pi=207'b100101011100110110111011111010110100111001101000001010001011100010000011100100110011111100010101111010010000011101110000100011011111101011110011010011011001101000111010000101101100001111000101111110010000011;
#1 $display("%b", po);
# 1  pi=207'b011101000011110010111101001011010100100110101011000010011110100010110101000001110000010000010011111010111111101101101000011100100011110000110111011010010101011001101111000010000100011100101010000000011001111;
#1 $display("%b", po);
# 1  pi=207'b100010011011010100110011110010111010011110100101011011101110010111010000110110011010110010100001000100000101101001111110100101101011110010110111110000100010111000101010001000011111100001001111001110000011111;
#1 $display("%b", po);
# 1  pi=207'b011100101001110100101110011101101000011001101100100010010110001010011110011011100011110101100110000100011010111000010000001101110010001101010011011010110010000111100100110011000011000001001100110110011111101;
#1 $display("%b", po);
# 1  pi=207'b000101010110111011101010001011000101110110101101000001000001001100010101101011110000001101100010110000101000000111101011110011010000011110000000110001110110011100010111111100010101010101110101111010001100111;
#1 $display("%b", po);
# 1  pi=207'b101111010001000001101111111000101010101000111000010000011111111000101110010111011111010001000000100110010001111000111011010011010111110100110001000011100001110010101001111110010100110011101010000010000001100;
#1 $display("%b", po);
# 1  pi=207'b111110000010011111010010111010100000101101001001101111000011011010001001110010011001000100111010000001101000011001011110111100101111011011010101101010000010101101010111010000111110011001000001000101110000011;
#1 $display("%b", po);
# 1  pi=207'b101101110011101111101011001001100001011000101101001110001110111100010110100001110100111111111010010011100011110111101001100111000110111010001000010111110011101001111000110001110010000101010010000001000111101;
#1 $display("%b", po);
# 1  pi=207'b000110010011011001100010111100111110001010000001000001101110000101010100011000011010001111110001000111011001001001011110000011000111110100000010110000110011111111010001111111101110010000100010111000000001011;
#1 $display("%b", po);
# 1  pi=207'b010101001001110101101110001010011101001100001001111110000110100000011110100011111111010000110100001011011011100110001010010001011011111001000110101100010010011110100110000110111001001100110000000011001011101;
#1 $display("%b", po);
# 1  pi=207'b111001100100001011001101101010100001111110010101100100010011011010101100101001011111001110010001110000010001100100001100011011101101110001011100010100111110101011100010010010000000101100010111001101100001011;
#1 $display("%b", po);
# 1  pi=207'b101000100111101000111001010000001010000000110100001001010100101101101110101010111101100010001000000110100001000000000110000001100010110010000100010100110001110101100101001111010101101110111111111010000000010;
#1 $display("%b", po);
# 1  pi=207'b001001001000111100001111101110010100111101010111000011001110100101100100010111100100001011111001111111110110110110001101110110001001010110001111111100011101111011100001011111111101011101001011100111101010000;
#1 $display("%b", po);
# 1  pi=207'b000101010010011011001111111111110100000011011001001001100011001001110010100111110011010110000100101101001011101000000110100000010101011100000001111011101100010100101100011101010100111110100100010010001100100;
#1 $display("%b", po);
# 1  pi=207'b110010010011100010011011000111001000111010111010011000100111010011100111001111101100001100001111011101000001011101010011010001100001011001111111010101101110110110000111101101011101110010100011110100111100111;
#1 $display("%b", po);
# 1  pi=207'b111101111101001101111010101001000001011010100110110000000011000111101001011110001010010101000101000101110000111000101001111110110001001001001100000111111001010111010101111110110011111101101101011000010110110;
#1 $display("%b", po);
# 1  pi=207'b010111111011010010100001000010001111000001101001010101011010111110111010010111111101011101010100100101001001101111011101101101111110000000110001001010110011001000100101000001111010101100110100110010011010011;
#1 $display("%b", po);
# 1  pi=207'b100011010100010001111101101001111100101001111000111101000110100001000111001110011010001110010101110101010111101111001000100100100101110110111001011111101101001011000001000101000000101110110110011011100001111;
#1 $display("%b", po);
# 1  pi=207'b101000000011011100111100011101111110100110001100001011010100011101001001010000111000110011011100111001100110011010011100010100001000110110010111101110001010100000110100010010010000001110101000101111001011001;
#1 $display("%b", po);
# 1  pi=207'b110110100100111011110010100110101101001000010001100000100011100010000111110011011111000101101001110000111011101101000000011101001000011101111101101011100010101110101010011100110110110001011010100000001110101;
#1 $display("%b", po);
# 1  pi=207'b001101100000001010111110001011010111100001001001000110100011011000011100010101010100000100000010011010110011110000111011101000101011010101001010000010100110000111100010110110010010000010101011001110000110010;
#1 $display("%b", po);
# 1  pi=207'b001011111010000010110111000010000011111100000000101110010100010011101010110011110001011011001011100100110110101111111111101001110011101011010111110011111011001001001101010010010001000111000100011100011011100;
#1 $display("%b", po);
# 1  pi=207'b100010000101000010101001100111110101100110100101110101110100010111011000110110010001111000010110101000111011110011101101011110100001000111001010001110110011000111010010101000010011000000001110111001111001100;
#1 $display("%b", po);
# 1  pi=207'b011010000010100101111010001010111011011100001110001001001001111000000000001011101010101011000010111100000100011101000001001000110111101111011110111001000111111011011110010011100111011001110001100100010110001;
#1 $display("%b", po);
# 1  pi=207'b110000010101110100001011011000001110110011010101011110010010001111001100011001011100111111000000011001001000011000010000100000110001100110110001110001110000111100001100111111001000001100100010100110001100001;
#1 $display("%b", po);
# 1  pi=207'b001000001100011101110001100010000100111111010100000011111001111000101010001001100111101011000000001101110101101011111000110110111001011110010101001001010111010101001011011001111101110010000010010101000101111;
#1 $display("%b", po);
# 1  pi=207'b101011100111111111000000110000000111010110100110100100011010111010111011001110101010110011101001010110100111000001001000100111000011000100001110110111101101010000101001000101000110111110111110101010010101001;
#1 $display("%b", po);
# 1  pi=207'b101110010000010011010000110000111101101100010101110010010011111111001010100010010010000000010101010000001111100000001100000100011011110100110100111110100001001100010101011011111101000110011110100010100100011;
#1 $display("%b", po);
# 1  pi=207'b111001100001001000100111101001000101010001010110001111101011010001001111011011011010010010111100010111001001011110111101111101110001110111010110110111111011100001000001100111000000111110001100110101011001101;
#1 $display("%b", po);
# 1  pi=207'b100001011111011101101100100101101110111011010111110101100110010011000100100011001110110110010110001100000011011110000100110001101111001000010101010000101110100100100101000010100000000011001001101010111100100;
#1 $display("%b", po);
# 1  pi=207'b101011001000000101010110011000110000111011001010100001100101101000010000010010001000000000010011101100010101011110001011000110000110100011001001100100110011101010011100001111011101101101010011011110101111010;
#1 $display("%b", po);
# 1  pi=207'b100010101010100111011000000100110010100100001000101000111001001111011001110101110110000111000011111001001110100101000110000111101110000000100011000000100100101101000101101101101110101100011101011110010011001;
#1 $display("%b", po);
# 1  pi=207'b011011100011011110110000100101101001001000011101110011100100100111101000011001000011111111011011000111110100011111110111100101101111100100011010110011001100011101001011110001100001000001010010010110000001001;
#1 $display("%b", po);
# 1  pi=207'b101101100101101101000111010100110111010011110000000000010100100100111010011011001011101111011011011111111101011010101101001111000111001101000111000010100110101011110001010111011001010111010101001010010101101;
#1 $display("%b", po);
# 1  pi=207'b001001011000101001100101001111000110000010000001001110111100011011010010001111010100100101001100001011111101000011001001001011000111100011011001001101111111101011011000010100110111111110001010111000100001111;
#1 $display("%b", po);
# 1  pi=207'b110101011010011100010011111010011101011001110011100010101000101001001010011000100110101100011101101111101110001000111010100000100000101000000110001110010101101000010001010010000011001101000000010011101111111;
#1 $display("%b", po);
# 1  pi=207'b001101001100100010101011111010000100110101101010010110110100011101010110101101010010111110010001111011100001110001001001110011101000100001111111000010011010011011101011100110011110101101110111111011000011011;
#1 $display("%b", po);
# 1  pi=207'b100110001100110101010010110110100101110111111011100000010000101000000010111100110101000011000110111001010011110111000011111101111101111000011010010011101100100010000110011100010011110111101110111101111110011;
#1 $display("%b", po);
# 1  pi=207'b011100010011011100101111001111001111010011011011000100010010100100001011111011111000100101111001111100010000110100001101011010000100111000101110010111000101110101110001010011011010110001100010111101010101010;
#1 $display("%b", po);
# 1  pi=207'b001100110111110110011110100110111110000011101001000110000111011110010001010001111101011111100110100101101100111010100100011011000001111100101010101000111100110110111111110010010001001001011000010011110110100;
#1 $display("%b", po);
# 1  pi=207'b100011000011101001100000010011110011110101111101011110110100010100000000011111100111101000001011011010111011001010001111101101110101101111111001001111100110011011101011110111111110001010111111011111001101010;
#1 $display("%b", po);
# 1  pi=207'b011001110101000100110001010001100011000010100010001101000100000000100011011011101111111010001010000100000100000010010101001011110000000100100100001001011001101110010101110001001011011000100101110101010100101;
#1 $display("%b", po);
# 1  pi=207'b100001010010111111011011110110001001011100011010100100000000010011011110000101000000110101100110011011011110010000010110111001001010011100111000011000001100010111111010110110011000011010101111100100110010010;
#1 $display("%b", po);
# 1  pi=207'b001100101110000101111010000010110001100100101110010011111011001000100001000110011000010101110100100111101110111010010110110000010100010011000111001010010011111111011000010111001110110100000000011001000001010;
#1 $display("%b", po);
# 1  pi=207'b100101010100110011101101010010101000111000111110111001010011110011110011001010101011111011001101111101011111100111101011000001110010011101000000110010010000000010010111000111010110101010010100100110000100010;
#1 $display("%b", po);
# 1  pi=207'b001110000011111110010110110100100010110011111011001100101001011100001101010101110101000010010000000010101011100111011110110001000001010100000111010100000110010001010110100111000001011011111011110000010001011;
#1 $display("%b", po);
# 1  pi=207'b111101001110101010110000010100001111001010100001010101110110000000010100011010111011100001010010001011110111000001010000011011101011001001010010010110011000110011000101011010111011100011001100010101000000110;
#1 $display("%b", po);
# 1  pi=207'b111101100001001011001100100000110010101101101010110000100000101110011111101010011010010000111101000011001000101110001001010001000110100110010101000010011011000001000000101010100000100011100010110101011101110;
#1 $display("%b", po);
# 1  pi=207'b110100000100000001110101000101011000001001010101100100100100111110011010100011101000100110011011000000111010110101100011011110001000111001011000110010011110100100011001100000101010011100011000111011100011111;
#1 $display("%b", po);
# 1  pi=207'b110110001100001101101001001110011011100100001100110110101111001111010000100101010100010111001001011111100110010000001001110101101010000101111101010000111000110000010101110000010001100110100111110101101110000;
#1 $display("%b", po);
# 1  pi=207'b100100101100011111101001010000000011110010101100110010110011101001100001110100111010100101011000001110000110100000101011011111001010111101000100101010011010100000000010000101000011110001100101110001110110101;
#1 $display("%b", po);
# 1  pi=207'b000100010001110101111011010010111011001110110111111001110010001100011100000001001100001010110110011011010010100001101001101001000100000100101100001101111100011100011011111011101001111000111010100011001110100;
#1 $display("%b", po);
# 1  pi=207'b010011101001011110111011000110101010110010000010011111110000000000011010100000000101101101100000010100001110110101001100111101101011011011111101110000001100010101001101001101000110000101011101010000010010101;
#1 $display("%b", po);
# 1  pi=207'b000011110111111010101111100000111100110110011110000010111100101100100000011110010101010111011110010011011111000111011010101001100111111111010110111001101011101101101100101101000011110000011111010011101110011;
#1 $display("%b", po);
# 1  pi=207'b111100111010000100101100001000011100011000001100101100011111100110000011010111011100010000111001000001100001001101010010000101010000011110011001111111000000000110100000011101101010110101101111111100110001001;
#1 $display("%b", po);
# 1  pi=207'b101000011111011001111101001001011101101111010011110001001101000111110101101110000011100011111000010111000110000100000110110111001011001110110101001110100010011110111001110100111101000100111000110000111100100;
#1 $display("%b", po);
# 1  pi=207'b000100110111011001101101000101000001010000011001010111000100010100001110100111011110011010111001001110111001010110100101111110000011000001100101111101011100100110111111010111010011100110001011101001101000101;
#1 $display("%b", po);
# 1  pi=207'b000100101000011011100000010001110001100000101000100111001110110110111111111010101111111100100101010010110000110001100000000001100111110101111101111101101000111100110011011100001111000011111110000101100111011;
#1 $display("%b", po);
# 1  pi=207'b010011101010111000010111010110001100110000111010001100100110000011011010010010000100010111010000010110000100011101010101001010101011100011011000001010000010010001100011100011110000001101100010111011001100100;
#1 $display("%b", po);
# 1  pi=207'b010111010101010011100100101101001011101110001010000110111010101110010110101110010010110011010011001100001101110110100100011101100000011110011011111001111000010101110101111010000000100100111111000011010001101;
#1 $display("%b", po);
# 1  pi=207'b001001011101011010111110010110010010110010010110101111100111100000101011101001111101011010011100100000101011000100011100110111101001010111100100000000010111010101010110111111110010010101111001100000100011001;
#1 $display("%b", po);
# 1  pi=207'b110111100111100100001010100011010100011001011111101010110101011101110101011111010000000001100111000000100000011100011000011110111000011101100010111010001110100110010101110100110000101110010010101111110100001;
#1 $display("%b", po);
# 1  pi=207'b111100001010011010110100011011010010100011101011001101001100101101101100001101100000110100011100111101010001100100000101111001001011000001111000110100000111001101010110101110001111010001010000100110001011001;
#1 $display("%b", po);
# 1  pi=207'b010111010100110001010101000100101001100110100100110001110001100011010000011100001101110111101100101010001110100100110000111110011000000000000101110010101000010011011100011100001111000111100011001111000000011;
#1 $display("%b", po);
# 1  pi=207'b000001100100111000001111010011110101101000111111010010000001100110000000011011010001101100000101100010000001101100000110100101000001000101011110011001000000011110010011001010111100001110100011000110101111111;
#1 $display("%b", po);
# 1  pi=207'b010111010100000110101110010101011011011000010111000000010000101011101100011010100111100010100001011000001001101110000111010011001110101001001111110111010011010101110110010111111000101100111010111011101111000;
#1 $display("%b", po);
# 1  pi=207'b000010000111000001110101110101000111000011001010101010101100101111100101000000001101100100000101111101111001000110110101110001101010000010001010011111100000110101111111111111011000001100011111100110000010111;
#1 $display("%b", po);
# 1  pi=207'b010100000001100000111010011010000110111011100011000011101000100011001001001110000110111010101111111100000010000101000101110111000000101010011000101101110010010101010000001011000000010000110000000010000000011;
#1 $display("%b", po);
# 1  pi=207'b100000100101100111101010111010110110000010011100011110001010001000100001110110000010111110101011011111100101110110000000110010111101001110011000100100100001000111101100101111000111111101111100110110000010100;
#1 $display("%b", po);
# 1  pi=207'b000111101100101011010111010101011110101010100101110100101000110111011101111100111100011100110100000000010000111010100001111010001100110100101100110100101001010110110011010000101000111000100100101111101101010;
#1 $display("%b", po);
# 1  pi=207'b011111111101111011100100010101010100111101011011100000011000010010111011111011010000011111000101111000010101100001001111010010101000011000010010100100001101010110101110101000111011111101101001111010111110110;
#1 $display("%b", po);
# 1  pi=207'b000000010010110100011110000100101010101001100100011111100011110110100101000100111000011011111111011101011001100000111100100100110100000000111001100001100101100000111010101011100001111101011111100011100010000;
#1 $display("%b", po);
# 1  pi=207'b101101100110011111001000011101000000001001011010100100101010000100110010000100100101011111011001101010000110010110010001111111000101010110111110001000111110010010111010110110110110101001111001101001010101010;
#1 $display("%b", po);
# 1  pi=207'b110111001111111111001011100010000100110101110001011011011010001000011000111101111010111001101100011111110001100010101001010101101111001001110111101001011010010100011111100101001111000010111101111010001110111;
#1 $display("%b", po);
# 1  pi=207'b010110101011001111100001001101101100010111100010111110001111001011110111100111000011010111001111100111000111010100110101111111110001100011110100100000110001101000000010000100001000101010011010101000101100010;
#1 $display("%b", po);
# 1  pi=207'b111101111100100111010010010110110001001110100111100111001001000011010101101110000010010000111101110010000011010011100101100100101111011111100100001111000100001101011111000011110100010100101000001111101001000;
#1 $display("%b", po);
# 1  pi=207'b010101111110101011100110101001110000111100100111011001110011001111011100100011011100001101011100111110111110100011100001011010000000000101100000010010111111000010111101000101011110101001010110000110100011111;
#1 $display("%b", po);
# 1  pi=207'b000101101100111001100011101001101011110000000110101111110010010000011101010001100101100110100110000110110101011111111001111000101011110001101011101000100100011111101100101001111010101101110011001010111011100;
#1 $display("%b", po);
# 1  pi=207'b100111111101000000111111100111001100111010010001000000101100001100110011111110111011101011001010110110000101100001000111010010000101010010001100010100101011101101101101011000100110100000110000001101011110000;
#1 $display("%b", po);
# 1  pi=207'b100110001111001010100001001010101111101101101100111010001000011000000010000010001110010111001110000100000100000011011100000011101000000110100111101101001110000110110001010100000110001011100011011110101101010;
#1 $display("%b", po);
# 1  pi=207'b000011101100010011011011001110010001011001011001100011110111110000100001100101100111001111010000100110110111000001110110111100100000010010000111010000100100101101100111010100100110001000001010001010101101011;
#1 $display("%b", po);
# 1  pi=207'b011001001011010000101100111100001001011100110011100010011101001111110100001111001100101100100111000011010011010100000011110100100110011101001111010110101000101011010100011000000100011111111000010110011000101;
#1 $display("%b", po);
# 1  pi=207'b010010011000101000111001110001011011001001010000110110001100100011001010010110001000000101111001110011101000101001111001010010111110101010110101010101001000010010110100010100010101111010010111101000000011010;
#1 $display("%b", po);
# 1  pi=207'b001100110011001011100111100111101001100000011011100010100110100100100110010111011111010000111111001100101110100000000100010000110111110000100110010000101001000110010100100110001101001100010000000011001000111;
#1 $display("%b", po);
# 1  pi=207'b001000001111110111111101100010000010001011000110010010001100101011001001000001011001011000011001001011111000001100111011001100111101110101011010101001001011101101110110001110011010011100001100011010111111001;
#1 $display("%b", po);
# 1  pi=207'b001110000101001011001100110110111000110101111000100110101101110011000010101001011110110011110000100000100010111001100010001111101010001001101011010111010110011100100100001101010010100110010010110000110100100;
#1 $display("%b", po);
# 1  pi=207'b111001110111100101100101001111101000000010110010111000010110000000100110100011110110000110110111111010110100110000100101000000011011000101101011101011010011000110011111101001111110000001001011001011110011001;
#1 $display("%b", po);
# 1  pi=207'b001001110001001011011100110110111111001111100111111110111000100100010010110000000001001010001100001101001001011111101000111001110110100100011111111011011100011010100110011011100100101010001101010010110011011;
#1 $display("%b", po);
# 1  pi=207'b011101011100110000011010010010010111001100001000000001110101010101011100000110011000000100010101101101011010000101101001010111001111111010100011110001101000101001010001010100011100110010110001000000100110110;
#1 $display("%b", po);
# 1  pi=207'b100100001101001101100001101001101110111110101100001000011100011001111011011110100110101101110110110000010111011110011001111010001011010010100000001110110000001110011100011111101011011100010100001011100111001;
#1 $display("%b", po);
# 1  pi=207'b001111100000110001100111100000110111011111000100001001111110110111110110001110101100100110000011100110000010101110010010100110010010110110011001010010101001010011111000010101010111111100110010100100010110111;
#1 $display("%b", po);
# 1  pi=207'b101010001101010001110110001011101111111101011010100010100110001010100100110001101111101011010111111111101001011001111001101010100111110100100100101100011100101110111011001110010000001110110100011101100011111;
#1 $display("%b", po);
# 1  pi=207'b001100011001110011110010011101100010101010011111001011100010110001110000010010001000111000011100010111101111011000111111111111001110000000000111000011110011000001101001000100110000101011010101111110100000000;
#1 $display("%b", po);
# 1  pi=207'b001011000110010010111011001110100110010101110000011100011110010010111110010101000010110000100001001001101010101100101010001010001000110011010100001100010010101111100010010111000110010110100011001000100100000;
#1 $display("%b", po);
# 1  pi=207'b101010001101000110101110110101110110110111110110101111001101000111110100000100011000101101101111000111110101010001010100100101110001101111111101000101110001110011110101101110101011111001010000001000111100110;
#1 $display("%b", po);
# 1  pi=207'b111011000001101011101101010010100010101000111000010111000110100001000100100010100100010110101001000101100010110001100101010000001110000011000100110110011001010101111110010100110001000000111010000001100101000;
#1 $display("%b", po);
# 1  pi=207'b010010101111111010010000000001011010110110100010100100110111111100000000110010100110111001010010010111010111110111100000010010011011110110000010001110001111101110100100111101110100001100100110100101111111100;
#1 $display("%b", po);
# 1  pi=207'b100001010011100101010100110000011000111100101100001110110111101010010010110001100111011000101000000100000011100010011111001110101010101111111111011011110001011100110100011100001010100101011010010010011010110;
#1 $display("%b", po);
# 1  pi=207'b110100100111001100100001111001110101111010101011101010010011110001001010001011000010100000110011110110011111010000101001010011001100000011001011101010001101010011110010010000011110011010111010100001110111110;
#1 $display("%b", po);
# 1  pi=207'b000111100000001100010001000001011111111001101010111011100110000010110110000010001110101011001100010111110110010010101011110101001110110010101111001110101100110110010100000000011000110000010000100111001110101;
#1 $display("%b", po);
# 1  pi=207'b101111011000110010001100110101010101110100000110010101100010010111111110011011011000010111000111000001000101101000001010010000110001001101011010101000011110101101110001001011110110100101101011111100111101011;
#1 $display("%b", po);
# 1  pi=207'b100011010011100001001101011101000001101011001101000010100101100100111111011010111100011010100111100100101010010101000000001111010010001001000101101111000001111011000001100011010010010101101001100001001101000;
#1 $display("%b", po);
# 1  pi=207'b101110011100010100001110010100010111011001000011101111111010101000111101000000101001001001101001001011000111101110001000000001100000100111101110011101110101010000001010000100111110101101001100101001110100000;
#1 $display("%b", po);
# 1  pi=207'b110111110101100010101010010001111110101000011101111110111110100100110001110001100111001110111100110011100111100111111101101110011010010010110000110100111101011110001111000101100001110111011011110000010100110;
#1 $display("%b", po);
# 1  pi=207'b011101111100010110010011001100110100000110110010010011000111000100001111001011010010010110010011110000111001010001000111010000100000100100111111100101100100100111011111110011001000000110001100010111011101111;
#1 $display("%b", po);
# 1  pi=207'b011100101001101110101101011010001001110010111010011100010001111011001100000000110111010011000110101100100100111101101110011101101011011110111000011000110101110110101100000001111011101110110000110000001000100;
#1 $display("%b", po);
# 1  pi=207'b100000110001000100011100010010010011100111001010000100100011010011110101101111000110001001010010000001110100101110110001011001111010101010110111001000100001101011000011000101101101111001010001011010010101010;
#1 $display("%b", po);
# 1  pi=207'b101101100110001111110011110011010110011001010101101110001100100111110011000010011011011010000110011101001110001100010111001010100001011000011111001000100111111101010111101011100010100011001000010011011101101;
#1 $display("%b", po);
# 1  pi=207'b110000010101011000001011110111000001000010101110110011001101110001011110110000101011101101000010101000011101101000000010100111101100100011100110001011100100100010011110100010110010101001011001100110110110001;
#1 $display("%b", po);
# 1  pi=207'b011011000110001110100101110011110010011101000100101001110110010111000110101001001101011011100011100101101000010010000011001111110000011001000001100100011010100111001101010111010100011100111110110011110010000;
#1 $display("%b", po);
# 1  pi=207'b011101110111111110011001011010100001110111100001011000011110010111001101010100001011101011001001011000011100011110101011010000110011001010000111111110111110100101101011011110100110000011100111111100110011101;
#1 $display("%b", po);
# 1  pi=207'b100101010110111110111011010111111010111100000000100100000011011001101111101110111100110110111111111110011011101101010001110100111100111101010111111010101000111101000100100001100000100100111001000000100111101;
#1 $display("%b", po);
# 1  pi=207'b010001010010111101011000010101011110100101111010110011001111011001001011010011100000001010110110001110110001101100101101000100110010000100001000001100001111100111000111000110101001010001001110000001111010111;
#1 $display("%b", po);
# 1  pi=207'b111011000011000010000010000000011001011100100001001000000100101111110110011101011000010110111110111100000100100111100111111000110110100000011110001011110011001111111010011001110001000010000110001100110000100;
#1 $display("%b", po);
# 1  pi=207'b000101101100000101011010000011010101101110011011111000111001111011100011111100011000100110111010000000100101001000101101000001111010000011000000000001110010011000101000101110010110101110110101101110001111101;
#1 $display("%b", po);
# 1  pi=207'b001001001101010001000011011111110001111111000100001001100010101010010100110111011111100010100011001111101001100001000010111011010001101111110100000011001001100100001010000110001110100100010011000011110100000;
#1 $display("%b", po);
# 1  pi=207'b010111110001110101111110110100101000110110011100100000001010000000101110000001011101000100001100001111011101111110101010111110001101110100100001111011101110011111111001010000001001100001010010001000000000111;
#1 $display("%b", po);
# 1  pi=207'b111011111101011010100011001110101111101110011001101100100010000100011000101000001000001010110011111100010011100011110001110001011111101001010010110110001111001110000100000111011001010000101101100011011111010;
#1 $display("%b", po);
# 1  pi=207'b011010101110011101100001100100101001001100100000100110000000110100000101110010110111111001110111010011101000101000100010000111001001001101110000001101000011000010001100001011000110101010111100110011001100001;
#1 $display("%b", po);
# 1  pi=207'b111000111111001111000111100100111110100011101000000010001000001110001011100101111000010000001111100101000110000001100011000011011111110111010010111001010110000101110010110001110001000011101111001101101010111;
#1 $display("%b", po);
# 1  pi=207'b011000111100001111111001011010010010011001001100010111110001010010011011110011111010001011000000011001000001111101001001001101101110101000100101011010001000110011100011011010111110101011110001100101100101001;
#1 $display("%b", po);
# 1  pi=207'b001001001011110101000001000110110000100000000100011010101111101010110111001000110010100010010101110001100001010000111001000001000000011101001100010011000010000000101111111111110011011011101001010011011000010;
#1 $display("%b", po);
# 1  pi=207'b110101011100100000010001010101110001010111101110000010110000111101110011110000010000110111011100010101000010101011101010001110001000000010100001011101111101001110100011000011000011101001101110000011011001010;
#1 $display("%b", po);
# 1  pi=207'b111000011000100011001000110010101111101011011000111010111101011100101010011110100100010110101001110111001011100111111110001000010000000011001110111011110110000100010010011010010010000001111110111100110110010;
#1 $display("%b", po);
# 1  pi=207'b111001010111000010010111010000110111100100100001011011110001110011011100101111000010000000110110010111100110010011000101110111110101011001001010001100010111100011000111111100100010001011011001111100001010010;
#1 $display("%b", po);
# 1  pi=207'b111010010111101101000000000010101000010100110011011010010110000001010100001000010100111011001110111011100100010111000011111111110110000110110001101100010111110101111001101101101010000111001111001101111101100;
#1 $display("%b", po);
# 1  pi=207'b100001111110000011101101100001110101010000000110111000101110001111011111110110111111100101011110011011000101101111100110101101100011100000011001110011101000110101000011011111011110110110111110010000100100010;
#1 $display("%b", po);
# 1  pi=207'b010010010000011001111111111110100011000011011010110101101011011111111011101100000000110001100111110010110011011000101100001000100100000011000111110010110110001011111110100110111101100100000101000111011110010;
#1 $display("%b", po);
# 1  pi=207'b001010111101101111111010001111111000100100101010011101100100111101010011100111001111100001111100110101001100010011010001101101010011101111010101101000010100101111101001001111011011111011111010101111100100101;
#1 $display("%b", po);
# 1  pi=207'b101111110110101111110010110001100111100100001110010111010110010101000011001100010000001111010100100001001111011100011111100011011010001101100001101010011101001101000000001001111011001100100011001111010000001;
#1 $display("%b", po);
# 1  pi=207'b110011011001100111110001011000000101110101111011000101110110010001101001000010110000011110001001000110001000111110011110101100111101111010000010010111110001101111010000111111000011110100011111010111011001010;
#1 $display("%b", po);
# 1  pi=207'b100011100011011001110010010110110110001110001011111000000010110101100111011111111101100100010000001010010100101010111010111101111101100010001111010000011100010111110110001001010110001110010110000010110011101;
#1 $display("%b", po);
# 1  pi=207'b000001110101110010001000111111101111001010100011010100011010011001101010010100111110000101010001111101011000010101111000000101111001110100111110111010001111011011011000000101001111011110000100011010011001110;
#1 $display("%b", po);
# 1  pi=207'b100101010100001101110000101100100100010010011101111110100010101010011001011101100000100111100000001000011100001100011010011100011011100010000011100100011011110001001010110000000110101100001000110011001011100;
#1 $display("%b", po);
# 1  pi=207'b010000010001010110111111001111010000110001110001000111011101101111111111001100101010111000010001010110011111000111111000000101001001010100011000110101011000111001000110101001011010111100011100011010010000011;
#1 $display("%b", po);
# 1  pi=207'b010001101000110001101010011010000000000110001101010101101100101100100000111001001110100101010101001111011001011001011110101111111100101010100111111011000000010001100100110110000100001111001001101101100001000;
#1 $display("%b", po);
# 1  pi=207'b110001111000011010001011110111110001100010110110101101111101101101010001011110101101001100101010000101101010001111000001010000010011010011111100101110100000100111110100001110011101101011111100100100101010110;
#1 $display("%b", po);
# 1  pi=207'b000001110011000000001110110000101011101000000110000010001001000111010010111101001100101011101100100100111010011111010111011010011011010110111010111101000001100010011100010111000001001101010011110010001011111;
#1 $display("%b", po);
# 1  pi=207'b111001110101011100100000010110100100101100000100010111000100111110011110001001001100111110111111110110010010000101010100100101101010100110100001011001010100100110011001101001001101110000100110000000010011100;
#1 $display("%b", po);
# 1  pi=207'b100011111001111110111101000101011110001010101001110111011110100100111100100000111001000111110010001011100110111101011111000001111110001110111000011111011110001010101001010000000111101100111000101101111000111;
#1 $display("%b", po);
# 1  pi=207'b110111110011101000111110110000101100110110001100011111001111110011010101100101111001110110010100110001010011011011111111111011001111010100100101111001010010110011010100010100111101000011100111001011110001111;
#1 $display("%b", po);
# 1  pi=207'b001100000111101110110101000001101011010011101110111000001011011100111000010101111001111100000001110111000100011000010111010110011010101111101111000100110001001011110101101100101010001100101101011100110110101;
#1 $display("%b", po);
# 1  pi=207'b101110101011010000101000011110100011010000000010111011100100100100110000100100111111101000000000011001010001101001100101001111110101010001100100101101110000101110111011100001101100101110100101010100111110000;
#1 $display("%b", po);
# 1  pi=207'b010111001000001111010110001000110010001111010010111010100011101011110000001000100000110010011111110110000100010110001011101101100110110010100010100100011110100111000110010001101011011111100001000111101101110;
#1 $display("%b", po);
# 1  pi=207'b110001111111110100001110111001010110110100110011110101100011111111100001001110100101001111001010010010010011010101110110111010001011011110011001001100101111101011000010111011010101111011001100100101110000010;
#1 $display("%b", po);
# 1  pi=207'b101000110111010111011011000110101010100001111000011000101001110011110001000000010011011111100100010001110000001000010000101011010101000011101000010111101101001101001000000001101010010011010011110101110101000;
#1 $display("%b", po);
# 1  pi=207'b101110001101100011010100101111010001001001101100100011001101000110110000000001101011001100100100111001010110010100110011001111000010110100101000111000011000001010001101000111000111000100111001101001101110101;
#1 $display("%b", po);
# 1  pi=207'b110011111010001110011101000010000001111001000100101000100010100011110010101001100110101011110111100000000110000100001110010010100111000011101110000100010011101011100000000110110110110000101001101000110100000;
#1 $display("%b", po);
# 1  pi=207'b001110011011101111110011100100010101010001111101001000011100001100110001011001101001000100110011110000011000000111110101100010000111001001011100100111011101001110110011111100001010000111000011001010100111111;
#1 $display("%b", po);
# 1  pi=207'b001011111110011001010010001011110101101011010001011110001100110000011101001010000000111010010111100110101101110011001010111100111010010001111010001110000111111110011110011111101010010111000100010110101000100;
#1 $display("%b", po);
# 1  pi=207'b100100101011101000110001101111110000111110111110010001000011111001001100100010011101001101100011010110101000100101110100101101100011110111010010011111000111011111111000011110111110111000101010111100110011101;
#1 $display("%b", po);
# 1  pi=207'b011001001110111010001100111111000101110110000000111010110011010110110101011110001011101011010101111010110101100010011100001011110010010101111001111110101000011010000011100000110110100001000100001011100000000;
#1 $display("%b", po);
# 1  pi=207'b100101011110111000111110001011011101111001001000101101001000100011001101101001101101111111011001110110100110001111000101001100011111000100011011000011001000110011010011111101110101101111110100000100111101011;
#1 $display("%b", po);
# 1  pi=207'b110011000110111001001110111101110011100001011001111010110111000111100111011110101111111011010010001111001101011011100101011101100110000111110111111010000011101110111011110010100011100111110110110000001011100;
#1 $display("%b", po);
# 1  pi=207'b111110111001111010100000001000100111010111101110111101000001100110000111101111111000100001000001000010001011010100110011011001000000011110110101000001101010000110110100101011101110101110011010000000000111110;
#1 $display("%b", po);
# 1  pi=207'b001011110000100111011110011000011101100000001111001110001010001000001110111100001010011110000110111010100111011011101110101111100110000111101110110000001010100011000110110111010011010101110110101101100100010;
#1 $display("%b", po);
# 1  pi=207'b001111101010001001100110101001100111010100101100010110000111001100101101010001111000100101100001100001110111010111000010100101000100010000101111000100111110110110000000100000100101011110001000101110110111010;
#1 $display("%b", po);
# 1  pi=207'b100110010100101001110111010000100100011110011110101001001110011111010101010011110010101010000010101111111110001101110010101100001101000001111100011111001000100000001100010011001100100101010010111001000111010;
#1 $display("%b", po);
# 1  pi=207'b010011011110100110010101011101000011101001011101110110010101011000001010111101000110001000101010111011000010111111000011010100111101000100000001001111101011011100000001111111111010010111001010101010101110110;
#1 $display("%b", po);
# 1  pi=207'b001001111011101011010011010000011001000001001010011101001100011010111011000011100011011001110100100110000001001111000010101110001010110011010100010101010100000100101111010101110111000100111110001011011111010;
#1 $display("%b", po);
# 1  pi=207'b010110110101100000110101100100111010100100010111010011011111100110101110001100011000011100110011001001001011110100011010001111000111111011000010111100100100011110010101001110101001110110010011110100001001000;
#1 $display("%b", po);
# 1  pi=207'b010010110011011000011111110011010101101110110100100100001011001101011110110001101101011111100111101111011011100000010100101011001111100100110000001011111010101111001001101100111100001110100100010101100010110;
#1 $display("%b", po);
# 1  pi=207'b111000110100101011011111000010000000001010101101111010010000111010010011011010110101111000001010011111010010100010111000010011001011111000110110100011101101011000101011010000110010001100111100001010010011110;
#1 $display("%b", po);
# 1  pi=207'b111011010011101001111011111000110101001111101001000010111101110111111000001010011101111001011011011111100000111100100100111100111001100010101000001110110100001110101101101101010101000001111011110011110110000;
#1 $display("%b", po);
# 1  pi=207'b110010001011010001100011101011101100100011110010011100110001111011000101110010000000101100100001010110111001000010111110001110001011010001011001010000101111000100010011110000111000101111011000000100101011000;
#1 $display("%b", po);
# 1  pi=207'b110000010001011111110001000011110100000010010110011110010001011011100111011011100010110110100101110000010010010111011000000000111110100110001011110010001111011010110010101000001110001100001100001111110010011;
#1 $display("%b", po);
# 1  pi=207'b110101001000001001001000111011011100001100110100100000011110101100011010101100000010101001111000100001111011011001001101111011011110100001000101110101000100111100001011100110010101101110010010001011100110110;
#1 $display("%b", po);
# 1  pi=207'b011110000000101010001101010010100110100100010100000011100111011110000110101000100010110001011011111101101110000110001101011010011001001001101110001111011010101011100000011101111001001010111100100111101100101;
#1 $display("%b", po);
# 1  pi=207'b110010100111010101010100001011100100100011001100111111011011110010110110110101000110100010111011001111100010101010000101011110000000000111011111011100100100100000010000011001111110111101110000110010110010000;
#1 $display("%b", po);
# 1  pi=207'b011110101100100111011001111000100011100011010110100011100010001001001010100110010101110001011011110110011011110000111100100011011110100010111111101010101111101101110010101010001110010010110010110100000101110;
#1 $display("%b", po);
# 1  pi=207'b101010110110111111000000000101011011111011011111011110001010010011010110100000000100010110100010011110001110101001000110010110100000111110000001100100110110110011010011111101011010000010101001100000001010101;
#1 $display("%b", po);
# 1  pi=207'b000111000010100001111001000001011111110110111010000011100010111000011110101001101110011100011110100000010011100110011101100100110101101000011100010101010000111111001110100100001011100001101000100010000111110;
#1 $display("%b", po);
# 1  pi=207'b100111100111011000011001010110011101100100101110001111010011100110000011000010101110101000010010100010000011011100000010011000011010000100000000110000001011010101011010001110011101111001100010001110100001000;
#1 $display("%b", po);
# 1  pi=207'b101011101000011001010111110010001111011001001101110100010101111111111001000001011010011111011010000000100111001110101011000001111000011010110010000001000100111000100110011100001011011111110100101111001001011;
#1 $display("%b", po);
# 1  pi=207'b000100000011011011101000011010110000011000011110010010111000111010011011001110101100011011001000101001100011001010111110111101100010000100101100001000010111000111011110101101001001001110001011101111111110000;
#1 $display("%b", po);
# 1  pi=207'b011010000000010000101100101001111110010101001110001101010110000011111111100101010000000100101000010000110001110011010010101000010110011010001100010101000100101101111101101000100000111001011001001101101001000;
#1 $display("%b", po);
# 1  pi=207'b110100101000101101000111101100101000100101100111001100010001100110100011000010110101001001111110100010010011100101000010001011111101100010010011000111010101011011100100010110001110111000100011111110011110111;
#1 $display("%b", po);
# 1  pi=207'b101111100010101111000001101000011010010101101111000111110010011001101000001001101110011011101101000011111110001101010101101011110010010111001100000100000111010000111110111111010110001011101100010111110000101;
#1 $display("%b", po);
# 1  pi=207'b111010010001101011010001011001000001011001001000111110110101110010010001011100110101110010111000101101001011111110110100110010110001001011000001011011101100101110110101110101010100100000100010110111001110001;
#1 $display("%b", po);
# 1  pi=207'b111110101110011010001000010111111000101001100101111100110100010010011001011111110110101101110010101001000101101001010000000010100010111111101000010111110010111001010111100100101110111010010101110001100011011;
#1 $display("%b", po);
# 1  pi=207'b110111000011010100010001101101101111000101011100111001011101111001001110001001001110100000011011011000011101100001101011100001110110110101111000100011000010011110001110000011011001100110110111011110101001001;
#1 $display("%b", po);
# 1  pi=207'b011001000110001101000011000101000001110001100011111000100110111100100101011011000111010100111101010111010101101000111110011101100011110001110001011111001011110011011111000011110001100000110010010001110110101;
#1 $display("%b", po);
# 1  pi=207'b000101001111010110110101110111001010100101101111110110001000100101101110010100000100111110000000100101111001111000001010011011000001111100001111000110110110001011110010111100001001011111000001110000100100011;
#1 $display("%b", po);
# 1  pi=207'b101111011111100101110011001010010110011101111100110111101100010101010010101101101011000111110000101100110111100011000111100100101001000010011101001011011111001111110011101110010001010111001101010111011000111;
#1 $display("%b", po);
# 1  pi=207'b111000101100000100000011110010001011100011100100001011010011101100000110001111010000100000110001111000111010101111100100100111101101100000110110010011111101010000110100010101011010001010110111101010101011100;
#1 $display("%b", po);
# 1  pi=207'b101011010011100110111111110001100101010011001111101001110010110100000001110001111001101001000111101100010011100001010010001011001010011101111101110111000011000110001111111100000010101000111000100000010010010;
#1 $display("%b", po);
# 1  pi=207'b101111010101111000010011011110000010101000010010001001110111010101011011110101000001000111100111110111110100100111100110101010011110001000100100110110001000001101111100001111110111000010100000000111001000000;
#1 $display("%b", po);
# 1  pi=207'b010101001100000101110100101011010100110000110011011010110011110001111101101100111001010100110001100011010100101010101011100111001010010010100001110110100110010010110010010101100111001001100000011001101001101;
#1 $display("%b", po);
# 1  pi=207'b101100011101010110101101101011011110110101111101111101001001011110001010101101001001100100011100011110011100111001011100101101110100001000100011110011111111110010011010010001000011011110000011011111010010000;
#1 $display("%b", po);
# 1  pi=207'b001101111000000000100000100100001001110101101000110011001110110010000100101100001011001011100010001011111000111100111001111011011100011001110111010100110011110011111001101111100100011100000100011000011010101;
#1 $display("%b", po);
# 1  pi=207'b111000110110101011111010010110100000000100110111000000111010001101011011100010011110001001111111111100111000001000001001100011101011011011100101010110110101101110101001110100100001001110000011101111101010011;
#1 $display("%b", po);
# 1  pi=207'b111110111001010000100010000001110101110011110110011110110100100110000100110001010101000110101010011101101101011001111000101111100010000011000110101111010100101101110100000001101010000010001001111011000101010;
#1 $display("%b", po);
# 1  pi=207'b111010110111111011110011110111010100100111100100010100001000010111001010010110100101010010111110110100010101001001110010100101100101110110100100101001111110101010001011011110101101111011100010100010110111000;
#1 $display("%b", po);
# 1  pi=207'b000011011010110001001110101101110111110100111111010011111111110011100010011111010001001111000001111001001010110100001010000011001101101011100001110001010111111011010110110001001011100001010110101000101001110;
#1 $display("%b", po);
# 1  pi=207'b101111001111110110000010100100000000101110101011101110110000111101010100011011010001100100100100110011011000010110011000011110110100011111010101101001100101010001001011010100010100011001100000001100110101011;
#1 $display("%b", po);
# 1  pi=207'b011000001101110011010100001010000100110000100000001100011101101011100100110000010011000101111010000111001100100111010000000110010111101011001110001100111000000101010000101100000000011001011100001011000000011;
#1 $display("%b", po);
# 1  pi=207'b100100000010000011011110000110111001001101100110100101011000111001100001010010111110001111111001110000000000110000001100101110101010111010110011001111100001000110100101000100101001011110011010101100111100110;
#1 $display("%b", po);
# 1  pi=207'b111100011001011110111101001000101111100010101010111101111000011010110001000000111100100111100001111001111000001000000011011100101111100100001101111010110101110100101001011111101000110111011110110101101101110;
#1 $display("%b", po);
# 1  pi=207'b101011010101110001111011010111011001100010000111001101100110110101001100110100100000000001001000100010100011010010100111011011000111100011111001001010010001000111111110010111101100100010111111100001001011100;
#1 $display("%b", po);
# 1  pi=207'b011100010010101111001001000011111010110100100111010010110111000000110011000110010001010001010001001001010001110100011011111100110101101100010100100010111110111101111101111111110001111100101101101001101010001;
#1 $display("%b", po);
# 1  pi=207'b101110101100100101001111001110100111101110100011000100110010010101110001001000110000101110110001001100010010011010100011001110010111110011100010100101000101010110110101011111101001101110101111101000111101110;
#1 $display("%b", po);
# 1  pi=207'b101001000001101000001010111010111100100010001100011110111101011111011101001101010001011001101110000001000010011010101110011111010101101011000101111111100000000101010001001100111110001010010100010000100101101;
#1 $display("%b", po);
# 1  pi=207'b111000000001001011110100100011000111001111110001001010011101101011100011010110101000101101110001000001101000011001110000000101010110001110111001101000000101100110100001010000111001100111001001100001111101000;
#1 $display("%b", po);
# 1  pi=207'b011011101101010011101110000101110111001001100000101001111111011110101000010111001000000100000101101101001110100111011100000000001000010110100011001111101100110001111000110000101101000110111110000011100001110;
#1 $display("%b", po);
# 1  pi=207'b101001000010100111110000011010000101101101001010100111001110110011101111101100011110111001110101111000110010111100011100011110111010000111001110100000010100011000110100100000110011001110011011000010111111001;
#1 $display("%b", po);
# 1  pi=207'b110001111100010101000100111101001000000001011100101111111010011111110101110001101010101010011001100010101000001100101000000010001100110011110111100000011110000001110010010110000010011111110101101011001000110;
#1 $display("%b", po);
# 1  pi=207'b110000110001100101010110001001011010000100011111100011111000110110000001011101111100111110011001101101110000111101110001001011110011001001000010010110010011100100101111000111010001001001010101001011101110011;
#1 $display("%b", po);
# 1  pi=207'b111010000000010100111000100100110001011111010001100010111001000111010010011011111010101011010001001010101100001010000100010010100001000011110010001000101100001110001011010001111100101100101110101000110100111;
#1 $display("%b", po);
# 1  pi=207'b001111110101100101111000101110010010000110010001000010010101000100010101101101010111011001000011100110110100100111110000110110100111111100110100001101000101110011101011111111111111100010111101000000011101111;
#1 $display("%b", po);
# 1  pi=207'b011100110110101011010000011101111111111001110101001001100101101110000000110111010000100011110111001101010010001101100001011011011010011101100010010101110100011000101101001100100111101000010100100011000000000;
#1 $display("%b", po);
# 1  pi=207'b010111110000100000001001110000100101000011000010110111010001011110110111111100101011010010000110011110001001101101001011010111010110000100111111100100110110000001001101100011000011111101110110010110100010111;
#1 $display("%b", po);
# 1  pi=207'b101110011111011111110010100110111100000110000000011010101000001110101011111000101010001011100110101100010001000110101001100111100010011001100110100100010111100010111101000100100100000110100000011001110010010;
#1 $display("%b", po);
# 1  pi=207'b111011110010001000111100110010101110001000101001000000111110100001111110101001001010000010011010001111011111110010010110011001100101010111111101110101001101001110100010101100000101111110111000111011010010100;
#1 $display("%b", po);
# 1  pi=207'b110100010101110111010011101010100111101100101101010111010101001001011100100001001111111111010100010110101110111010010011001010001100001111010001011110110010111000010100000101000100100010101001011111101010110;
#1 $display("%b", po);
# 1  pi=207'b000011001010001110100111100000111110111101000011000111000010001111000010010111111100110011111011101110000000011010100010101101110011101111101011000010010111100001101000010110111001110000010000010110010111010;
#1 $display("%b", po);
# 1  pi=207'b110100111101111101111001100010001001100001101010101100111011001101111101001000010100001000010101000001011010100101111101101010111110110101111000100101011111101101000101000001001100111110001110110000000101101;
#1 $display("%b", po);
# 1  pi=207'b101101000011000000010011010110000011000111000100110100110100000011010100111101000000100111110010010010110100100110000000110100000110110000100101000000000000001110101110010110110101010111010110010111111001101;
#1 $display("%b", po);
# 1  pi=207'b001111101100010001100001100010011000111100111111101001111110010011110100100110010101101000000011001001101100001100101000010100001010001001000100101111100101011010100110011000101100111110111101100111100010010;
#1 $display("%b", po);
# 1  pi=207'b010110101100000111010101100010111110110000001011011001001000111111001010101010001101010010010110111110101111101011100110010100011110001011101010001111111100011101000011100010001000101101110111010111010001111;
#1 $display("%b", po);
# 1  pi=207'b010001001001101010011100100101101110100100101000110010101000000001000100000001000110010011000010100111100001100011100001010011111011010010111001100010101010100001000100100111001110001100100111010010110101111;
#1 $display("%b", po);
# 1  pi=207'b001000001101000101010110000111000010011011011001001011000001000100110110110100111110000011100101001101001101100010111110101101110111100100101010111000001011101101000111111011011100001111001110001010001011100;
#1 $display("%b", po);
# 1  pi=207'b011001110001011000111111111010100000111111000110000101001011010010000111011101010110100101011011101000101001001011000010111010100101001000111010000100000001010111110110101101010101110100001010110001111111110;
#1 $display("%b", po);
# 1  pi=207'b100000111101011110010110110011100111010000101001111100001001001011101100110110111110110110011111110011111110011001001111100110110000101001011100110010001101101101110100101011110100111011011011010101001001111;
#1 $display("%b", po);
# 1  pi=207'b010110101000111110000001110010101111111011001110001111000010100000111110000111111001101100011001001010101011011000001011000001000011010111011100101001011011010010101101111110101101110000100100101110001010100;
#1 $display("%b", po);
# 1  pi=207'b100110010000110100111101011110110100111110110101000101111001110101011100110011100100101001001010011100011001010110010000011110101001010101001101010011101011110111100110100111100111100000110101110111011010110;
#1 $display("%b", po);
# 1  pi=207'b111001000110011111000000010110000000011000101101001000011111010101111100010111110011000011100001110000100101010010001110101101011101010110101001001010000000000000010000010010010010010100101011010011000011110;
#1 $display("%b", po);
# 1  pi=207'b011011001001011000000101110010100001011101100001101100100011001101001001101110010001101100110010011100010101101011001000100001111100000100010110000100010111011011000001100010111011010110100001110101011001111;
#1 $display("%b", po);
# 1  pi=207'b000111001011101110111110100110110100001110110001001111100101110010111000010110111111010010101100010001000010011011011000110000000001011111110000000000011101111100110010011010101001100101010111001111101001010;
#1 $display("%b", po);
# 1  pi=207'b010110010110010101001000110011001101011110110000110110011110101101001001000101111101101001111101111110001000111111011000001101101010010010000100111001110111001010010000000110001111100100001101101100011110110;
#1 $display("%b", po);
# 1  pi=207'b000100010001000001011110001101110111010111111111111100000110001101110011000000110110110000010101111000110000011011001001101101100100111110110000110001001011110101010100001000101101000110110000011000001101010;
#1 $display("%b", po);
# 1  pi=207'b100101110110100010101110110111010000110010000110100111101101111111101000101000101110100001110100100101100100010001000010101001100111100111100111011110010110110110101010110110111011111011011111000110111101000;
#1 $display("%b", po);
# 1  pi=207'b011100010110011010110001011101000100101101011011101110001001000011100001110001111000010111000111000111000111011111111111000110011111011100010000001110110010110010101001011001100011101011111001101110111000101;
#1 $display("%b", po);
# 1  pi=207'b111110001111000011011110111011100101110111110110000101111011100001001101100100101011111111001011010011100011011101001011011110010000111000110001011101011000011110010011011001001001011111001010111001000100101;
#1 $display("%b", po);
# 1  pi=207'b001110010110101101000011110111100000100000010100001101110010101110100010100101000010111100101001010011100001000100100100100111011000001101001110001111001001001011110001000101001100110000110000100001001010110;
#1 $display("%b", po);
# 1  pi=207'b000111010110000111100001111100010001000001100011100000011110011011111001111000110011100000000001001011100011001111101100100011101111001111001100010111111100011101111001000011000001001101111110000000100101001;
#1 $display("%b", po);
# 1  pi=207'b101100000101110000110100111110010000000011011101011101100001111110110110011011111111010101100100101010001101000001000011111110010111101000001000010001100100101000010101110111001110101011110111001001100011111;
#1 $display("%b", po);
# 1  pi=207'b010010101011110010000110111110110010000001111101001000001010111100110001001100011001111011110001100001001010000001001110011110110100110110000000101000111110011110010110011100010100001100011000111011110001011;
#1 $display("%b", po);
# 1  pi=207'b011001010100000001101110010111101111000011001011110011101110011100101110100111000110111000011101100110111011110110010011100000101101110100000011111111011101001100110011101000100000111010111000111010000001100;
#1 $display("%b", po);
# 1  pi=207'b101000100000111100000110100001110111100011100111100010100110101001000011010111011001101111101010011010000111100100000111011101000000100110110111101110101000110010111100010010011010010100010010110101100000111;
#1 $display("%b", po);
# 1  pi=207'b011011001110100111100101001110110100010110001001110111010010010110100000010111001101110001010010011101101010101011001100101101011110101000100001011000010100000101000101000011011101011011010100000011110110110;
#1 $display("%b", po);
# 1  pi=207'b000001100100011110100011111101111011000110101001100111000011001000101101010010110011101100010000100010101001000100110111001101011000010011000100111011011010111010101111001111000101010001010100111100001111001;
#1 $display("%b", po);
# 1  pi=207'b101100100101101111111011010101001100101001000101110010111110111111110001111100001010111111001010011010111010111001000010101010101100011101101100100011111111110100100110000111101101101000111001111100010010010;
#1 $display("%b", po);
# 1  pi=207'b100011100011010111110111010101010101101000010100010110011010110110111010100110101001001101100011100010101111001111010100001101101101011011011011010000000010100111111010111101001111110000101110011111111111001;
#1 $display("%b", po);
# 1  pi=207'b001011001111001010011111000011101011010100111010001101001110100110100001011000101101000110000011000101100010001110100100011010000101000100100101010010001001100111100100010101001110110000000101001001110000101;
#1 $display("%b", po);
# 1  pi=207'b011010101010111100100001000010110110100010011001101010111111011000011010000100110001001011111000100110110101000010011001100110101001111000101001001110010100111110111111100100010011111001010000000011111111110;
#1 $display("%b", po);
# 1  pi=207'b111111101111000111010101000100001101011100010010101011100000000011101001001111001100100011111011001011000011011001000111001011011001011001101111111101011010010000010111010110000101100111111110011011001001000;
#1 $display("%b", po);
# 1  pi=207'b110011100111001100000100110010001011111110111110110101000011101001001110001101110011000010001000101010100001110111011000111000101001110000111001110100011010000110110110011010100101001101110010010100000101100;
#1 $display("%b", po);
# 1  pi=207'b001010000011110111110110011100111001101110011101001000101000110101100100100110101101110011111010111111001011011011100011111100010101110100111101011010001110100100001110111010000001101101110110001111100110011;
#1 $display("%b", po);
# 1  pi=207'b110100000010001110000001110011001101100101010001100110000101000010101101100100010000101111000100101110100100100100000011000000101011001111111001110011010110100111000010010010011000100010101000110101001100111;
#1 $display("%b", po);
# 1  pi=207'b001001111110111001000101110000101110010101110110001000110011010010010101100100001000100010110010010010111010001110111111111000100000111010110010110101000100100100100111111010101111101100101110001000100010100;
#1 $display("%b", po);
# 1  pi=207'b001100110111111100101010001001001111011111011110010101110111100101001001011000000001000100100111001101000101011110100110011100111111011010100111010100011001011000111010110111010000101000011110110101011001000;
#1 $display("%b", po);
# 1  pi=207'b010000100101101010101000100111111110111111010001010100011111000100000010010101011101101011011001100100111111101000011110010100001011101000100010010101011010011100000101111110001111001011110011100111000100001;
#1 $display("%b", po);
# 1  pi=207'b001111100100110000110001001110001000101010110101000011000010101011100111110000001101111100011001100000001110001011101001010001010010100100001101110110101011000110101011110110010100110101100000111011111111001;
#1 $display("%b", po);
# 1  pi=207'b111100000011011101011010000000000110010100010010011101101100101001010001000111111000101010000100100111101011011111010111001011101110001010111101110110110010000010101010010001100110110110011111011011010010101;
#1 $display("%b", po);
# 1  pi=207'b011011101110001110111011000010011010110001110111110101001010101011001110101000001111101000000010111000000110110000100010100011011010010010001001110110100111000101100110010010010100000110100100110000110100011;
#1 $display("%b", po);
# 1  pi=207'b101001110110110000101010011100011111001010001100001100110110100001100111101110001010001011100001111110000011101110001110110001000100001010010010010010010010011011001101110001111111111011000101000110100101100;
#1 $display("%b", po);
# 1  pi=207'b111000101110000110110000111100111001001101110100001000100110011101011001101000100100101110111001010000110111011111001001010000001111111000101000010111001010001111111000100100001000111111001011000111011000111;
#1 $display("%b", po);
# 1  pi=207'b011100110010010101100011101011001001100111000011110100110000010011110001011100110101010001000111101001101100010010001011010110110010010110001000011101001110111011011011001101001001010001010000111100000001101;
#1 $display("%b", po);
# 1  pi=207'b110001011100111010011101000010011011111100000100011000001101111010110000100101111100111101111100110001000100011110010011100011011110010110111011111110110011111110010001010000111001101010110111010111011011110;
#1 $display("%b", po);
# 1  pi=207'b010101001000000001010100101100010000110001110001000001110100110000110011110000000111101111000001100001111101011101101000010101101000010000001001001011011000001011100000001010100100000000111111011100001000001;
#1 $display("%b", po);
# 1  pi=207'b000110110011110010101000000100111101011011000101100111000100111110011000110001111011001000100001010100011000100011100010001001110001101011010011111100000011100000011111011001011111000101100110111010011011011;
#1 $display("%b", po);
# 1  pi=207'b010110010001101101100001100101000101111010000110110010001001010000011110110000110011101111101110100110100101010101001010111110000100110111010110010101010000110100110101000111101000101010111000101010000000011;
#1 $display("%b", po);
# 1  pi=207'b000010001101101001010101100000101100100110000010110001001110100110011100001000011001111100110111111100111011100000011010111111001011111111110011001110100101011001001010001011100110111011000011110000111111110;
#1 $display("%b", po);
# 1  pi=207'b000111101110000110010001100110100101000101110100110111110110011110101111001100100010001111000110010010110111010000101111111011000101110010101011111101100110110101011111100110010101110001001000001011000010000;
#1 $display("%b", po);
# 1  pi=207'b111101100111111001011001111101110101010010100111001001011101111111111010001101000100011010000011110101000111101100110100001001111011100011110000100011001000111110100100011001111001110111101000100001100000101;
#1 $display("%b", po);
# 1  pi=207'b110101010011010101111111111011011100000010101001111000101000000101010101000001011011000001110001101110000010101100100001110110100010110010010100110000111001110011101011011111110100110001001001100110100011001;
#1 $display("%b", po);
# 1  pi=207'b101100001111110010010100101001111110001001101000111010100010101111100001001101101111000001010001101100011101101011101001011001100110011101010000001100111001110110101010000110011111010011111011110010000010001;
#1 $display("%b", po);
# 1  pi=207'b111000100011011111110100011100010100110111101000010001000111000000010000010110111101001100011101010010001001110100011010111011001110000010101110010111101101001000100011110110000110010001001110101010010011101;
#1 $display("%b", po);
# 1  pi=207'b010100100100001111100010010010000110101100011100011111011111001111100110110100001001011100000010101010110011010011111101111010001000010011111111001110100010111001011001000110110100010110011110001000010011111;
#1 $display("%b", po);
# 1  pi=207'b000010011001011110000010100110100011010010111001100010110111110010000010000110110011111001100100101011100000111100111101101001011101011011010110101111111000000100100110000110100011111101010001111001000101011;
#1 $display("%b", po);
# 1  pi=207'b000001100000011100011011011110101010001101010110100111001010111010111101110011000001111011001101100101111010011011001110110000010010000101000101001000101001000011000110010110000101100000010010100010010110100;
#1 $display("%b", po);
# 1  pi=207'b001011111100011000000101011110001101101110100010001111000100000000110001110011111001100110100010011010111010011111001011011110101010100010001010111101101110000111001101100011001110100101011101100101000110001;
#1 $display("%b", po);
# 1  pi=207'b001011001100100111001100100010101110101010100101110101001101011001111011111100100001010000100000111100010011100111101100001011101100110100011100010101011101110110000001111001111000001100001010111111100011101;
#1 $display("%b", po);
# 1  pi=207'b011110110111110000000010101100111001011110001100111000001111000011001110001100010111001110000110011010011001101111011100000001000011001110011010010011111101000001101110001001011100010011100111001001000011101;
#1 $display("%b", po);
# 1  pi=207'b011001101010101111110011001101111000100111000100000001011100100100011101000111101011100010010110101100010010010110001101010000000011011101100001011110011100000110111000101110110001010001110011000111001000011;
#1 $display("%b", po);
# 1  pi=207'b000101110100110010011111111010001000101111001111111110100000010010100011101000000111100001011101000100011101110101001111101111011011110110111111010011101100001101111111001011011101111101001000111011100110101;
#1 $display("%b", po);
# 1  pi=207'b001110100011101100001011100000000101001110111101011000011111111011000101101011001000010111011001011110111001000000000111011111111001101111001000111000011101100110110111111101010101100011110110101000111000000;
#1 $display("%b", po);
# 1  pi=207'b010101101100011001101111111101010101000100101110110111111111001100110110101111011011010011011001011000101000111110101110110001110011111111110000100110101010101000110100010110101100110110011011010100010100000;
#1 $display("%b", po);
# 1  pi=207'b110001001111011100110001100111000000111011110010100101110001111100010010100010000101110100011111110110100110011001101010001000000001001101001001010100010101100000100101110010011010011011111000110101101111101;
#1 $display("%b", po);
# 1  pi=207'b011111111000011010001000100001010100111101011100000100001010010101101000010001110000001000110100001010001011010011101010010010110110010010101100111111101000111011110000110110101101011111000100001010111100111;
#1 $display("%b", po);
# 1  pi=207'b010001100010111100011001111111011010100100000100100111001111001011111001010011110011101100101110010010101110010011110011111100100010111101011001110111100101110110001100111010000101111010110111111001110111010;
#1 $display("%b", po);
# 1  pi=207'b101001111010010011100101010010000101111010001100001110111101110100011110101011011111001001000011101001101000011111101101001111011001110111010010011101001010010000010011011101011010000100100011000011111101100;
#1 $display("%b", po);
# 1  pi=207'b111111111111001110001111011010111001010100110101111111101101001100111001011110010011001011000001000110101110011000101100011001000001001101100001010101000110010000001100001010101111010110111010101011111010101;
#1 $display("%b", po);
# 1  pi=207'b011001111101000100010110100000000100110011010101011010010101010100010000111111101110000111000100110011101010100100111010110010010100110000000011110100111110011011101010110100010110111010110001111001110010110;
#1 $display("%b", po);
# 1  pi=207'b101110001111100010010010011101101111000010110001000110111111111111101100000000010011110101111101000000101000010101011001010100100110010010000110110011110110000101001000111011010100011100001100101011000011110;
#1 $display("%b", po);
# 1  pi=207'b110110100000010001000110000011101001010011101010101010000100110101110100100100011110011000000001100000001101110100000010100111110100001010011100111111010010001101000111000111000100010001001101000011100001000;
#1 $display("%b", po);
# 1  pi=207'b001001001010110100111101011101000111011101001110011100111010110011101010001101010011101100100111010111011000100100111000011000111101011001110100110000101111101101111110001010111000101111100111011010110101010;
#1 $display("%b", po);
# 1  pi=207'b001000010101000101001100011110101110011110000001010001011100001010100011011100101001010011011010010000111111011111001111011100001101000100110011010111111101000010001101111110010011000100011100001100100010010;
#1 $display("%b", po);
# 1  pi=207'b001101110010000111111001000101100010111001001011010001110100001111100111101001011101100100100001111011101011010101010100110000000001111001010011010000000111110100110111011111110101000010010001101010000101110;
#1 $display("%b", po);
# 1  pi=207'b010100000010000010110110010100001101111011100111101110100110101111100010001010100111110011101000001101111000110000010101001101111011010111100111011001101111010001001110010100101000010000010001000100110000111;
#1 $display("%b", po);
# 1  pi=207'b000101101101011010010000000010111001011100101100011110000011101110101010000111101110100110100101010101100011001000111001110101100101000100100111100110010110111001100101001001110101010111110111111101011100011;
#1 $display("%b", po);
# 1  pi=207'b011001100110100001111100011000110110001011101001111111011001110010001001101010011100000100101111010000000101000100100000000110011110111000001111110101101011011111100101010010000010000010111101110100000100110;
#1 $display("%b", po);
# 1  pi=207'b010111100001101100100111001001111110010001110100111010001100011110000000110100110110110110110101100111101000111100001101011111100011000101000001100111100001111111101110100100011100111000100110110100011001110;
#1 $display("%b", po);
# 1  pi=207'b110011011001111001001000101001111111110011101100001000000110110011001000101101110011010001010011011000011100111001001100010110100100000100000000000100010101010111010110010100100110111111001100010100110001100;
#1 $display("%b", po);
# 1  pi=207'b010110100000001011101010011101011101101000011101100010000000011100000110011101001010101011001000111101100001111100010101011000111110111100001000100001100000110110001010100101011001111101011001010000111100011;
#1 $display("%b", po);
# 1  pi=207'b011000001110111110101011000001001011001101110000001101100001010110100110010001000000110111100000000100101001111001111001111011101110110011100110110110100101010000011111011101111001110100111100000101100101000;
#1 $display("%b", po);
# 1  pi=207'b010111100001100011100100101101001010100000100110001111000101010011101100000101111110110001111110101110110111011011011010101010101111011010111001011100000000100101010011101001110000000100100101110111000000010;
#1 $display("%b", po);
# 1  pi=207'b101010001000110011011101011010011010010001000011011010010110011100100100000011011111100000011001110101001100001110101010011000001000101000101101010011001000010000110100100111111100001111111011100110101110010;
#1 $display("%b", po);
# 1  pi=207'b011110011110111110011111111010011011010111100101001010110110010111001100111110011010100000011010001101110000111001100011010111011111010111110111001100101100101111101011001000100010001000001000000001010000001;
#1 $display("%b", po);
# 1  pi=207'b111000011000001001110011010100001101010110000101010111011100110101000100110110111000000000110011111001100000100010110001011101011010111101100010111111101010001010111110000000101100110001011000110001111100111;
#1 $display("%b", po);
# 1  pi=207'b100001011110010001111001010011111000111000001110001100110010111010011100101001000100001110100111001100010100110010010100110010011001010001010000000001101011001000111011111101000100010011011101100100111101110;
#1 $display("%b", po);
# 1  pi=207'b111000000111101000101011010011100101110001001110010110010110000001100011101100000111111000000000011010100001000000010110010101001000000001111010100010101001111011111101001000010001100101011000100111000100010;
#1 $display("%b", po);
# 1  pi=207'b011000001001000001000111001100101111110111110011001101110011101100111101100010001000100010101011111010101100011010001110001101001110100001100000101011111101100110001111111000100000110011010111110110110010111;
#1 $display("%b", po);
# 1  pi=207'b110000100000001000000001100110011101111001110000101001111000001110110111111000100011101111111001011000000110100010000010001011011010010010110100001111100111011011010011101011000111101110001000100101111110010;
#1 $display("%b", po);
# 1  pi=207'b001111010110111010110100110010000101111011100010110001101110001100100100111010010110111101010110001001110100101000000000011101101101010000111101111111001101100110110010100100011100001001100100010101101101000;
#1 $display("%b", po);
# 1  pi=207'b111001001000100011100011000011000000000111011110100001110110010000000000111101111111111011100000000110110001110001110110110100111101101001100010101000111000010110000111110011111011011100000110001111000000100;
#1 $display("%b", po);
# 1  pi=207'b101011110111010110000101001000100110110000011111111110101000000100100000000001110011101010011011011001011000000110100110110110011110110001010010001111000111010001100000000101010111110101010010010001000100100;
#1 $display("%b", po);
# 1  pi=207'b100110100100111110111101101100001011101110011011010001101110000000111011011010111000010010011101110001001101000010111001111111010011011001101101010000100000100101100010111111100111111001001001110101101101011;
#1 $display("%b", po);
# 1  pi=207'b001011110100110110100001001010111001000001000010000001000000000011011101110010101100111000101100011000100011110111110111001011101011000101011011110011101010000111100101111111010010011111011000100000111101101;
#1 $display("%b", po);
# 1  pi=207'b101001000011000110001001001011100111111110111111011110111000111100001111010100010101110011110000101010110100001010110010111101011100101000010010110101011110101100100111000101110010100111000011000110000101110;
#1 $display("%b", po);
# 1  pi=207'b100000011011111101110000100000001100101100111100110101011100110110010000101011110111011100010110001001000001110011111111011011111110111011000100100100110001110111110110010000110101011101100100111011010011101;
#1 $display("%b", po);
# 1  pi=207'b010101101001001101101101110110100000000011110111001100001111100000001000111101101000110000101100100011011100001111111001011111010101010101110000111000001010011001011001111001011001000110010101100110111101111;
#1 $display("%b", po);
# 1  pi=207'b100101111101011000110111011111011101101001011011001001010010001111101111010010000010001000110000001111101001110101101101010110000001010110011100101110111101110110110110010100101110000011101111110110000011100;
#1 $display("%b", po);
# 1  pi=207'b010011101100010110110010100001110010111101110000100000111010111000111110110011101101101100000111101110111111100100110001100001000111101111100101100001010010110011111100001001100111010011110010011011010101111;
#1 $display("%b", po);
# 1  pi=207'b011110110010001111110011111001010101111110011111001110111001001010100001010101110100010010001101101100001100101101100001101011101010010111110000111111100110101000011101010100001010111001101001101001111011110;
#1 $display("%b", po);
# 1  pi=207'b101101100111001001010001010001100010001111111000001110010100010001010000000001011000010000110110011000001100000001000000111011100010001111111110101101001101010001001001000001011111001111111001010101111010001;
#1 $display("%b", po);
# 1  pi=207'b111110111101010100000111011100101111111100101001001010111010001111011000101110101000010011101001000000100111111110001011000001001000101111011011110111010110010110110100000101001101111001001111100101010001001;
#1 $display("%b", po);
# 1  pi=207'b010001111100010110101001100001101110110100100110001010010011011000000110011000010010010110111111001001001110110011011000101111111000001010000101011001100011000000110000110100010101000101110101111000010010110;
#1 $display("%b", po);
# 1  pi=207'b110010011001101100001100010001111001101001111011000001010111011100000011010100100101011111001110101100011100001000010000111010010010110011011001010001000110111100110110110000101100101010110000100111010010111;
#1 $display("%b", po);
# 1  pi=207'b010001100001101000000011011101001010100010001101001111001010101111100110000001111011011011000101010011111010000111100111010101100100001110110010001101111101001100001111101011101011101000111110100110100111100;
#1 $display("%b", po);
# 1  pi=207'b000110001000101011111110100100110110010111101000100001000011101100101000111100101000100000000100110100011100111101010100100001011001001001100111111011001010110100100001111000011101001011010110111010110001001;
#1 $display("%b", po);
# 1  pi=207'b010000011101100010010100101000011110101100111111110010100111101100101111001100111110110010100000110011110001000000001110100110101110111001010100010101011010100111101000011110001000000000011100100000011101101;
#1 $display("%b", po);
# 1  pi=207'b010101001011110111000110000010000110011010000011010011111110100000101111011010011110010001110111101010000000111001011000100100000101011011101000010100001110111001101111111011011011001110100111111100101010010;
#1 $display("%b", po);
# 1  pi=207'b111001111010001100110111011011000000011111000001000101001100100011000100000010011011110110111001101100001110100001011111111011000011100011010001001111011100000100101010101100000000000101010110011001111110011;
#1 $display("%b", po);
# 1  pi=207'b000000111110111100011001000101011100100110101011010000010100000000011000010101100111011101110110010101110001000010010100001000001001101111111100001100100011001010101001101001010011101101111001100001101001101;
#1 $display("%b", po);
# 1  pi=207'b101110110011001000100001011001010001011111010010000000110110001110111011001001000101111100001101001101111100010100111011011100110001100101010100111101011011000110110011110001000011000010101011110011110111011;
#1 $display("%b", po);
# 1  pi=207'b110110000110000100100000100011100111100001110100001011100110100101111001101110001111100000001011100001010001011001001010000101100000100001101111110001010100010011000100011001000110111111111100110100101101111;
#1 $display("%b", po);
# 1  pi=207'b101100111001011010011000111010100100011000111100010111010101001010001101110010100011011100010101111011100000101011011010110100000011011001010001001111111111010001100111000101101010011111101111110101000111101;
#1 $display("%b", po);
# 1  pi=207'b001001111111100011111100100001010111100010101001001111001111001111010101010100000011000001001010110100001001000000000101110111100011010001011100100111000011100000100001100111110110100111000000111011100100010;
#1 $display("%b", po);
# 1  pi=207'b010111100010110000000100001010111000011010011101111100100000011010100101010101010101100011001001110101000010000110010011101100101100010110000010111110100101101001101001100001000000001010000101011101111010001;
#1 $display("%b", po);
# 1  pi=207'b100001011011000011000001110001001011101111100000011101110110100011100101111100000000111001010010010111010111011100110010010111010001100001011101000111011001111111101101000010000001100011101110001110110011111;
#1 $display("%b", po);
# 1  pi=207'b011010111101110111111000110111000011111110110011101000000001101111100000111110001011001011110110101111110011011111000111110001110101111101011001100011111100001110000010000010001111010110010001001000111001001;
#1 $display("%b", po);
# 1  pi=207'b000011011000011001101100000001110011100110001000101000001101011100001101001000110110101010000000001101101110100011011000000100000010101010111100001101000011110111000111100011111111110000011101101101100000010;
#1 $display("%b", po);
# 1  pi=207'b100010011111011000000000011000100101110100110011100000001011001110001011111001000110111010111101100101010010011011100010000011111000000011110010100000000101010010110010000100010101001100111000000001100011010;
#1 $display("%b", po);
# 1  pi=207'b001101110110011100111111011001100000100100111001111000101011001011110110110110110010000100000011111001101101000100110101110111000000110010101100100010001100110110011010010001001001000010101110111011001010111;
#1 $display("%b", po);
# 1  pi=207'b001101000011110010011010000101011000011011100011100111001000000001111100100111100111110010110100101110000100001110011010101100110001111100110100010011010111001000000110110011011100100010000101110000100010101;
#1 $display("%b", po);
# 1  pi=207'b001101000101000001010110100000110100101101000011111100110010110011011001000100001011011011111001111100110110001001011111100101101010000011001011111101011011111001010101101001100111000101100100001101010001110;
#1 $display("%b", po);
# 1  pi=207'b100101110100111110001100110101011010001110001011110100000111011000101111001111001011000110010111010001101000100100111011110110010010100010011000010011111111010100110100000110011011001000010010011101000000110;
#1 $display("%b", po);
# 1  pi=207'b011100001100110110001110000011000010100000011001000111101110001100000111011011101111001010101001110000110100000010101100011001111010011001000000000000001101111000010110110101101001100000100010011111011101010;
#1 $display("%b", po);
# 1  pi=207'b101110100010011011101110110001100001010010011001101011110010010000101000110000001110010100110110111100110010011110010001001101110001100010000000011000101010100011001010001000010011000110000001001001100111101;
#1 $display("%b", po);
# 1  pi=207'b011010011111110110001010010101101111000010010110100111010111111011110100100001101001000001101000111101111110110111010010111000001110110111110100000111111110111010111110000100010100100000001100001001011110001;
#1 $display("%b", po);
# 1  pi=207'b110010110101010001111111001100100000010101110110111011110011001011110110011101101001111100001100100100000000110011011110001111010101011001111011101111011001110010000011010001101000100111010010101110000000000;
#1 $display("%b", po);
# 1  pi=207'b001000101111110100010001110011010110101000010011000110001000010100011011100101100100101110011100010100100110010000011000111001100101010110111101010111111111111000110100010001101011110001010001000001110010100;
#1 $display("%b", po);
# 1  pi=207'b110101010101011011100101111101001010010010011110101010111010010010001000010001010110010110110001011100010000000100001101011011010100110010111000011110100000101000111010110001000110010001110100011010011001011;
#1 $display("%b", po);
# 1  pi=207'b010011100001001111000000011011001110001111001000111100110010111100101110001100011110000110000110111110010010011101011110000100111001100011001110101100010010100101111110000111000001001000000000011000111111011;
#1 $display("%b", po);
# 1  pi=207'b111110010100000010010000001111001001101110000000101010001101000111100100100101101011010011100001010100010110000101001111110101000000110000010001001010000011100011011001100001001100111000110111110100100111010;
#1 $display("%b", po);
# 1  pi=207'b010011000110011011100000011010010101001110011111101101011100011100111111011000001001010010100111101101100101111010100011010101001000110101110010100110100010111101001101111000100100010101101010100011011001100;
#1 $display("%b", po);
# 1  pi=207'b000101100100011110001101011101000110000101011000011100110011001100100011000110001010101010001111000111110100100100000011000111110000100000010110100100010100110000010100001001101010001010100101110010000011010;
#1 $display("%b", po);
# 1  pi=207'b111010010111111111010011111000111000001101111000110101010010011111010100101000010101100010100110101010001101001111100101101000011011111100100001001111011110100011100011011011110010101111100111110011111101110;
#1 $display("%b", po);
# 1  pi=207'b001001001110111110111100101100100010100110011101011111111011010001110100000000001100001111001110011111010100101010111110000111101110110010100010010010000100000110101111011011011011111010111110100111111111110;
#1 $display("%b", po);
# 1  pi=207'b010100111110000011101011010101011100000011010101000000000101000101111111101000000100001110101100101101001101011110011001100111101001110001101101100010010100110101011100110110100011010010001101000000011100111;
#1 $display("%b", po);
# 1  pi=207'b011110101100001000001001111111100010100100110011000011100000110010111101100000001011000110010010010000000010010100011001001100001101100110001111101000011100010100001001100010110110100111110110011001001011101;
#1 $display("%b", po);
# 1  pi=207'b111001100000000111011110001110010011110010111100010011001101001100110110011001101110101011111111110100111111110001011000110011011011110001110001110110001011111011000000001010100111101110001110100000011000011;
#1 $display("%b", po);
# 1  pi=207'b100011101010100000101100001101101011100100110001111111000110110111011110011100001000010011011100100100010101100110011100111011110100010100110101100010000011010100001000101000001100101001001100001000000111111;
#1 $display("%b", po);
# 1  pi=207'b100010100100010101010001011011100101111101000100011011011110010111111011100011111111111110111010100010011000010011101101000101011111001100110110011111111010101100011100011001111111100011110111001001111011101;
#1 $display("%b", po);
# 1  pi=207'b110101011111011001000011010110010000001010100000001100011010001111100110111110101101001001111010000110110111010111001000010100000000000001000110010100011100111011000001111000100100100101101010000010101011100;
#1 $display("%b", po);
# 1  pi=207'b011101010111000101110000000000011100100101001111100001001000111100100110000101001101111100000101001010011010111111000000000001010010100100111011100111100110101000010011000010111000001000001110011100011110100;
#1 $display("%b", po);
# 1  pi=207'b101100000110110011111000110000011111110100110101010100100100011111110000101100100100111101001011010010010111110110100101101100011011111001111000000000010011100100111110110110110001000110101111000100001101101;
#1 $display("%b", po);
# 1  pi=207'b100110000110100101111111110110011000101001110100100100111001001011010110110000100110101110110111011101011000001000011101011100111101101100100000001101011011011110011101010101010011000100000010111011111000010;
#1 $display("%b", po);
# 1  pi=207'b000011111000110000010011001000011001100110100011100000010101110110011011001101111001111000001101010101011000100101111100010010000000110011101000010101100101101111101001110001111110101111100111001101000100110;
#1 $display("%b", po);
# 1  pi=207'b000000110110111011010001110010011000010010100010001011101010001110001111111111110000011010010011000011000001111010011000111110001110111011110000100111011110110101001101111000001100100000011101011001110101111;
#1 $display("%b", po);
# 1  pi=207'b000011111111000111110101110011100011011100010101101101000101010101101001111000100100001100100111111001100000100111110011101000010001000001010010010100110101101011011010101100011011101001001000101010100110111;
#1 $display("%b", po);
# 1  pi=207'b111000011100011001001011001111010110101010111111000011101010110000100100011110001100101010011011001000010000100100001001000010101101101000011000100110110100110100000001010011001010101010011101110001011100011;
#1 $display("%b", po);
# 1  pi=207'b010110000110111101011110111010100111011111110111111001000101110000111001111100001010011000100010100100011001101100100011000001101010010010101001001011001001011010000110011000101011110110111111000011000010101;
#1 $display("%b", po);
# 1  pi=207'b110001100110011011101001001000110101010100001001011101000111100000000101101101000110010100101111101111011001111100001000000100110101101111001110010110000000011001001100011010011101001001101000010011101010000;
#1 $display("%b", po);
# 1  pi=207'b110100101001011000001011100110111101000011011111100000100110010110011000010110000111110100111000101001111100011101100101101110100111100100110011000101000010011001110111110001101010111111101011110110100111010;
#1 $display("%b", po);
# 1  pi=207'b010111010111110110101010111101100011011011111001100011001000110001010000011111101001100111010100001001001111101010110010111010010100000101101011010101100101110011100001001011100111100100000010000110111111111;
#1 $display("%b", po);
# 1  pi=207'b000100101000110001001011101101111101011111001100000101010011101001101101000101010100101111110000101010011110010011111110111000010111111010001110001000110101110111111101010100000110010010111111110101111001100;
#1 $display("%b", po);
# 1  pi=207'b011110010100011111000100110101100110101001000110001101000100010101001111011001010001001000011110010000011011010101011111111010010101111111101000011110111000110101110110110110001111000011100010001001101101000;
#1 $display("%b", po);
# 1  pi=207'b101111010111110100011101000000000001100010110111100010010000001101111101010100110111001101101011010001000011000011010011001110001010101010100000000001010000000010111110010100001000000111111101101111110101011;
#1 $display("%b", po);
# 1  pi=207'b110010000110001101010010110100010011010111010100011010101001111100101001111010101010110111100000101101110010000111101111000010101101010011111110110100100110100110110110111000000111000101000000110111101111010;
#1 $display("%b", po);
# 1  pi=207'b011001001100100111001001010101011010011011101101011010110001011100000111101010001101100110011010110111001000011000011100010000010001101100110010001100101000010101100111100101101011010110100101100010000111110;
#1 $display("%b", po);
# 1  pi=207'b111011100001010010001000111100100000010101111101100111000110000100100010101111100101111101010010011011010101100010000100010101111100011010010011100111110011010010101110111110000110100001010011110111110000001;
#1 $display("%b", po);
# 1  pi=207'b100101100011111101100011110101111001010100101100100110110110001000100001110111111111011010100100011100000110011001010001111000000000010111101100000111100011010001111001100010111101000011101001001101111100111;
#1 $display("%b", po);
# 1  pi=207'b101111111001011100101110010111111110010110001011000100010101001110001110000110101000110010100111111011000111010011000101010101100101111111001001100011010011000001111111110000011011110101001001001110001111010;
#1 $display("%b", po);
# 1  pi=207'b010110101010010000100011001000011011101111011000011001010111111001001000001111001000011100110001011111111010011111010110000011000011000101110111111001001011000011101111111010100100111110001100011110111100100;
#1 $display("%b", po);
# 1  pi=207'b011110000100101110010101011000001111010000001010011011001011010010100000010111101100101000010001100101010011101010100101111010111001111011101011000100000011000100111011100011111001100001010101100010110011100;
#1 $display("%b", po);
# 1  pi=207'b000000110010011011000011011011001101110011001111001000111010011011000111100110000111101110011111011001010011100010000100100010001010001011010010000000001110000100001000111100101111100011101001100100000111011;
#1 $display("%b", po);
# 1  pi=207'b100100101000101010100010110111011010111010010111010000110100001111101011000100100100110101000010111011111010010010011101100100110011111110000010101111000111001101001111000101111010100001100010111110001111001;
#1 $display("%b", po);
# 1  pi=207'b101101111010100111000011101000110101100010110111001011110001110000001000000111000011001010001110110011000010001001011001000101101011101001000101001111110101000000101010101101000101110011011110100101010011101;
#1 $display("%b", po);
# 1  pi=207'b010111011011100011000011110101011001001111101000110011111001111100111010100000100010001100101001001101100111111010110010011100111010110110001011100100010110000100001001111101000000111010011011111101000111010;
#1 $display("%b", po);
# 1  pi=207'b100101110101110011011011101111110100001101111011001011000100010110000011001100000000100101010000100111100010100001011110000011010100110010010000001110111101111111111011100110011110001001111100110001010000110;
#1 $display("%b", po);
# 1  pi=207'b100101101110011101100011110000110001010001111100101000010001101100100101110011110110110101011110000100110100001011101010101010011100110010110100011101111010001000011100000011000100101110011110100011010100111;
#1 $display("%b", po);
# 1  pi=207'b111101001000001101001000010010101100000101010010110010000010100010000100111110101011011101001011100010100000111100011101000101110110110001111101101111011110101010000111101010011000110010110010100100111010011;
#1 $display("%b", po);
# 1  pi=207'b110010000000011110010100100101100110110011111001010010110110111001010110001111011001011110101111011000101001011010010111101011000000111111110001010111010001001111111001111001000011011011111001000110000001011;
#1 $display("%b", po);
# 1  pi=207'b100010011011000111111010111100100001110011011000110011100000011111110001001101101111001011111101110010100010000111001011101000011100011111010010111000001010011101010001010001010111011001000001010111000101111;
#1 $display("%b", po);
# 1  pi=207'b011010111000110111101011011100100111101001001010111011010110001101000100101101010100011011111001010011001010011100111111100110111000001011101100111110000010000010011010101111001000010000111101000010111100010;
#1 $display("%b", po);
# 1  pi=207'b110011001011001101111000111111000001000100011000001111011000010001000000000011110011100111011000001001000111100000100111011010001011111100101000100111100101100011100001100111100100001101011100110010000011010;
#1 $display("%b", po);
# 1  pi=207'b011100000111110111110010011111001100001111101110101110111000001000111010000011111100110011100100000111111011111010100100110100110000001011010000011010111011111010001011000101111001100111001011001000111010011;
#1 $display("%b", po);
# 1  pi=207'b000000101001110000100110010011101000011001000100101110000111011110100001011010001001100110001001110010111111101010001110011010011111000111100111010001110010100010001110001011100001010010111110000000011100110;
#1 $display("%b", po);
# 1  pi=207'b101010011000010100110101110000011000000110010000101001110000011000101010001101101111110100111000100001101000011001000010011100010100010011101101000100001101001010001100101001001010110111111110101110110001011;
#1 $display("%b", po);
# 1  pi=207'b001010010011000110001010110100100111111111010111110100110010010100100110111010001101010100110110111110011001101101011111101011001111101100011011101011011010000100000111111111111100001010110010101101010100111;
#1 $display("%b", po);
# 1  pi=207'b101101100111110111110010101101001000000100101110010010001111101010100110111101010100110111111001110110010000100110111111001100000000010100011011001000010001001010001100011111001101111111101011001110001100111;
#1 $display("%b", po);
# 1  pi=207'b100111110101110111000111001001111011100011010010001101011000111110001010100111110001001101011000101011011101111000110001110000010001111001101000111100101011110011001010001011010111100011000111010100111101010;
#1 $display("%b", po);
# 1  pi=207'b010110111001000001110011100000001111011010001100011100011011111100011000011101111101000101011100001101001101000101011100011111010000001001101111100010111011000011010111011000011111010001011110000100001000110;
#1 $display("%b", po);
# 1  pi=207'b101110001101001101100100000111001100000110000001010011000111101011101111101000101111111100111101010000111001100111000100000101001011110000011101100101101100110010100000101110100110000011110011001110111001110;
#1 $display("%b", po);
# 1  pi=207'b010010100011100011111001010001010010111111110000100100010101000101010011010110001000100101101000001100010111101100011101011111111111111100100100001011011101011110110110110101000011000000110001111100110101100;
#1 $display("%b", po);
# 1  pi=207'b010010001001111001101111100110011000110001100000000011101101101100100011101011001100011110110100000101010001100100011110101001001000110110000000101011001110011010101100001111110101110011001001000001011011100;
#1 $display("%b", po);
# 1  pi=207'b011010000110011001100001100000010010101111001110100111000101001010000101101110001011111001001001111000010100000011010100110111000111001000100010001111111010011001010110000001101011000101010100111101110100000;
#1 $display("%b", po);
# 1  pi=207'b100001001111100001001110011001110000010000111011000110111001100101101001100110000110011100100100001000011000100001001111110011111011100011011001101110010011001001011011010011111010100001110110010010101010100;
#1 $display("%b", po);
# 1  pi=207'b010011001001001101011011001001101101100101100011001110100100001010001110101010100111101011100100001000010010101010100000110000100101001101110101101001001100111101110000111110101001110111010110100101010000101;
#1 $display("%b", po);
# 1  pi=207'b100110101011001000011001001000000000010110010010000000011001000110110100001111111110010101101101101000011011111001111011111100010111011000011011110010011010010110110011101110010011001011110011100110110000011;
#1 $display("%b", po);
# 1  pi=207'b001010000001111110011000000011101000110000011000110101111011100010101111000001110011000010111110111000111101101000011000000010110001110111000111001100111100101101111001000100011110100011000110101110000010011;
#1 $display("%b", po);
# 1  pi=207'b000001000101010100001110100100111110000000011011010001001111001100110001111110011000101100001010100011000000010010010010111011100011111101101000100111110110111010110000100110000100101101000001000011110111101;
#1 $display("%b", po);
# 1  pi=207'b011010000010011110001111110101101101101110011110010011110110010011011101000110000000101111010011010010101011001001001011110101100000001010100001011011010111000111100010000000010000001110111101000101110010000;
#1 $display("%b", po);
# 1  pi=207'b011011110100010011010000111000000111110010100011111011100110110111000011011110011001011010011001101101111011001101111101000011010010010100111000100000110001011010011111011101000110101110111001100001111011000;
#1 $display("%b", po);
# 1  pi=207'b110000100001111001110100010001110000111001110100101011000100001001001101100000000110101001111101100101010100001000100001100101111110010010101110000011111111111011110000011011100101110110001110110110000011000;
#1 $display("%b", po);
# 1  pi=207'b101001011101001110000001000110010010100101111111111010111111000101100010100001000100100010010110111001000011111101100010101101110010110010000011010110000110010010001011101111001010011100100011001101011110000;
#1 $display("%b", po);
# 1  pi=207'b000100111110100001010011100111001101101100111001101111010100011101101000100110000001010100100110110010000010101111001010101010011001001011001000100111001111110011000110111100111001001000101110101011000111011;
#1 $display("%b", po);
# 1  pi=207'b010000101111100001110000110111000101000010000110110010110100111000111100101100011001010101111111001010010011101010000000110110010110111110010100010100010111010101000111110101011000101111101001100000101110010;
#1 $display("%b", po);
# 1  pi=207'b001010110000101111011011100001101101001100010111111011110001011101100110011100101010011000101111111110011011111000010011110011000010111010001000010011111000111111101110011100001110101110001011001100010100111;
#1 $display("%b", po);
# 1  pi=207'b010001010010100101101100010110101110011001010100110111010011100111100000101101001100010110010110110011000001010101111001100111011100101011110011101001000011010111011111001011010011101101001010110010000000111;
#1 $display("%b", po);
# 1  pi=207'b110111111000111010101000101100011011001100100111111000001100111000111100011011111011001110000000000101011001111111001011011000000011111111110000110001100000011110001011010011011001011010000110101001111111111;
#1 $display("%b", po);
# 1  pi=207'b000011000001001011000111011101111011110000000000001101001000001010100011010110111111011100011100000101000010000100110111111101000100010100001000010101110000010010011111001111011100111011011011111001101101100;
#1 $display("%b", po);
# 1  pi=207'b110000001010000111001011011110101101110100001000011011101111101001111110101000001010111100001000101111011111101101010000111111110000110010001100100111100010101001111111011001110010100000100100000110101100111;
#1 $display("%b", po);
# 1  pi=207'b010001101001010010000100011110110010010011011011101010000001000000010000101111101000010000001101111010111011111110101011011111111010100010001001010110011101111110011111010011110101001110100111111010100011000;
#1 $display("%b", po);
# 1  pi=207'b010011010011110010001000011100001010010111110000110100000101110011011111010010001000011001100110101111100000011111010111011111001110111110100011000111011110110100010001110101111111100101011011111101100100001;
#1 $display("%b", po);
# 1  pi=207'b101110001111110001011100101110110100100010100010000100001011101011110110101110100001010111100100001101011110101010100010000000100010101111111110000101010100011011000101111010111000000010011110110101111101001;
#1 $display("%b", po);
# 1  pi=207'b010100000000011000010010010001001100110100110101111101001001100011111101100010011000001001000011010100010110000100101000010110010110001010010111010011111111111001001100100011010000111110111010000101101001011;
#1 $display("%b", po);
# 1  pi=207'b001110100111100010100110110010100101001010110010101110010100011010011010010000001000100011010010000101010101011011010011100010101111111001011001110101111001110110100110010001011110000001001110101010001110000;
#1 $display("%b", po);
# 1  pi=207'b101111010000101110000011101111010111111110011101101011111101110011000111010110111010010110011110010111011011101100011111100111100010110011110000001110010000111001101000001001000100110000100111010010001101010;
#1 $display("%b", po);
# 1  pi=207'b100101010111101010100000010010011111111101110100010100010011100000001111110010110110100011111000000010000110111000000101111001001001110101100111111001000010110011010011110100110110000100100010011010101011010;
#1 $display("%b", po);
# 1  pi=207'b111011100110001000010100100000010110110110111111100111010110011001111100101110011011110101100110000000110001100100011011001000011100001111101100001001110100111100111110010010110110101101101010100000101110011;
#1 $display("%b", po);
# 1  pi=207'b011110100100101101011110010110100011110001001111101010101011111101011101110001100111101000101011001001111001100010111011100010000011101010000000011011010110111111011110011110111010100110110001011000100000001;
#1 $display("%b", po);
# 1  pi=207'b101011010110001010001010000101110101111010011000101010000111001100100100111000110000110111100011000001000110000010001111100001101110010001001110101110011000100100101111110001100100101001000000100001000110110;
#1 $display("%b", po);
# 1  pi=207'b010001100000001011000110000000101000100001100101101110010110100111111011111100001100110101000101111010111100010110010111001111100000011011110001000011100001011001010100101010011100111101010000100001000011000;
#1 $display("%b", po);
# 1  pi=207'b111111101101000100010111110100101110110111101100010110011110110111101001010001101101011110110110101110100100010111010110001010011110010000110100000111110001110101000110000001100011101101111010011101100011101;
#1 $display("%b", po);
# 1  pi=207'b001100101111110011100110010001001111100011111101000101010110111110100111001111110010110001010010001000110011110001001110011000100111010000100011110000100001110001111101101010011100000000000000101100001000101;
#1 $display("%b", po);
# 1  pi=207'b110100011100000110001111001101101111110101001101101000011101010110110000100100010011110101010100101110111111011010001000111110100001101010010100011000000101110011011100101101000011111111011000010011000110111;
#1 $display("%b", po);
# 1  pi=207'b011000010001100100000000001010101110110011110111001001100100001111110111011000000001101111001100001011001100111111000100110011101000101011001001100111110101100010000001110101001000110011000111001100000011011;
#1 $display("%b", po);
# 1  pi=207'b100000111001110000011010101001110010101100110101101010100011000011010111111010001010100111010001110000110101110100000100011010100111100110100001100101110011001011101011011111001001111101111110101101101101110;
#1 $display("%b", po);
# 1  pi=207'b001110001100001100110100001010001111001110101001001101101101101100000101010011100110100111000011100110011101000111010010111010000110100011011000000110110100010000110111110001111000101011000001101101110010001;
#1 $display("%b", po);
# 1  pi=207'b111100100001000111001110100000101001010110000001100000111110010100110101010101111111100010001000100001000001100101101010000000010100110101010111001001101110101111101111101011001100001100011111100001010000001;
#1 $display("%b", po);
# 1  pi=207'b000011100110101100111100110011000011110111000110010111110110100001110110010010100011100101110101111110011110101110001111101100000111111011001111011100111110111100010111100100100011100010111100100000100000001;
#1 $display("%b", po);
# 1  pi=207'b100100101100111010011011010000010000100001001010111001100100011001100011001101011000111111110011100011101110001111110001101111000001010100101000011110000000110010101010111101000001111100100010011111000110000;
#1 $display("%b", po);
# 1  pi=207'b101101011100011010110110010111101100011100110011010001011001001010001000010011101110101101110101010110000101100101100110000100000001010000011100100101011000000111011111111101101000011000011011001100101111010;
#1 $display("%b", po);
# 1  pi=207'b000010101101011101011011001011110011111000011011000010011101001000000011011111110000011100100011001110101010101100111010100101001111110000111001001101010110110010101111000011100111011010101000001001000101110;
#1 $display("%b", po);
# 1  pi=207'b100000001100011100011001001000000100100100110001111111110000010010011101111111100000011110010100001011010101101100111010000011010110011101110000000001010100100010000010111000101110100011000001101011111111010;
#1 $display("%b", po);
# 1  pi=207'b010010111010011100101010001011001110100000110110011100010111100110100111111000100101001010111100000000111111010111010110110001001111111100110011011110110001010010101010101010101111101100010001101010101001011;
#1 $display("%b", po);
# 1  pi=207'b010111000001000100100010111000101010110001010110110110000100000011011000111011101101100000101101100001110110000100101110001011100001011100110101101100000001111100011110110001111101000010110101000111010011011;
#1 $display("%b", po);
# 1  pi=207'b011101001100110111011100111001001111010011110000101001000110111001111101000100100011110110101001001110100110111000110111110001101010011101110001001010000100111111111001110100010111100001011101000101101001111;
#1 $display("%b", po);
# 1  pi=207'b011100001111011101010000111101001011101111000000111101000110010111100000100101111001110011101111011100000100011101101111001100100011011110110011011111101100110101011111010111100000011001111010111001110100001;
#1 $display("%b", po);
# 1  pi=207'b101011010011111110100110000100110101101011000011111100101100011101010001010100110101110001010000110010110110110010101100011100011110111010100111001011110011101010011001010100001110110001011010110010010000110;
#1 $display("%b", po);
# 1  pi=207'b011101111100010110011011101000101110000001001011110101000111100011001100110011000110010010011001011111101111100000001001111100001001100000101010001001100111011100101100100101101010101001111010110000100011111;
#1 $display("%b", po);
# 1  pi=207'b100000100011010100110010001000010000111000101011011100010010101111111111111100100011111010101101010110000100100110100010000011010001111111111000011110111111000101100110100111000001111100001000111111011010110;
#1 $display("%b", po);
# 1  pi=207'b111110010101101010010011001101111001100000010000100101100101000010000011000111101100011011010111011101010000100011011101111001011100000001001001110100010000110101100100111001011100001010001101110110101111011;
#1 $display("%b", po);
# 1  pi=207'b011110010101011110011010011101100101001010101011111110000011010111010100101101101111101011100000110101001111011111011011111001001111011110101000000010001110011110101011111100111110010100001100000010111101101;
#1 $display("%b", po);
# 1  pi=207'b100110011110110101110001100010011001000010101000011101110000111011110101111011101101100001010110111010110000101001011011101100111011000000110010111100010000011011110101111110100010001100110001001100110010000;
#1 $display("%b", po);
# 1  pi=207'b111000101010111110101110000100100000001001001000110100001010101011100011010011011100011001011010011011101110001001100110111010010000110010110110101100010100101001000111001101110100100111101000101111100100111;
#1 $display("%b", po);
# 1  pi=207'b001100110100010101111110011010111011100010100111100101110011010011010100101011110001101001111000101101100100110111011000100100000111010101000110011010100011000110100101101000001111111111010100011100011001110;
#1 $display("%b", po);
# 1  pi=207'b000011101010000001001101010101001011101010100000001010111001100011011100001010010111010000001011110010100010011100111000000000100011011111000000110110110001000001000010011101110110100110001100110010011001100;
#1 $display("%b", po);
# 1  pi=207'b101101000011111001111000010001101000101100000001111001010110101101110001010111111111010110111000110010100010001110010001111010011111101001100000100010000111101100111100000110000100111011111000001000010111001;
#1 $display("%b", po);
# 1  pi=207'b011000001101111101000011100001011010111000000110010111001001111110100010011011101000101110110111110101000000111011001001100110010100010110100111010000100100000101001101000100110011010100100011001010100011011;
#1 $display("%b", po);
# 1  pi=207'b100011101000011100101010101000001110010000101111111100010011110010010101100011101010100010001010000101001111111010000010101010000010001110010011011101011110110000000001110101001011101000110010111010100001011;
#1 $display("%b", po);
# 1  pi=207'b111000111100011011101100001110001111011111010010001110111111011001001011010110100111101100011001111110000100100000111001011001011011001011110100011100111110101010100110110101111111100110010010111100000110011;
#1 $display("%b", po);
# 1  pi=207'b011010110101111001001010001101011011100000001111111111011110010110100110001101110100110111010000001011011111010111111000010010001100110110010010010000000011110011111110111100010101111001101001010101010111101;
#1 $display("%b", po);
# 1  pi=207'b010100000111101110110101111110111010001111010110010100110010110001111101111110010101010001100101011001110010101110110111111111111111010000010100110010001010111010001110111010111111111000000011101011001111000;
#1 $display("%b", po);
# 1  pi=207'b110100100111110111001101101000110101101001010010111010100100111111000110000000101111011111010000101101010110010100101111100100011000010100011100100110011010100101001010011110101000010111110111000000001001010;
#1 $display("%b", po);
# 1  pi=207'b000010001010001001110000111010110001110100100000000011110110000101111001101010111011101110100000011001110011000000000001101000111011011010100001101101111000111010010110110000100101110100111111100001110101111;
#1 $display("%b", po);
# 1  pi=207'b011111100000001011111001111011010111000110011000010010100110011101101111100000100111010101000100000100001011110111100100011001110101000010101001111100111110001101110100010111101011100101010000011110011000101;
#1 $display("%b", po);
# 1  pi=207'b111000101110110111010000110111011000000001000110111111010011110101110110101110011011000111010110101100100000111001100110001011110011001101100100001010001101111110100110011000010111111110110010000000101000011;
#1 $display("%b", po);
# 1  pi=207'b101100011011101101001110111011011110000100000011101011001001110001010011001101100000110111011000111110011001100100100111011111100101110101110011100011000100101011110110100110101010000001000011110011111100000;
#1 $display("%b", po);
# 1  pi=207'b011100011011101110110010101101010010111010101010000001100001101111100110100010100101100000110000000011111000000010000010100010110100101011100000110011011101101000111110101111111000001101000110000101101001110;
#1 $display("%b", po);
# 1  pi=207'b111101001011011010110010011111001010000110100011100011100110011101001010001101011001010111110001101110001101010010010011100100111001101111100111110110101001010011000010000010000010111100101010001001111111101;
#1 $display("%b", po);
# 1  pi=207'b010000000101101011100011011110010101110110000110011001100000000001000000111011111101010010000001001100110101011010100101010100101111110100001000100011111010011101001100110100100111110010011110011010100110010;
#1 $display("%b", po);
# 1  pi=207'b001111000010101110010001010001101011110111011010010111000101100101100101000001010111101001101010011011000001101110000001000100011001001110000011010010000101010000101010011000100110101101000110110011111001001;
#1 $display("%b", po);
# 1  pi=207'b001111001001111101010101010010000110110000001010011011011110111010010011011011011001110100001010101000100101111101000110000101011001000101111100010000110000010101111000100101101001101100101100110001110111100;
#1 $display("%b", po);
# 1  pi=207'b110100101111111100001100101111100110010001001010000011100001011010001111101101100111110000010100010010010100001010111011000101010111010100001111001000110001001100101110101110000111110101100010110111010100010;
#1 $display("%b", po);
# 1  pi=207'b100000101011001011001111110101001010001101011010110101001011001101110100000010101111110101111110101010011100000101011001111100101101100110001100001011111111100011101110110011110001110011110100110010111110010;
#1 $display("%b", po);
# 1  pi=207'b001111011110110001011111100010101110000011000101111111111001110100001100000010011000010111111000110010011110100100111111000011011111110010101100100110100011100010011110110111100110111010100101110111011011011;
#1 $display("%b", po);
# 1  pi=207'b101110110010011101010011001000101110100011010101010010111001001100001101011011101011010111110011011111101111111100000111110000101111110010001110001100001011001101010101000011000110110101011011011110100101101;
#1 $display("%b", po);
# 1  pi=207'b011101101101011010011110011111011010010001001110110011100011100100001001010100011110111100110101101111101010100010100010110000010001110101001100100110111001011000010000000001100101011000111000110101100010101;
#1 $display("%b", po);
# 1  pi=207'b001100110001111100011111111100101100100000110110111100100101111101001010010100011010111011000100001101010000010011101010000000011001100010001110000111011111000001111110010101010011011011101110011011000001011;
#1 $display("%b", po);
# 1  pi=207'b010010001000011010101001111010001011000000000110111010110111001110110011011001011101100011000011011011000001110001000101001011001111010101000110001000100000001111000101101110101011111000101001100101010000100;
#1 $display("%b", po);
# 1  pi=207'b100011001100011110011000001100011101010010101001111010010011001101001001010100110011010101001100001110100111000011110111010110101111100111011111110010010110011110011000001111001010001000110000010000110111010;
#1 $display("%b", po);
# 1  pi=207'b111001110011000011010011110010111100011110010110111110100010000111011110111100110111101100100010111011010010000111111010000111100010000110011100011001101101011000101111011100111111100010001111110010110111110;
#1 $display("%b", po);
# 1  pi=207'b001001100111110110010100000111000100000010101011011010011010001011010111011010110111011001011011111001100011100001011001110001111110001001110111011010110101011111110100111110101101001111111011110100000000010;
#1 $display("%b", po);
# 1  pi=207'b010010000100101000001100111010101000110111001100111010010100001101010101000110000000011110000100010100000000110100101001100001010001000010010111010000110111011110111001100001110111100111100010011010110001010;
#1 $display("%b", po);
# 1  pi=207'b011101111110010100110011110101010011010010111100001111111101110111000011001100101111110110100101101101111001001000000111000010111101101100101101001101110000011011010110110000010111100100010001010001110001110;
#1 $display("%b", po);
# 1  pi=207'b000111111100111110011101010110000001101000000101010100011100101000111100000100101100101110011100100000101111101011110011001110111110011011111101100111000111001111111000100001101110000011110110001110100101001;
#1 $display("%b", po);
# 1  pi=207'b100010111100110101001110001101010110011101011111110110000011110001000000100110110010010111010010100100011111010111000001110010100010000110000101110001111110001100011111110111000110101110110010010001010010101;
#1 $display("%b", po);
# 1  pi=207'b011100001111110101101001011011101111001001001101111011001000101101100110101010010111001110100001100001101011110011011110010110000111101001110000011001000000001111101000010011011100101110001100010100100000101;
#1 $display("%b", po);
# 1  pi=207'b100101011011010001000010010110101011010000111000111101001101000110001111000000000111111110100101001001101100001100111110101101110000011000110111001111010110011001010001110110011010100110000010110111110000010;
#1 $display("%b", po);
# 1  pi=207'b001100001000111010010110011010010001000101011011110111110010101111010110010111101000011000111111100010000100011010111001110000110011100001001001111000001100110011001010000000010101111101010011010001001010111;
#1 $display("%b", po);
# 1  pi=207'b010010000011100010010111111011100101000010110110101100110100111010000110001000000101011000001111010100001100010111011000001100101101001011110001000011011010010010001000011110001111111101111100000111001001110;
#1 $display("%b", po);
# 1  pi=207'b101110001001001011111000100001111111011100110110010001001001110100011110000011011101010000110000000010010000011100101000111100100010111110101011011011111110010001110101001110100111000110010010011001111011010;
#1 $display("%b", po);
# 1  pi=207'b011111110000100001101010110011101011011101110001100101000101101111111101000000010100101011111001100110111111111110011011111010001011001100100110101101011010010011101110011101000101101011101111101011100001011;
#1 $display("%b", po);
# 1  pi=207'b010101110110010101101100011000010010010111111001110001111001001100001101100010010111110110111010001010101111101000100101010000000000000111001100101101011110110101100000001111011010111101111111111001010010100;
#1 $display("%b", po);
# 1  pi=207'b011110101001000011000110011100111100101111111011000011101100101001010100101100100000000000100010100000101110000011101111111101100001111101000100100000011001101101011010011101011101010011100111000010100001000;
#1 $display("%b", po);
# 1  pi=207'b101110110111000111111100001110101111011010100000111111001100011111100100111100010110000111010100110110000010011011001110110110111110100000111010100100100111110000010100010110100101011110100101010001011100110;
#1 $display("%b", po);
# 1  pi=207'b010000101000101010110001011000010001110110000011111100101001010011100101011110001001101011011100110000000110000001000111100110011010101110100010100010101100110001100010010111100111010111000010011000110010100;
#1 $display("%b", po);
# 1  pi=207'b000010001011101110110110011110111010101111110001001000101001111101101101001110001100001000110111101011110011000101110000000000100111110111110100111101111100100100000101100000001100111110011111101000111101101;
#1 $display("%b", po);
# 1  pi=207'b000000111010011011110111101111111010001100000010000001011100010010011100111100001100001001100001010010000000100101001011101011111001000100001001111101100000011011011111001101000010011001100100010011001100101;
#1 $display("%b", po);
# 1  pi=207'b011010100000000100001001101010010011100111010101000110101001100100111101111000100100100100011100000110101111110011011100111001011111111110111111010000101100111111111111010010110011001110111110111011110011000;
#1 $display("%b", po);
# 1  pi=207'b000111011100011100100110011110001000100100100010000011001011101101000010101111010011100101000010111010101100000111111101101000000000100001000101110000001101110011110001100011011010011001110100101111011000110;
#1 $display("%b", po);
# 1  pi=207'b110101101101100100111110011001100100100011100111101000110011010010111111001100101011111011001111001101010100010111101000010000101001000001101110000000100010101100000011011000111101000011010001110110100111100;
#1 $display("%b", po);
# 1  pi=207'b000101110000010100000001111101101111100011100010001010101100001111111101111000111000100110001001101101010110000111101011001110011001101111010000000011101111101000010001011000001110001000101111111111110000010;
#1 $display("%b", po);
# 1  pi=207'b101111011011111000001010100000111100110100100101101101000101011001100011111010111101010111100101101010001001010010001111100100100011011100010110100011001010100111101100000110011000010101000101001101101010000;
#1 $display("%b", po);
# 1  pi=207'b111001101001110110000100111101001101001001000011010001010011100100111111011001011100010010111011111100010111010000001011001001010111101010110011101010010111111111101111100100100111101101001101111101000110111;
#1 $display("%b", po);
# 1  pi=207'b010110100001110100001101100001001000110100000110011110011100100100110110010100000111010111000100111100101011001001101110011001100000100010110011011111000100110011110110010110000010101111101111101000110111011;
#1 $display("%b", po);
# 1  pi=207'b101001110000110001010100101111100010110111010100011001110010100001100110001010111100100000011000011010011101010110000111010000011010010101011101101000111011010010011100111001111010101110011110010001100101101;
#1 $display("%b", po);
# 1  pi=207'b110100110011110110011110011111101100100110011110110011010101000000001010100011100000011001110001010110101101101100111100001011100011111110010010011110001100110100111101100010110010010010000110110111011110001;
#1 $display("%b", po);
# 1  pi=207'b000001100001111001111011101111101111000010001010100110101001100011101110111001100010111001000001011111010001100101101010110111011100000001101001001110000111010010110101001000011010000010001101001011111000011;
#1 $display("%b", po);
# 1  pi=207'b001110011000001001011100111111110000110001111101111000110011000100001011011110111101110011101000100001011010110101011010111011011101111000011001000111111110101000110001101011101010100110101010000010111000000;
#1 $display("%b", po);
# 1  pi=207'b101100110101000010000100000001011110001111110111100000101001100010110101000111011011000110110001110100001001111111010000101111101101100110000011010000110001100010101100101101110011110011111000011001000101010;
#1 $display("%b", po);
# 1  pi=207'b011010100010011011010100101100000111011100101000101111010011011001001101001010010011110001100100001111111011000100011100001010011111111111101010001110000110010001010110110011010001000001111110011000000110101;
#1 $display("%b", po);
# 1  pi=207'b001101000110010101000100100111010001100010101011101001000001000011010001001111111011011100001001111000111000110011111110110111001000001101110111101100100111101011100010011011001001010111001100011110101100110;
#1 $display("%b", po);
# 1  pi=207'b010000101101100011101100100101011100111100001000011001010010011001001101001111000110101011000010101100100011011100111100001101100010100100001010110100100100000101100110111111001010101101100010000110101000101;
#1 $display("%b", po);
# 1  pi=207'b010001000011011010000101010001111000111111011110111010011010100101100000110000110011110011010010100000000101011000101101100011001011101010100011100111000011011101011001100110100111010100010100000000100100000;
#1 $display("%b", po);
# 1  pi=207'b110100111101000000101000110011000110010110101001011010100010101011100101100000101011110110110101110111001111010100101101000000010111001110000101001000010001111101101111010111110000011010101001111111010001101;
#1 $display("%b", po);
# 1  pi=207'b100111011101100000111101100110010100111111101001000001111100000101001001000100100010011000101000001001001011100100001000010010010000110110011111011011001101100100110010101101000110101110111101111110001001001;
#1 $display("%b", po);
# 1  pi=207'b101100110100101101110101111110010100111010101100101001100011100011110001001110000110100111111000011000110011000110011101011101100001111111000000110010001011011000000101111010111100000011011100011100101000010;
#1 $display("%b", po);
# 1  pi=207'b001111011000100100110110110010100001111011101001011011011100110101001011001100010000000100100110110011100010101001100101111111011111101001100110110000000010000101101111000101011101010000100010100111111111110;
#1 $display("%b", po);
# 1  pi=207'b101110110000100110000111000001111011000001001101011111111111100110000101101000000000010011010100011100001001010011111001101001001111110010001000110101011011001011010111100001110101110011010010101100001011000;
#1 $display("%b", po);
# 1  pi=207'b011001100110101111100100010010010000011000101100001100001111110111111011011111100101000111100010111110000010011110100000010100001110100010000011001011001011101111110100101000100101011111011010000101001111101;
#1 $display("%b", po);
# 1  pi=207'b010101100111111100111011111111011000101000111110111011100011001011011010110001010010111010100111010001100001001011011110110111011110101000101101001110011001111011010101101100100001111010110111000110101110011;
#1 $display("%b", po);
# 1  pi=207'b101010111000001001010100011000001111000010100111001111000010100111000101001101110011100101110000100000100000101111111111101011110111110011110111111000100110110101111110000101010010011011001100100110100110010;
#1 $display("%b", po);
# 1  pi=207'b001000111111001010111100110110000101011010010101101101110101101101111101100011011101100010011011001111001101001110000101101111101011111111101001011010010100000111001100011001111110011110001000011100010001111;
#1 $display("%b", po);
# 1  pi=207'b110011011110011011001100110010111110111111110101011010000001111111111100111001011111111100111010001001100011000101001111001110111101111010000100001011011001101110110001110110010011001010010100011101001011100;
#1 $display("%b", po);
# 1  pi=207'b111111110111101000111111000100110110101101111000001000001111111101000000010011001101000011101100000101100100000100111000000010000001101111101111101001010001001010001001101100101101100100110000110001101000101;
#1 $display("%b", po);
# 1  pi=207'b010010010110111000011110011011111001000001011111101100001011110000110110000101011001110000101101011010010000100001010110111011110001100101100111001001101110011110010010111101011111011011001100011001101000111;
#1 $display("%b", po);
# 1  pi=207'b000111011101011111100000110110110000001011111111010011111010001111110110100101001101110101110011010010111100000111111100011010100000000101100000011000001110111110110110101011100001100101111000001100110001110;
#1 $display("%b", po);
# 1  pi=207'b000100011110110101110100011110010001110010011011111110110111010101010000001101010100000101101000011111110011010011011111110111110001010001111101111010001011101100011111111110111110111000101101110101000001110;
#1 $display("%b", po);
# 1  pi=207'b010101101111110100010110101010101110110000110100111000111100010011001110101001011101001110001010001100101100010111110111111001011101011001111000101001011100101010000010100001100110011000101010000010000010110;
#1 $display("%b", po);
# 1  pi=207'b111011101001110111100110011001011101011110110011110111010011001100000000100100011001011000100111100011001110010110111110010101100111011111011100111110011001101100010101111010001100001010011000000000001100010;
#1 $display("%b", po);
# 1  pi=207'b000110011101110110010101010011111000100110101000010011001100001010001001011100100010100111110000101001001110101011100100110100011001111011000100010011101101111000111010100010010111001010111111001101011111110;
#1 $display("%b", po);
# 1  pi=207'b010001001001000010100101101011111111110010010110110001111011100100110010110110001110100111101111100111101100110111010001010000011100000000010011011000001101100011001101100001010100100100011000001111100000101;
#1 $display("%b", po);
# 1  pi=207'b000010001001000111010100000001010010101001100011111001110001110100100010001011000110001001100010110001101001001010111011001111111101110101111111011001000110011111000000101011001011100110100101111000001101100;
#1 $display("%b", po);
# 1  pi=207'b000011011111000110010111000111110010010111011001011110000100110001110101011100011001000110100111110000010010000111100001001010101011011010011000010101000100111011010001000111010111010111010011001111111111011;
#1 $display("%b", po);
# 1  pi=207'b001000111100011110101111000111000100111101001011010001010010010001010001110100010100000101010100011011001100000111010011101110101101100000011000010011000000100011101111100001111111010001111010011011010001011;
#1 $display("%b", po);
# 1  pi=207'b000000100111101111110100100110110000000111110010110100110110000110110010111000110011011110010100100111101100101101000000010100010010001000100110111111110001001001001011101111000110000010010110010001011100111;
#1 $display("%b", po);
# 1  pi=207'b010001001101100000000011010011010001100111011011100001100101100000110111011100111010000100111010101001000000001110111001100100110110110011111001101011001110000011010000010001110011000011100111101000111100000;
#1 $display("%b", po);
# 1  pi=207'b011000111011000010110010011111001110011111111110101100111110101000011000111011010110111000011011010110111010010001001100010100101101001101111011100011010110000001110110100110110111101100101000010001100100110;
#1 $display("%b", po);
# 1  pi=207'b111110001111111000100011110001100001101011110101010010101111100111101111001001011100000010101001101001010001100010100000000001100010001000010000001000010111100111010110101010110000010001111001101101100101110;
#1 $display("%b", po);
# 1  pi=207'b110110000000010110000101111001110101101100110101011111100001000001011101011110001000000100000010111011100100101001100001011100010000010011111100011111010110010111111011101000111000011010110001010010011011001;
#1 $display("%b", po);
# 1  pi=207'b101110001111001011100000101111010001110010110100101011100110000001111101011000010110011100110101101100011101010110111100100101110000010101100110110011001000111001110101100011000111100100101011100111010000010;
#1 $display("%b", po);
# 1  pi=207'b010111100010011010100111110011100011000110100010100110011101111010001001100001100101001101000111001111110011000101001100011100100001010100001111100111010010101000010010100101101101001011000011100100111010101;
#1 $display("%b", po);
# 1  pi=207'b111011110000101110111011111011011110001010011000010100001100111111111011000010011100000010010101100110000101110110000001101011001010011001111100110100011011101001010111011110100101100111111100011100101111011;
#1 $display("%b", po);
# 1  pi=207'b110110110010100001010010010011001001100000001000000111101001110111011110101110000001001110010011001110010010000110111011011001110111001011001011100110111010000101100100111110101100111101100100110000111101110;
#1 $display("%b", po);
# 1  pi=207'b010010001100001100000000001100111100101001010010110100000110000101101011011100000001101011101011100001000111001101010001010101000100000001000100100110110011010111010100001000101001100101001100001110001000000;
#1 $display("%b", po);
# 1  pi=207'b101100111010011100100001110111101001101001110000110101001111101010011101100001010111110101101000001101011101011001001111101011110100110110110001001010001010011000000010101100101111011001101000010000100111110;
#1 $display("%b", po);
# 1  pi=207'b001111001011001001111010111111010101101100000101110111011110111001100111010010111101011111000001101011101000101001000011010101100000001101111101111110001010100000101011111001011011110010100100011111000001101;
#1 $display("%b", po);
# 1  pi=207'b010011100010100101100100101001100011010011101101001110100100100000110110101110110000001000101011011100110100111111000110111001101111011011001010010011001100110111101101010100010110010111000011111000011010110;
#1 $display("%b", po);
# 1  pi=207'b001110011011010011100110001001100110111101111110100011100110011110011100001110000101011010000111010011111100000001110001001110010011000101100100101011011010010101111101000100010111101010011111011000111101101;
#1 $display("%b", po);
# 1  pi=207'b101000000010010101100011100001011011000100111011100100110000100010001101111011011000111001000010100110101000110110001011001101110011101100100110101001001000101100101101010100111010000101011011010101110110010;
#1 $display("%b", po);
# 1  pi=207'b101101001011011110011010100010011111101001111101111010100101011101100010100000101111111110000101110001001110000011101011001110010101101001000000101111001001110000111101111000001010101000101111011101001010100;
#1 $display("%b", po);
# 1  pi=207'b100111001000000000001110111011010001111011111101001101001010100000100100110110111010101000001000011011111110110101110010011000100010010100011000000101010110101110001011110111011100001001010001011111000111011;
#1 $display("%b", po);
# 1  pi=207'b110111010111010010110001111101100110000110001111010101010110001000101010000100111101000011001010110111110010111000001110010010010110110001110100011010101000010011001101011011101100111100101101010110011111111;
#1 $display("%b", po);
# 1  pi=207'b101001111101101011000110000110100001100010011111011111111011010001101101001001001011000010100010101011011011011111000000111111011100010110001010010011011000001000000011010101000011101100101010011011100011100;
#1 $display("%b", po);
# 1  pi=207'b100110111011010000110000000110110011000010111101001000001000010101111010011101101000000101010011000001011100100111011011010110100010011001011010111101111010000111111011111001001110111100110111001101111100010;
#1 $display("%b", po);
# 1  pi=207'b101100110010000011100011011010011000110111101111011111000101010111010101010001001101110110010111111000001011100001000011100101101110001010111101001110000100101100001111011100110001111010111110001001001001101;
#1 $display("%b", po);
# 1  pi=207'b100010100100000101110000100110100111101011001000111100110011010100110001010001000110101110110011111101110110111011011011110101011001110110111011000000000010101111011111100100111001001010100111001010010000111;
#1 $display("%b", po);
# 1  pi=207'b111111110100111101011100111010010011000100010101011010100101101011001011000000000001110101010011001000100000000100110100100010101000101101010011001011111111011110000010100000011101000101000011000110100000001;
#1 $display("%b", po);
# 1  pi=207'b011110111010010101111101010001111101100000000010000000001100010010111111011101011101110011111110001110000011111000010011010101110101110101110100111000101010100111100010010011100010001110100001100101000101011;
#1 $display("%b", po);
# 1  pi=207'b000010101110010110001000111101100010010010011101000000101111010010101110010011001011111100000010111101001000111110100000010000111100110001011101110110010111101111000101000100110011010111010100000011001001111;
#1 $display("%b", po);
# 1  pi=207'b110111100000111001101010000111011010011111001010000110001110100010001100110111111100001111110001100110110110001001001101100101001010110111110100011110101001000101110010111101010111000011010011101100110011101;
#1 $display("%b", po);
# 1  pi=207'b111110011000010100010001110010001101000101111011111101011000111101110100010111011100111000111100111111111001100100110001101100110111000100100101111000011111100010111111110011010110010010100111111100100100011;
#1 $display("%b", po);
# 1  pi=207'b100110101111100001111110001011110100000010110011111010010000111110110001101110000001110100100100001101111101010011110100000011000000011111101001011000010010011010101010111101101110001111011000011000111010101;
#1 $display("%b", po);
# 1  pi=207'b001111101001100111100011010100100001100000101011111100010101000001111100010111111001011010111101111111110110101000011011010001000111100000111110101111110110010001110001001110011110011000110111100101011110110;
#1 $display("%b", po);
# 1  pi=207'b010110011111000000111111101000100000111101010100011100011110110101000100000101110101101100000111000111011000101000101101011101000000000110100111010101101000101001000111101010011100100110010110110001000110000;
#1 $display("%b", po);
# 1  pi=207'b111011100101010010010101011100111101101100001111000101100110001111100000000111111000011000010010110011000100111001101101101101001011100111100110011000110010011100010101111000010101011101011011010110001110110;
#1 $display("%b", po);
# 1  pi=207'b000001000000111101001111000111010000111001110001000001001110110111101000010100001000100100101011011001001100010001011100110010110010001001001010011110000010100111011010101000100100110011110101111100101010101;
#1 $display("%b", po);
# 1  pi=207'b101101000100010110101000111001000111000110010101110110011001110011001011010111100100010010000101011000101110111001110001100001110110100010010001011111110101011011000001100011010000010101111010100001011100010;
#1 $display("%b", po);
# 1  pi=207'b101011100110010000101110000011101110101000010110100000100101101011000011010000010110101000111010000001000001001000110000100011000011010000111011000111001111001010010110111001011001101110110000101000110101000;
#1 $display("%b", po);
# 1  pi=207'b110001010101010001010111000100010010111111100111001110100000110011101000000101011100100011111111111000100001110010101000100000111110011010101100111100100101001010011101001011110010111011010001111110001111110;
#1 $display("%b", po);
# 1  pi=207'b010111110011011101101111111001001000110101000011001011100001111010000001100110010010011011010111010110001000101101101100110001001111010000111000111100111101011101110101100100100001110110001011101011001100011;
#1 $display("%b", po);
# 1  pi=207'b111010001000010101110101110000001111110110001110010111011100000001100101000000011010101011000011001000101000101111101100001100101101110010010001000101001101000000001010010101010001111000101001101010111111100;
#1 $display("%b", po);
# 1  pi=207'b010010010000001111111101101100010111100011000110111111101000001111000001111110001111000011111101001010000011001101100111001101011100101000100001111011000010110100010101110100001000111111110110110001100011100;
#1 $display("%b", po);
# 1  pi=207'b001100110010001011010101111101101101001000100101100011101000100111011101110110000111010110100001100100110000111110010001111111010111010000011010101011010111111010010001111101100001110110010111001110111000010;
#1 $display("%b", po);
# 1  pi=207'b011000011001010111011101111001111111101011100101011010110111001010100001011100010000000110001111111011111011001010100110101111011001100000100110000001100110011111011101111101110110001011111011100000000111011;
#1 $display("%b", po);
# 1  pi=207'b011111101001010111000110100101010100001000111001110111100110001110001100011110010001101000001000100001110010010100111101111001110110110000001111111100010011101001000010101110001011100010001111110110110010000;
#1 $display("%b", po);
# 1  pi=207'b011000111100001000110110010101101111111010111111001110100111000011011000101100100111101001101011110000000000001011000111001110100011111111100111011000111100101110100000110111001100000000000111001111010101010;
#1 $display("%b", po);
# 1  pi=207'b100111010001001101011001010001010010111000101110100010101101010111100001101011101000100100111111111010011100011101111010101100111000011010000000110000110000011010111110111110000011000011111100100101010110010;
#1 $display("%b", po);
# 1  pi=207'b110001000100000111000010000001001010110001110000000000010110011001101100100010011110001110000100100110100010100101010011101101011100001111010111010100000001100010111101110010101111100011110110010001111010011;
#1 $display("%b", po);
# 1  pi=207'b110011001000010100101000000000010001101000001000010000100000100001110010001111011000100001000010011010111111100010001011101010111000100011001110101111000011011111010101111001100111010001011001001001010011010;
#1 $display("%b", po);
# 1  pi=207'b100000000110110110000010110100111010001101101011011110010100110001101001110111000001100100100011101101011111000111101100101100011110111100000010001001110011101011011111000100011001000101101000011001101001110;
#1 $display("%b", po);
# 1  pi=207'b010001101101111000001101010110110001001000011101110000111100011000101110101100100010011101110111101100100010010110001000011001010111110011001000100011011010101001010110101001111110000111010000000101011011011;
#1 $display("%b", po);
# 1  pi=207'b000010001010101010111010110111000110110001011111110100101000101001110111101101011001000010110000010001111001001110001101010111000011111101101001011001001101011101101111001011000011101001011101001101101101101;
#1 $display("%b", po);
# 1  pi=207'b010110010001111100101000000110110011110001111010001010100111011101100110100100111101001011101110101011011111000001101110010110110101001001111010010100001000100011010001101100000001000001000000011011000111000;
#1 $display("%b", po);
# 1  pi=207'b010010011101011100011001001010111010110100010011110101011100000100110111010110110100010100011011101001110111110001111100000100100101110100111101111001000000101001100101110001001111011001011011110011110001001;
#1 $display("%b", po);
# 1  pi=207'b110110011101010001011101000011101111010010001010010010010001000101101110010101111111101011100010001000111000110110111100001101110010011001100101011100010100101100000111111011010011101000001011100110110000011;
#1 $display("%b", po);
# 1  pi=207'b000110000110101100110010100011010000011011101000010100000001100100001111001010010000111111101011000101110110010010101111001000100110000010111010110111011010110101010011110000001010110010111001010000100011110;
#1 $display("%b", po);
# 1  pi=207'b001111111010111111110011110010111101111001001110011100100110100010010100010110001010011010100100100110001011001001011011000011010111101010000100011011011111101111111111111110010110010001010110110111110011001;
#1 $display("%b", po);
# 1  pi=207'b010100111110011011010111001010000110110010001101010010101010010010011001011010111010111001100100100111110110100111000101011110011111011110100011100100010101101000101000111110111110110010000100010011110100111;
#1 $display("%b", po);
# 1  pi=207'b010010111000000100000000101100101111011011000110111100001011011101010011101111101010001110010001011100100001011111110101000101100101110000100110100000001010011011010010100110010111111011110010111010111001100;
#1 $display("%b", po);
# 1  pi=207'b110100011101010111001100010100011001000111110110100001001001011011000001011100011000111111011000101010111111111100011100110110110001011100011000101001000100011100111110000010101101010101000001110001001001010;
#1 $display("%b", po);
# 1  pi=207'b000000101000001001000101100100010111110011011100010000111101010110111010110111000001011011011010001110111001000111011010001001111000010111010111111111001000110001000101110001100000011100110010101110101010111;
#1 $display("%b", po);
# 1  pi=207'b110001001101011001000111001011101111001100100010100011000110110000011001110011111000101100111000111100011111110011101011001110110101010010000010110001101000101100010101110011101000010101110110100010010110110;
#1 $display("%b", po);
# 1  pi=207'b011010010010111001101101011000000111010101001111011101100111100100011101011010101010100010110000011111001000000010011010111001111010011111110111110000000000110111111101011101100011011110011001100101111110111;
#1 $display("%b", po);
# 1  pi=207'b111010100011000010110000100101100100101111101011010100011001010110001111101010110011001011100111100101010010010110110010000100100101000111010110010110001111101100101011101001100001101100100000100011001110011;
#1 $display("%b", po);
# 1  pi=207'b011100010010011001101001010011111101100111100011111010010010000110000100011111110110000111010110101000001110001001111110010001111100100111111010100110010100000110000000111011110111101110000110100111010110000;
#1 $display("%b", po);
# 1  pi=207'b101011111110100111001000011011001100010000100100000000110000000011111001000000111000111110111101110010000101110011010001001101011010111100000010100100100001011100110101100101101001010111101111010000100101111;
#1 $display("%b", po);
# 1  pi=207'b101110110000010111101011000011100011100101001000010000001010110110001100101010111111101100111110101011111101001110011110011101010000111101100110001011100100111010101001000110000101101111011010111001001110011;
#1 $display("%b", po);
# 1  pi=207'b100010010110100111011000100011111110000000001010110101010110110011111010101110100000011100100001011111111010110100110010010100100111000001111001011001110010101000101001000110110010010010011000010111101110110;
#1 $display("%b", po);
# 1  pi=207'b001110110111010000100010001011011110110100110111100001001000111101001000100101001001111100110011011000111100100110011111011100100000000111111100011111011010100101101101011111110101100001110110011110001001100;
#1 $display("%b", po);
# 1  pi=207'b000010111101111100101101100100101100000110010101100101101011001111011010111001001010000110010111010101110111001001101010010010000101010100000101101111111000001101110000010001111110001111101101001101100100011;
#1 $display("%b", po);
# 1  pi=207'b101100110100010010111111001011110100011011101000011110010111001010100011000000000110100011001001010000110001111010001110010111010110111100101100001010101111001000001010000001010101101001011111100100101010110;
#1 $display("%b", po);
# 1  pi=207'b101010000001011010010111000100110110001001100000001101001010101011100010011101111110101010110111000110111111101000101110010010100001110101111000111010101100110111000111011001101011101011100011000101011111011;
#1 $display("%b", po);
# 1  pi=207'b110100000011001000100110111111101111011111101100110111110110001010100101110010001101101001110111000100101101011011111101011111111110010101011010101001111001101011001000001111101001000111001011000100101010111;
#1 $display("%b", po);
# 1  pi=207'b000101001110001001011100110100100100000001100000111111111001001110010100000001100100000001110011001100001101011101011101110001010010110110100001000111001001110011111001010000001011101111001001001110011000011;
#1 $display("%b", po);
# 1  pi=207'b011011011110001000101000001100101110000000101101000011100010000000000001111110010000110101111001010001111101011001011000101101100100111001000101101101110001110110100100101011110011011001101011110101001001101;
#1 $display("%b", po);
# 1  pi=207'b001111010110111110100110010010010111110010001111001101100110100010000110110011000100011011011010111101101011000111001101001010000000101010000110110100100110100110001100000110010111110101101001111001111110111;
#1 $display("%b", po);
# 1  pi=207'b011100001010110010100010100100000010010110101111000110100000100001011110100110110111000000010110110100010111100011100010010110010110110111100011011001100001111111010111110111010011111110100101011010001110101;
#1 $display("%b", po);
# 1  pi=207'b001100001110001010111111100111000010111011000011000011100001111011111111010000011000110101100011001010011101001100000111011100001000011100011100001011000001010011111001010100101101010101111001111010110111101;
#1 $display("%b", po);
# 1  pi=207'b000101110001101010101101010000011101111100111001010111000010010011011100101000001100111100111100001000101111001011010111111011001000111101100101111101001001001011010001110110001111001100001011110010111100100;
#1 $display("%b", po);
# 1  pi=207'b000010101100101010001000110111010011011001000110011110101000111110000110011100100001110111111000010000100011111101000000101111000100001010011101011100001111001011100110111110110000011010101101000011101010110;
#1 $display("%b", po);
# 1  pi=207'b101001000111111000101111000000000000110010111000010001111111101110011001111010000010010101001001110111010011100000110111111110110000101000110110111100101110111011101110010110001110110001011110111110000110101;
#1 $display("%b", po);
# 1  pi=207'b011111011010111010110001100001011101111000000000000011100001010101001101010111110011100011101110110101000010101100111000111110111110111100001001101111110010001010111111010010000100000010110000001101011001111;
#1 $display("%b", po);
# 1  pi=207'b110101100000000110111100000111111111001110011110111100011111110110111010010110001100100001011000101001001000100100111111011000110000110100111011011010000101001101111111001111111110100111100011100111010100111;
#1 $display("%b", po);
# 1  pi=207'b010000101100110110101010011100011001110111110110001011100011001011001011101101101110110011111000011111010111011000111101001000000111010001001001010110101100001101100001111100101111001101111000011111001010001;
#1 $display("%b", po);
# 1  pi=207'b110000111011010100101011100100111010101110011111110010011100100000111100101011100101011010001010010010101110000000011101100101000111000011100111011000001000100101000110000101011100100101001000111101001110001;
#1 $display("%b", po);
# 1  pi=207'b000000000010110000110010111010111111110100100100110010010110101100011011000110001111001010010001001111011111111110111110010011001111110110000001010010100010001001100100011011101111010111100111000001100011000;
#1 $display("%b", po);
# 1  pi=207'b100010001110101101110110000011100001011010111111000100101110111011010111010011110111000000010001001100001000100010101010001011101110100101110011111000101100111110010110001100111000100010000011000011100011101;
#1 $display("%b", po);
# 1  pi=207'b011010011001100001001101111010111110001110100100100110110110110111011101100100000000101111101100100100100101101001100110101101101101010010101001111011111100000110001011011001011010001010001101100111100000100;
#1 $display("%b", po);
# 1  pi=207'b011110001111011110110110111001000000011000100110011110001011111101010111010001010010100000110111101001100010010100011111100001010000111101111001010101101100001110011111001000011110100101111010011100011011001;
#1 $display("%b", po);
# 1  pi=207'b010000001110010010111000010000111001010100111110110010001111110001010101010101001000101001010010100110111100110010101101001001110001100100111001110111101010000100111110111100111111101001101010000011111101001;
#1 $display("%b", po);
# 1  pi=207'b000000000110101111000100111101000100111101001101100001111101110111100001111101110000111011111110100110011001111001011011111110010000011000010011101001110001000000111001100010100100110101000000001001101100101;
#1 $display("%b", po);
# 1  pi=207'b100011110101000011001000101110101000001011001001110011101110010011100001001010111001010100010010010111000111000011111111111010101001100001100010010100101010000000100010000010000100001111110101011010100011000;
#1 $display("%b", po);
# 1  pi=207'b110000011011011100011010001011000111101111001111010110011010001000100110110000010100110011111111111111010000110111100010001000111110100010110010010001011000101110100110011110101001010001110100100010110110010;
#1 $display("%b", po);
# 1  pi=207'b000110000110101111000101010111011110010101000010111101111111011011011101110000000011101100011111110110100001111101110000100110011000100011011000101001011010010001001010000100110000001100111001101011110011101;
#1 $display("%b", po);
# 1  pi=207'b011010100010101111010100010111100010110111111100110101001110010101110001011101110111111000000010000011000111101001100100100000101011001000100101100001000101111100000000011100101010000101010101000000110100100;
#1 $display("%b", po);
# 1  pi=207'b010111110101000000010001101010010001001110100111110010101111001101001110101011000010111000111001011111011000111111111101110100000111001110010011100001000000011010011110011101010101111111100101011110000101001;
#1 $display("%b", po);
# 1  pi=207'b001000110010100111011001011101101100100101010101111101101010110011010100010110000011010110100011111011010011111111011101110100001100011100000101011001110110001001111011001110101110000000110100111100011111111;
#1 $display("%b", po);
# 1  pi=207'b100111101010010101001001011011000110111010001101100110111110110000011110010011100011000100010010000100111000111100111000110000001111010111111100100111000011110000110111011111101001011001000101110000000110110;
#1 $display("%b", po);
# 1  pi=207'b110001001001010000010011111101001010001100010001110101001111100010010011110010101100111011100111001000100111011100110101010101101100010100100001010111000111100101000110110000010010011100010000011110001101000;
#1 $display("%b", po);
# 1  pi=207'b011001111110011111001101110100101000001110000110011010011001000011000000001001011001011011100011100110010110000011000011010100100100000100101001110111110011010001010100000100000001100001010100000000110110000;
#1 $display("%b", po);
# 1  pi=207'b110100111010111010100011011010001100011010101110101000011011010111001010111001110001000000101011100000100011110111011111101111111101011101011101101011100010100001110010111101010110111100111110001111111110100;
#1 $display("%b", po);
# 1  pi=207'b011110111011001010101001011010011000101000101000110101100000010100010001000111010110000011111011001011101111011111010011000001000111110111100000100111000000000000100101100011010100100101100111100011111110011;
#1 $display("%b", po);
# 1  pi=207'b110010010000000011100011101101101110001010111000111110101000110010110011010011000110011100011110100111000001110010111111100011100101101000011100111010010011010001101000111111111111101111001101010000100001010;
#1 $display("%b", po);
# 1  pi=207'b010001010000010111100011110101100011010111110001111101101100100001000011000111001111010110010110011011100110010111011011011010100000000111100010000010100100110110110111101111100100110000110111010000001000000;
#1 $display("%b", po);
# 1  pi=207'b010010010110101010011101110001001110011001010100001110001110111101111000101111100110110101111101111011011101010110111001110010110011011100010000100100001111100001010010111010011111001110000111000101010001100;
#1 $display("%b", po);
# 1  pi=207'b000001110101111111101001011101011010010011000111010010111011111101111000100101000010000010000011010010110101101101001010000100110111110100111011011001100110001101101111111100011000101101000010010010001110000;
#1 $display("%b", po);
# 1  pi=207'b100011001110010011110101000000110101101111000100001001110110110001101000010111101011011101000100010000110110010011001001001101000011110111011100100100111111110110010110010111111010101100011001000101010111010;
#1 $display("%b", po);
# 1  pi=207'b010001010100010000110000111000000111001010000011100011001100110111010000011011001100111000010010011010110010110011110100110101100101111101101110011110100000100010001111101110111010000111100111101011011010001;
#1 $display("%b", po);
# 1  pi=207'b011110111010010111100100011010110101001010110001010011001100000000111110100111000001000100100000010000111101001011101000100010000001010100000011100100011000111001001101110100110111001100101010010010110111010;
#1 $display("%b", po);
# 1  pi=207'b010111011111011100000000001011111110110101110110011110110001110110011011000011111000101101010001101101000000110000101111010010111001010011011101001101101111011010011110110000100111101011111011010010010100111;
#1 $display("%b", po);
# 1  pi=207'b000111111111101111101110111011000101101111101111110110111101011110000010001000011010001110001011111101001101011011001010101100111100011110001011001011011000000011100101010110000100010000001000110000001010010;
#1 $display("%b", po);
# 1  pi=207'b011000101111011011000001011101100001111101100111101110101101001111010011100001110100001000000010000011110110101100010100101001101001001100101010000010000010000000001010010000000000000000101001001001101001010;
#1 $display("%b", po);
# 1  pi=207'b101000111001010000000000101101101001100001111011111011000101001010011101000001111101100101110111011001010111001001000000010110001111110011011010010100010001000000101111111011110000011100010110010101011001001;
#1 $display("%b", po);
# 1  pi=207'b011001011001100001010110001111100110010110100011011011100101001010100000101111001010100110011011110010101111111000010010010001011100000101001100011111011111010001100000100101101111111100000010000100111111110;
#1 $display("%b", po);
# 1  pi=207'b100011000010101111010010101111100000010110011000100010001000110100111001101100110011001101100000001111010011001010011000001001010110100001010011001110000111000011100010100101010001111010100111011100010101001;
#1 $display("%b", po);
# 1  pi=207'b011001111111001011111010010101011011101110100100000001100010010101110100001111100111011101101100011101001101110101001111001110111110101010111110001011110110111100000101011010110111010000111000100010111100011;
#1 $display("%b", po);
# 1  pi=207'b110001010110000111101010000111100001100111000000101101111010100000101000000001010101100100010101110110001001100010000010000110110110100001000101011101000111111000111100110010100111011100000100010110011111010;
#1 $display("%b", po);
# 1  pi=207'b010011000111111110010001000111011110000100011110101001000000110111011110011110010000101110000001001010001011101000010111100101001001110100110110101110110101101111110111100000010110010110101101001011100000110;
#1 $display("%b", po);
# 1  pi=207'b111111011100011100100110111111110110010111111111011110100100100111111111111100001100110001100110111001101100011100101010100111101000110111001101110000110100110100110011011010001111111111100111100010000111100;
#1 $display("%b", po);
# 1  pi=207'b000101100101011011101000111000000100111110101111100000100110010101110011011111110011110001101010110000001000100011111000111010101001010011101010001011100000000110101001000110100110101111101111010001111111111;
#1 $display("%b", po);
# 1  pi=207'b001010000011100010011111001011001010011001100110010111110011010001001101101000111100001011000111100101010101100101000000100000111110110110111111110001101101101101000101001100001100011000100101110100010110110;
#1 $display("%b", po);
# 1  pi=207'b000011011011001010011000110101000010100100111011000110001101111011010011011110100001001101001000011100110001011100010111110000010110110001001111011001111110110110011001011101001011111101000101101001100000000;
#1 $display("%b", po);
# 1  pi=207'b000000011110101011111111111100100111000001010000010100101011101000000101111110111100110010111111011111000001000100001010111110101101011100101000001100100101010001010110101000011110111010001010000111100111011;
#1 $display("%b", po);
# 1  pi=207'b001101111110101011001110101111000001010000000110100110011010011010001001100110110001111011100001001101010101010011111011110011000010000010010011000111011010110110000111011111100011000101100011010000000100001;
#1 $display("%b", po);
# 1  pi=207'b101111101101010001110101010011000100001011010111100100110110110010010011011111011101010111101001010110100100111100001011011011101000000011100000000010111111101110111010001111111100010000100101010000111100101;
#1 $display("%b", po);
# 1  pi=207'b000110101011110101111100000001010011000000000110001001110000100000010110011010100000110001100100110000101100110001100101011010110001011101001011010100000010110111001001110011111110010110110001010100110011110;
#1 $display("%b", po);
# 1  pi=207'b011111010100111010101001100001101110011010000111010111110110011101111110111101111101111111111111111000111101011010110001101010100110000001011100111111000001001111010110101010001000001011001011111011010000100;
#1 $display("%b", po);
# 1  pi=207'b100010011101010000110011011111000111101010110011001001111110010110000111010101000111000100101101010100001101011111111101101000101100100001001111000001100110100101100111111101000001111010110110110111010111010;
#1 $display("%b", po);
# 1  pi=207'b111100010110001110000110101101100110010001110110110100100110101100011001110000110100011100100101010000011110100010111011101111000110111110101000110110110111011000111111000000001011001001001111110100101001101;
#1 $display("%b", po);
# 1  pi=207'b010100101101001101001011001010111010101001001110001111110001010010111100010010011011000100011000010101011101110110111001011111110100001011000110011100100010010011111110010100000111100001100111001000010000001;
#1 $display("%b", po);
# 1  pi=207'b110111001111100011001010010011010010100010100110111010100001101100101000010100101101110101011000101010110010101111100111100111001110100111101001011011110001001111100001100101000001100011001011100111011110000;
#1 $display("%b", po);
# 1  pi=207'b110001111000111000110000110100010110101011100110111010111010110000111110101010110001100100100100111001111100001001000001000111000110000000110111101000110000100001110000111010000011011010111100011000111101111;
#1 $display("%b", po);
# 1  pi=207'b011110111111110010011001101100101111010001000010111111100101011100100100110000011110110011011100001000011001111111001111101011111000000101000111000010000001100010100110011110111111010010110010000001000111010;
#1 $display("%b", po);
# 1  pi=207'b000010111111010101011001100000000100111010101100010101110110110011011001011111101010100110010111011111101000110001110000111000011000010001100010101110001010111100011011110010111010110100100111110000011000110;
#1 $display("%b", po);
# 1  pi=207'b010111111001000101011101110110100001110011010110110011010011011111010010011000111100011111101010111011011101101011010111000101101011111101100100010101111110100101100101110000100110001110010100011010011101101;
#1 $display("%b", po);
# 1  pi=207'b111110010101110011101111011011000101110110001011001100001000001001000000111000011010010111011011011101100111101101111111011000010100101110000100101101000001010011011011110000100110011010100011000100011000100;
#1 $display("%b", po);
# 1  pi=207'b011100010100001111111100011000111111100110100110010101100000000100001100010100011010010110101001011101001110110101100000011100010001110100010001111001010101010011101000101111110001000001100110001101010011111;
#1 $display("%b", po);
# 1  pi=207'b110111101001010001100110001011101011110011011010111010011010111001010111111110010000111100111111101100011100010101001111000110100110011101011100000110000001100110000100111010011010101011111100111011010001000;
#1 $display("%b", po);
# 1  pi=207'b111100100010001000101000000011111100010111111110110011110011111101001010110001011101001011100010111111100110100100011100101010011000001101010101000110110110011100101001000110110000111110101001011111011110010;
#1 $display("%b", po);
# 1  pi=207'b111101101010011111000101001100100011001110000010110101010111011110001010110100010111110010111010111110111001011111100001111010110001011000010100100001111010000110001100001001001011011011000101001110110011010;
#1 $display("%b", po);
# 1  pi=207'b111011010000111011110110000000100011011110000101001111100101000010100011011011110001011011011000000000111011101011000101111000010100011110011101000110000000001111001000001100000000110111000000011010000001111;
#1 $display("%b", po);
# 1  pi=207'b011110101111110000111100100100110010000000111011010001100011001000011101111101101110100000110001110110111111001001000101000001011100100101110111100000101011110001000000010010011001110110110010111010010001001;
#1 $display("%b", po);
# 1  pi=207'b110000011101001100000010001111111110100110010101001110001110100111100000011000010001101001001110101001010111000100001000101100010000001110111101010101111101011111101010010000001110010000111000101001010111111;
#1 $display("%b", po);
# 1  pi=207'b111000110011110111001110100110011101110111101100001001100010110111010010001110111001100101011000000111101010101000110000010001101010111001010100001100111100011011000011111110000100010101100110000100111010101;
#1 $display("%b", po);
# 1  pi=207'b010010000101000000000101100101101100110101010011111011100101001100111001111010011001110001101010001101010000101001001100001001110000111110110000110011101001011111100011010110110101010111100111011001111110010;
#1 $display("%b", po);
# 1  pi=207'b111010111111100000101010110010110011010101110000101001011010010010100011101010011010011110111110011010101100110111011010110010001000110010100101101000010000110000110011100101101111110100101101110001110000110;
#1 $display("%b", po);
# 1  pi=207'b010101010010011000010001001011000000111100101101011010010010010000111001001110011010110010000111101101100101000001010000111010001100100101110000001011110010100110000101000011101000110011110100011010110100100;
#1 $display("%b", po);
# 1  pi=207'b010101001001000111000011100011110011001000110101110001000110010110010101100001010111100000010000010111111010100111000001000110100110110110101000001010111101001101111011001011010111111100111001010011011101011;
#1 $display("%b", po);
# 1  pi=207'b010000000100110011100001110101011111100100111000000100011111101001010011111101100111110100011110101100111000111111100011101110000111010110111001001111000010000111101011000010110100110100101110001001010010100;
#1 $display("%b", po);
# 1  pi=207'b011110110110000110011101000111000000111111100111001000001001001011111111101110000001110101001010110111111101001010010001001000001101001010111000000100100111110000000001011010000110010000000101010111001010100;
#1 $display("%b", po);
# 1  pi=207'b111100101000011101110101101011101010001110010110101010000100101100010110111110111101001011101011101111001100101001110100101001111110100011110010110110110010100010100110000010010010101100010110011101101001000;
#1 $display("%b", po);
# 1  pi=207'b110001100111101010011110010101011010001000000001100010110100001011111100010010100111010011011011011000000011100111010010000011100011000010110001000001100001010100100100000101100101000110011110100000000110001;
#1 $display("%b", po);
# 1  pi=207'b110000011110100010000000110001110000010110101000111010100101010000011101101010110000100000100001001111000000111000100101101110000000110001100000000111000010011101000100011101001001111000010100111101100110001;
#1 $display("%b", po);
# 1  pi=207'b110100000000100101101100110010111111000111101110110111010110101000001111101100111000010001110101111000011110110100111111000101110011101000111111100011000001000100100011101111100001001111010010000111111100101;
#1 $display("%b", po);
# 1  pi=207'b101001100101011000111101100110001000110101010000000111000110110010111100101011010010010100101110010101010010111010010111011100010111110000111111110100111110100110000100101011111110101001000111011111110110101;
#1 $display("%b", po);
# 1  pi=207'b000011001010101101011101100011111110100100000110000011111100111110100010111000010110010101001011110111111001101111000100011010101011110110001110101101110110010111011010110000111100000011000101111001111111100;
#1 $display("%b", po);
# 1  pi=207'b001110011110001111110000011100001101011000110111110011110100101001100010100000011001010010111100000111110011000000110110010010010101100100111111000110100010100101100010110010110001110110010101001001101010111;
#1 $display("%b", po);
# 1  pi=207'b101110011011010000111101100110111001011001110101001010111111010110110001100010101010010111100101101011010001000110000111111011100100011010001000111110001011101011000110011011000111111100010110100111000011001;
#1 $display("%b", po);
# 1  pi=207'b101000100110011000010101101101101001010110110101001011001101000100111011000011010100101010000001101010101111001101100000100101111011010001100000011101011000000111000001011000010010010010000101001101110111011;
#1 $display("%b", po);
# 1  pi=207'b110111011100011001001010000001110010010011110010011010110110101101000100110100010010111001101000100100010010100101011110100001110111110110010010110101111110011001001001011101010110011010010110000110111011111;
#1 $display("%b", po);
# 1  pi=207'b101110110010111000001100100011010011011010000001001000100111010001111010110000000011000110011010110010011101010101001100111011011111111001110010100000101000011111000110001111000000100100010010111001000100110;
#1 $display("%b", po);
# 1  pi=207'b000011110000001110011011011000010010110111000001000110010001001110110100101011100000110110100110011010111111100001101001111010110001010001100001000110111011100001000010001001001100001000100010110000001011001;
#1 $display("%b", po);
# 1  pi=207'b000010111100010111111010110010111000101011000110001100100001110000101111101001011101010100011001010111010000010111000100100000011001101000111001110100111100100011100010100100110011111001100101001000101111000;
#1 $display("%b", po);
# 1  pi=207'b110111100011011100101110101111111100001011000110101010111000100111000001101011010010011110011010100000010011110111010110010111110001000010010110000100000011010111111101110110110000101001000000101100100110100;
#1 $display("%b", po);
# 1  pi=207'b101010011101110111011000001100101100000100010101111111101000100001110100011000000011110011000011010110000000111100101011001010010111001101101110001111011110110011010000110100111011011111110101010000101011000;
#1 $display("%b", po);
# 1  pi=207'b011000110111101110000110010001010100101011110000001111111010111010111011111111101101000010111101100101010011010011110010010111011011101100110100011001100100011111110101110110001011111000100101010001100000011;
#1 $display("%b", po);
# 1  pi=207'b110001000011101010010010010001100000101001010001101110111101010001000010000101101110111011010010100100100011010001101011110111001101001111100010101011001001010111010111100110000000010001000011001000010010111;
#1 $display("%b", po);
# 1  pi=207'b111000000111011011111001111110110111111010001011101011010101011001110000011111010010110110001110111010011010000000000000100111100011010101011011010100001110010110011101010100011010011000110000001010001000111;
#1 $display("%b", po);
# 1  pi=207'b100000000100110101100001010011001000001111100001111001100111100000100100110011101000010001111111001000011101000111010011011100010101101111110100101010101001010111001101101001000111000110110011010110110110100;
#1 $display("%b", po);
# 1  pi=207'b110000111111000000100011000100011101011110001100000000100011010000110110111001110110111000000011110010101001111111101100000010100111000111101011001001101001010000110010110010000111000000111110111110101010111;
#1 $display("%b", po);
# 1  pi=207'b110001011000110001000101111000010111010011111000000000000100111010011000011010000111111111110010110010000001000111100000010100100011100011100011100111000010100101001010101010111110111101101110010000010101011;
#1 $display("%b", po);
# 1  pi=207'b011001001110110001100111100110011100111000101011010111011110100001100010000100001110011101110010000010111111101000010101111011010101011100100111001011010111001111110101000010111011000110101111000000011101010;
#1 $display("%b", po);
# 1  pi=207'b110001100101111001101101111001010111101100111001101110110101001011000010111110101110100100100100011110111110001001101010000101101001101001111101111010110010111101001000010011000011000010010111011000000101010;
#1 $display("%b", po);
# 1  pi=207'b110010110110100110101000011010000000100100011101100011001001100111100001010010100100010110111011100010101111000100110010010001010000011010000000111000000100100101000001111111001101011101001000111110001001100;
#1 $display("%b", po);
# 1  pi=207'b111100101100000011111001111111000100000000100100100011010010000101101010001111000001110000100110001001111100000101100011100110111011011011001100001010111111000001110101001000111110001101111011011001001101010;
#1 $display("%b", po);
# 1  pi=207'b111101101101011111100001011001100111100100100111010110100010100110001101100001101010001111101111000011010100011001001001110100011111000101101011111110011011001111111111001001100100101110100101100101011001011;
#1 $display("%b", po);
# 1  pi=207'b001011010000001011001000101100101011101010101100000011111101100000100110000100001000011000110011010000101001111100100010010100010010110100001110001001101101101111010000011111111110011100000010110100101110111;
#1 $display("%b", po);
# 1  pi=207'b011100101001101100101010001100011100100110011010110001101001011000001010101110011100010011010011011001100001100111011110001110001110001111010111101010010000101111000111100101001111010101111100100101000001011;
#1 $display("%b", po);
# 1  pi=207'b000100001011111110100101100000011000101010100111101001000110011110011110010110011011000100101110110101111110111000101110101110010111110000111001001011111000111101001010111101100101111110100011101010100111000;
#1 $display("%b", po);
# 1  pi=207'b011010001001011100010100100100011101100011011111110010100000111010000000000001101001111001010001100011000111100100010011110010111011111010100111000110100111010101101011110100110010101101011101111111100100110;
#1 $display("%b", po);
# 1  pi=207'b100110110100011111100000100111010101000110101101101000100001011111100010000011100011010101011001011100010000011010000011100110111001101011000101001110111101101110100011001000001010111100001110000010000011111;
#1 $display("%b", po);
# 1  pi=207'b100001101110101001110111110001010110111110110000010000110100010111001100001000000011110000110000111101111000000011000010100010101001101001000100101011010001001001010111111010001011011111100011010111011100100;
#1 $display("%b", po);
# 1  pi=207'b011000100110100010000001111000101101011100110101110011011010000000111000100001011001100001011010010100100001000100000010011111111011111101111100111001010001110110010101011101001100100100001110110011000011110;
#1 $display("%b", po);
# 1  pi=207'b001110000001111100011000111101111001001001101010011001111011001000001101010010111001000000101011110111111100010011010111001011100110110100100011000001010100010101000010010111111111111100000001110111111110110;
#1 $display("%b", po);
# 1  pi=207'b101000110110011011010001011011101011100111101010110111000101011011100010001001110010001010101111111011010111010000010101111110110001110000110100011010010011101111000011010001111010010001000100011100000000001;
#1 $display("%b", po);
# 1  pi=207'b110011100000101111100001011010010100010110000010110011001100100111011100001000110011110010000110110100110001100100011111001100000101001100111111100001101011100010001100110000110010001000010111110110100011001;
#1 $display("%b", po);
# 1  pi=207'b100000111011111101011101011111011111111101001110101001111101101010110100111101100001011000111000001110101000100011111101101010101000001100100000000111011110011011110110110110110100100000110111111110010000010;
#1 $display("%b", po);
# 1  pi=207'b110110101101010000101101101011110111101001100000010001110110001110111001110110001110111011010001011110110000011000001000100101101110100110011100111100110110111101011000000110101001000011101100110011110100101;
#1 $display("%b", po);
# 1  pi=207'b101110011111011111000011000011101001100101100001001101011010010110010111101011100011110100001110110011100000111111010000010101010000101110111110011000100010100011100000110111111011010010101000100000110100100;
#1 $display("%b", po);
# 1  pi=207'b000010000000001001110010001111101001110010010011000100010111110000011101111010010100001001100010101011010001000111100100011100100011101000000010110111111110000101111001000001010011111100000011101010100110101;
#1 $display("%b", po);
# 1  pi=207'b010010000010011011000111110101101001110110110111101100001000100100110100110101001011100111000111111111011001010010111000100001010110111011001101100001100111101010000110001100110010110011000101001010011010011;
#1 $display("%b", po);
# 1  pi=207'b100010111010010110010100000000011010001001111011011000010001101000111011111100101011000111000000011001111100111111111011010000111000101100010111101111111000011101110000110001000010100000010100110111000011010;
#1 $display("%b", po);
# 1  pi=207'b111010011001101000000010001100100100101010110001100011000100111111111001011111110010110100110100001100110011110101100000010100110101111100000001100011011100010000111010101100010011111110011101100011101011111;
#1 $display("%b", po);
# 1  pi=207'b111011101001100111010110110011100111100110010010101010000011100000010101010101010111001000011010100110110000101011100001010111111111000110100000001111101101010000111000000101111101110100101000110101011001100;
#1 $display("%b", po);
# 1  pi=207'b010011010010100100101011111111010011111100011000001011111101101011100100000001010101001101101100110111001101110000000101000000100001110111011111110001001011110110011011100001100100111010100110001101100000101;
#1 $display("%b", po);
# 1  pi=207'b100011010111100110111110100010010001011111001001001001100101001001011100001110100011000111001111001001110110100100110110001011110110000010010111101110000110100011011010111000111000111000101001101001000010011;
#1 $display("%b", po);
# 1  pi=207'b100111101000000010000010111100000001011100011100001010001111110111100100011011011001101001000010010110001000110010101011010001100011100011001001100110000100000000110001011000110011101010101111010110100100111;
#1 $display("%b", po);
# 1  pi=207'b110110111010101011100001111101101100100110001000001011001100101010000111111111010010100110000111100110010011101101110001010110001111101100001101110010101110000100000010000000011111000000001001010110011111010;
#1 $display("%b", po);
# 1  pi=207'b101000101001010001111001011010111100100011100001110111111000010010110111001111100001011011100011000101001111100110100001111011111111100100100011100011101011111000110100011010101001011011100100001000011111101;
#1 $display("%b", po);
# 1  pi=207'b110110000001110111111010000001011100101110000000011111100101001011011110100011010010110111001000101010110110000110110010111101011111011010000101001011010111101111100010001011010000101001010101111111101000101;
#1 $display("%b", po);
# 1  pi=207'b100100100010100110000011101011110010110011110101100110100000100000110111010110101011010110010001011000111101000011100101111111011010010101100100111010001101100111001000100101110100110010001001010101111011101;
#1 $display("%b", po);
# 1  pi=207'b001110101011100111111011011100010111110000000110001010111101101111100111000011010001010101111101111000000101000111000001001011011001000111000110001010010001011100011000100000010110000011011111011110010010000;
#1 $display("%b", po);
# 1  pi=207'b000001110011111111001101111010100101101100110001001110111011011101110001110100011100001100101111111001101110001111001111011101011000000001100001100101001101011101010100010110011010001111110001100000001101000;
#1 $display("%b", po);
# 1  pi=207'b011001111001001011001111000001000001111011101101100101011111011001100011110100000010111011110110001101111000011000001111000100000000100100100111100000111011110110011010100001001101100110110111101010011010010;
#1 $display("%b", po);
# 1  pi=207'b011110110010101110000011111111010110010011100011010101110000001001001111010101010000001100100100010011011011101100101101110010100001010111001011100000010001100000101001001000101010000011011101001111011011011;
#1 $display("%b", po);
# 1  pi=207'b111110010000011011101110011011010011011000001111001010110110111110111110011010000001101100101011110001101100010111000010000111110100001111111000000100001000000010011101101000010101111011011100111010011101001;
#1 $display("%b", po);
# 1  pi=207'b001011011010110100100010001100101111110000101110100001010011001010010010001001110001000101001101110101111001000010111110110100100001100100000101001000110111001000111010111010110101110110000101011000000000111;
#1 $display("%b", po);
# 1  pi=207'b100111010000110001011110010011011000100000000010111111111000111011111100111100010100110100111011001111111111001011101100100110111110010000010100001101010010000010110111000001000111011100111100001110001001010;
#1 $display("%b", po);
# 1  pi=207'b100101011100010000011101101101111111000100001101110100100000111101111100000111100010101011110010110110010001100100111101110001000101000011101010100111000000000011001001100111101010110100000001010001110000100;
#1 $display("%b", po);
# 1  pi=207'b010000011001011001100111100111101110001000101001100001101010101011001110101001101101011011010101001000001110010010100100100101001111100110111101101000000001001011010001011001111111110100000111011111000101111;
#1 $display("%b", po);
# 1  pi=207'b110110001111000010001010001111000011011001101010011100001000111101001100111101000110011101110100001001100011110100111011010101010011010110001110101011001101001000010000111110001110001111001011111111111010101;
#1 $display("%b", po);
# 1  pi=207'b000110011001001110111110001100100111010111001111001101001001111001001000100010010111000110010000101001101111000001000001110010000111110011101101100101001111011101111011101010001100110011111001110100010111101;
#1 $display("%b", po);
# 1  pi=207'b011010000111110010000010100011011100010110011111110101111011111001011001010100101011100111010010111111110110000010101100111010010001000110011100011100010110011101000011111100011011100010011101011111011101011;
#1 $display("%b", po);
# 1  pi=207'b001010011001101100110010111101000001100000010010011100101111100110100100010000110010010001010000101010111011101111001100011000001000111000000001010110011010100000101011011111011101110001001101000001100101010;
#1 $display("%b", po);
# 1  pi=207'b011011101010010001000000100001010010011111100001010000011001000000111011110110011110011100011001110110011001001010111101011001011110001010111000101100110110000010011110110000100111100110000100010010110010011;
#1 $display("%b", po);
# 1  pi=207'b011101100100110101000010010001011010101010011000100110011110010001100111110011010101011010010100101010000101010011110111001000100111110000101110010010011110000100101101011000010100100001011111110101110100011;
#1 $display("%b", po);
# 1  pi=207'b110011011110011010000001101001110110111010000001100001111000111111110000110111000110100101101010011001001011100000111010000110100101111100010000011110100110101000010010011101001011111111111110001110010010100;
#1 $display("%b", po);
# 1  pi=207'b011010011101001101001000110001010001001011111000011101010101110010101010010011010111110011001110001111001000000100110011110001010100100101001011000110111011010011001000011010100101110001110011010011000011100;
#1 $display("%b", po);
# 1  pi=207'b010101001100101000100000001100000001000111010011010111111010010010111110101010000001100110110010000011111000100110101011101101011111001000010100110110101010110111101001110111111110011001011001010010111000101;
#1 $display("%b", po);
# 1  pi=207'b000000100100000011100110000001100010010001010000101101001000100011101010110010110000100001100101101001101010111010111011010011110110010010101010111111100101001101001011001101111010100100011010011000000000100;
#1 $display("%b", po);
# 1  pi=207'b101010101011100111101000101000101000100100011001110011001001001000110101100011101010100011110111110001101001010111111101101010111010111100011001000111010000101011100110110010110101010111111001001000101110111;
#1 $display("%b", po);
# 1  pi=207'b001100111001111011100110010010010110011011101111000110100110111111000110101100000111111010100110010110001101000100000100011100111010101110001100110001001101111101100101010011010011001100101011000010110011100;
#1 $display("%b", po);
# 1  pi=207'b000000111001100011110101110100110000010011011101010100011011000011011001110111000000110011110011010101000010001101011101111000010000001111001100111001110101111110011000100101111111110101000010100001110111101;
#1 $display("%b", po);
# 1  pi=207'b000110110101110111001100010001000111001010101111001011100110111101000110001101001010011111000011111101000100110111101000100011110110000100011011001111101100000111101100110111010100000111111011010100100101111;
#1 $display("%b", po);
# 1  pi=207'b010100100001000101101001101010111111010000011111000011100100011010011101101010111010101100100001000100000001100110110010001110001000110010100111010000111011111101100101000110110011110000000010110100000011011;
#1 $display("%b", po);
# 1  pi=207'b110011010101110110010010110101011010001011100000101010111000110110101010111101100111000101101010001110001011111010111010101100000001111111101001000010011010011100011111001101011101101001111111111111010001100;
#1 $display("%b", po);
# 1  pi=207'b010111110111101011101111010001100101100010110100111100000111111000100001101000010010110100010101111101001010111111001100001100100000011110111100000111010000101110000010000111011000100001111000011000101100111;
#1 $display("%b", po);
# 1  pi=207'b010010001111101110111011100000000101100110111001010001010101110000111101011101001011101101101100001010111000110011011000011010010001110010111011110010011001001101010001101000111010010010111111111101000010010;
#1 $display("%b", po);
# 1  pi=207'b001010010011110100011001111110101100011111110011001110010000100110100101111101000100100010000111011011100101101111001011011100011100110101001100101001110111010010110001101001101110111110110001111011111111111;
#1 $display("%b", po);
# 1  pi=207'b110100101111101011000100010100100001010111111010001100010000010100001111101111010001000000110001000010001111101001010101010011010101110001010001001110001101011010000000011110010100100011101111111100111101111;
#1 $display("%b", po);
# 1  pi=207'b111100000010101011110101110101100010101011001100011000101111010010001100100101011000110010101110001010100100111010110001111000001101110011111111110100101100100000011010111111010011110111111100101001001101100;
#1 $display("%b", po);
# 1  pi=207'b100011111101111100010101111111111000101101111100101111000100101000111000011001110100010000101101101101000101110110101011000101110111000010100010000011111111000010101111001010110100110000101101011001001010010;
#1 $display("%b", po);
# 1  pi=207'b111100000010010000000100010011011001110100110100001101001011110100111010111111101111000100011101100101010110100000010100110110001101000101001110001101001101000110010000110111100010100110010001001000101000100;
#1 $display("%b", po);
# 1  pi=207'b000100001110010010111101000000101110000001111101111011101101011110011001011110101001010000001101111101100010010101001101011100110010101001111000010101011010101000110001101110000101101010111101110011000000001;
#1 $display("%b", po);
# 1  pi=207'b110000111101011010111010001101110100001011000011010001010111100100100000101100001011001101001111011110001000001011101010110001101111011010011100111010000100111110111110101111000100101111001110000000010011111;
#1 $display("%b", po);
# 1  pi=207'b011100010010001101111110110100010101111111100111111101111000000000100111100001110011011111000010101000011001000010100011001110000001010101011010101100111111111011101111001110000001011000010011001110100010011;
#1 $display("%b", po);
# 1  pi=207'b100110001011100010011100000001001001001011000111110000010111000000101100000111001101001111100011000000100111110001111010010111101110010110010001010110001101101010101011000101100010000001110000111100110010100;
#1 $display("%b", po);
# 1  pi=207'b110100001010111111001100011001001111001111000010110111101011011010001010100100110001100111100111101100010011101110001001101111011001111011100000011000100100010110111000001001111010001110000000000011100111011;
#1 $display("%b", po);
# 1  pi=207'b011001000111100100110001100111001011100001010100010000011111010100111111001100111010011010111110010001010010010011010010010001100100101011111100100011101101111000111000011001011001000001101011110010001111111;
#1 $display("%b", po);
# 1  pi=207'b010111101010000100010010100000000101101000001101001110110011001100100011000001000101111111000000111001001100111101101010100011000010010001101110000111010011101001100011001010111101110100010011100100100011110;
#1 $display("%b", po);
# 1  pi=207'b110010110000000001011000110101001101000111000111100101111010111101010000011000100111100001110110010110011010100101100011001110010000000001111001010011000011101000010110001010000111110101010011100000011111110;
#1 $display("%b", po);
# 1  pi=207'b010101011010011110001010000101000110101001010111010101110100000111011101001110011001110000011010111010111011001110111000110011011110010111111111000001110111001101010000001010111010000001100100110101111000110;
#1 $display("%b", po);
# 1  pi=207'b000010000100000011110101110001101100100010111100101001010100001000101101101010011100010011100000011100110010001010110000100110100111110011000111010011110111101100100000000110001101110000100000001000000000000;
#1 $display("%b", po);
# 1  pi=207'b110010111111001111110110010110000101100001101111110111010010101001010001110000110100001000110010111100101001101011001011111001010001011000011111010101111001001110011100000010000011100010100101111001111011100;
#1 $display("%b", po);
# 1  pi=207'b111100001011000000010100110011110010101010100111110111110000100011100010110011010101101100100100100110000100111010010100111001000100011101111101110010101011110001001100101100111110010110000001101011000001000;
#1 $display("%b", po);
# 1  pi=207'b100010110001101001101000111010010110000101101100011110100000011111011000111000111111101011100001101010000110110010110000100110111110011111111011111000100001111110110000011010110001110011111010000110000101010;
#1 $display("%b", po);
# 1  pi=207'b010100110011111001101011010011010000110000000000000011100010100000100011100010000011111111110110010110011010000110111111111111001101101011001010100001111010011000010010101101000110000111001001010110000001010;
#1 $display("%b", po);
# 1  pi=207'b100000000011111101001110010110000010110101111011111001001111010001001110110001001001111110101010101100101011011110100100010011001001111011011100010001101011010000010100101110011110010111100101011111001101100;
#1 $display("%b", po);
# 1  pi=207'b110100011010000101010000100010111000110100000000110010111111110001110010011010101001000001100001111000101011110101000110001000111110001010100010011111001000011011011110001100110001100000000010000000100111100;
#1 $display("%b", po);
# 1  pi=207'b100011100011000011100110000101110011111001010001101110001110011010000001101110100100011110110110001100101100011110000100110100101100010000100010010000100111001010001101010010000001000100000011001010110011110;
#1 $display("%b", po);
# 1  pi=207'b011110011010100111110011011011000110011110101110011010011010000111101011111100010011001001001101110111010111011111111101010111001001010110111010000111111100101110000110101001011110010001101110010010011111100;
#1 $display("%b", po);
# 1  pi=207'b111100111000001011110101000101010011110101101000110101010111011011100111110000010011101110110110100010000110010111010001111001011110100110110011001111101000001100011101011011010101001010010100100011100011101;
#1 $display("%b", po);
# 1  pi=207'b011101110100110011011011000101011111000111110000011000010000100101001101100010110100011011100111100111101100000001100011001010100011110110010011011100110011100101010011011111111100100100110011010101100000101;
#1 $display("%b", po);
# 1  pi=207'b001111011011100111111111111001101101111010111111000101100101100011100110101010110100100111111101000111001101000000110010100111011011101111010111100111111101001001100001110010000111100000011001111110011100110;
#1 $display("%b", po);
# 1  pi=207'b011000110110110011100011010011001011110010001001011000001110011100011000100000101101101100111000010100000011101100010001101000000001001000010001000100111110101001011000010110110001111100000000010110101100111;
#1 $display("%b", po);
# 1  pi=207'b001011001001110000111010010001010110101000110010001001011110011010011101010101100111111110000010011110110100101110011010111111110110100101001000011100101010111110000011110011110111011011010010011000110100000;
#1 $display("%b", po);
# 1  pi=207'b011001011110001010101100101000000101101101011100001100100010111010101001011011000010000110101011111001000101101101000001100100010100011101001100110001100110001001101110001110101111110000101010010100110110000;
#1 $display("%b", po);
# 1  pi=207'b011101000100100000010100110100001111110110001000100100000000000010100010100010100001010101000100011011110001101111001100011110010100001100011011001001000111000011101101111111111011010111011110100111011100110;
#1 $display("%b", po);
# 1  pi=207'b010011100111011100101000011011001101100000100010110011000010110000011111111001110111101101101000011100001110101100100110011100100111111000101010011000001111000100001011010001101000010111110110010101011101011;
#1 $display("%b", po);
# 1  pi=207'b100010101001001000101001110001100011001101000010000100001100100000111111000010111001101110010101100000011000011111100001101100010110011110111010000000001111011000100000001101011001011010101101111001011110000;
#1 $display("%b", po);
# 1  pi=207'b100100110100111111101001010010001011100110111111110101000101101001110110000111101110011010100010011110010100100011110101100110111100110010010011111000110111000000011011010011011111110110100001011001001111011;
#1 $display("%b", po);
# 1  pi=207'b101001101111101100100001010111100100101000110000000100110011010111000110101001100110111010100110110000111011010110000101100111010000010000011101010010011111001000010111110011000001110001111001110001111000000;
#1 $display("%b", po);
# 1  pi=207'b100111000001110010110100111111100101111000001111110010111100010011110000001001001000110000011000110110010101111110001110001101111000111110011101011101011001011000111001110111010010100110111110100101011011101;
#1 $display("%b", po);
# 1  pi=207'b010100011001011000011000101101001011010010111011010101011011111001001000101001111111101011000101110010111100110101010011001101110101001010111111100110011010111010111110010111100011101100101010100000000010100;
#1 $display("%b", po);
# 1  pi=207'b011111101111010111010100111011100101001000000000100110100101111110100011000111001000010010011100000011010011011100110101010101010010101010000010010111011100011100110010010110100101110111010011001100001011111;
#1 $display("%b", po);
# 1  pi=207'b011010101101111110100001110011001001010001000001111110110010000111100101101110100110111100101011000001111010100010110011011100010001111010100111100100010001111011100000111101101110111000100100100111010100000;
#1 $display("%b", po);
# 1  pi=207'b111010101110101111101001000011100111111010101110101111011111010111110100010101011010100101010011110111111011110001000111011101001110100111001000011111000100100111100011000000010101001000010110001110000100100;
#1 $display("%b", po);
# 1  pi=207'b101101100000010000010001110110101001101100010111101010101101101010000110001000100100110011000000011100111011010111111111101010111000101001010101111110111101101011100000011011101011001011101000100010110111001;
#1 $display("%b", po);
# 1  pi=207'b010011100100101110110001101110001000010111010000010010011101100111010011000000110001100111011110110101101010000010011011110110001000010010000100001110110010011000111010110001010101011100100000101000100010110;
#1 $display("%b", po);
# 1  pi=207'b011001110101101011111011111110101011010101010111000001000011010100101010101101001101010001001100111011010100110100100000001010101000001001010010101000100101000111100011001001101100000100000011100110111010111;
#1 $display("%b", po);
# 1  pi=207'b000001011110001011010110001101111011101110110010010000001010111101001111000110001111101100000110000111100011000110010101010011101000111001010000100110101100011100100000011111110001110000101110000001000101011;
#1 $display("%b", po);
# 1  pi=207'b000000111100011011111101111001011110000111000010011000011001011101001100111000111110001000001000101001001100010010010100000100100101100111011111111001001101011011011110100100110011011010000010101101010100111;
#1 $display("%b", po);
# 1  pi=207'b000011001001001011110010100110100000111001110010101010110101000011100101101001101110010101001001111110001100001011100000110111011111010000010011111101001011010011001010101011110111110001000001110010001011111;
#1 $display("%b", po);
# 1  pi=207'b010010001001001001010001001001101011011110001110001110011101001010001000101111010011011010011000001100010111100101101000000010010000100111110000010010111001111011101110100011111011010111010011101101001110010;
#1 $display("%b", po);
# 1  pi=207'b101101001101011101100011101000100100010101000000101010011011100001111010010000000111111111001100110101110011101111010111110111101110111100100100010001100010001101011001010010111011000101000001101111111100111;
#1 $display("%b", po);
# 1  pi=207'b001110011111101011001101010111011100110100011100011001110010100011100001101110011110000110001010101011011011101110011111011001110000111110000000100000100011010011101110010011101010001101000010010011000101101;
#1 $display("%b", po);
# 1  pi=207'b100011010111100110101111000101011000010100001000011100000010001101000001111100101101100100011101011001011011110110100010000010110111110101101011010100010000001111111111010001001101100010101111011000100011110;
#1 $display("%b", po);
# 1  pi=207'b001001001010000110101011100001111010111000111101101100001000000000001100111110101111011010010010110111101110000010110110000110010010110110100010011010010010010110111100011011101011101001111110001000011001111;
#1 $display("%b", po);
# 1  pi=207'b110001001110010100011101111010011110011000011000010011011110001010110001001010010100111010101011011011101111000010010010001100100101111100011100110101101011100001101010011111000111111101001000101101001000000;
#1 $display("%b", po);
# 1  pi=207'b000111110100100001000110110110001100111101001010101100010001010100110110110000110110111010100010110001001110101111111010001110100011000100011101011110111111101011010110011110110101110100100000011110111100011;
#1 $display("%b", po);
# 1  pi=207'b101101001011100001011001000101011001001101110000010111111001100101101101010011000101101010000110110010001101101110011101001001000001110001111010101001010100000011101111101111111100000010010011110000111000111;
#1 $display("%b", po);
# 1  pi=207'b101101001101110101101100010010100000011111010101010101010111001000000111010011010110110101101101101011100001111110011001010010001011011100001000101011011101000000100111100110011100000011000111001010111110010;
#1 $display("%b", po);
# 1  pi=207'b001010101111100110001111111010010100100100110111111000101010100011011100010010111010110100111100000111110110101001011001101111111110000011100010101111010011011100110101110001110011011100010010110111110001011;
#1 $display("%b", po);
# 1  pi=207'b110111000101101000101101010111000100111010010101100101101100001011101101100011010111110010000111110100110000101101110110111000101101000000101110011111111001110100010000010001001011010111101111110000111001001;
#1 $display("%b", po);
# 1  pi=207'b101110100100110111001110100010011000000011000000100100010100000011111101000100111110010110011111101110100100010000110100100100000011011010000100111001000000110111000001100000010000100000010101110111000111101;
#1 $display("%b", po);
# 1  pi=207'b101010010101001001000000101100101110110010111110101011001101001011111111110001111111110101011101110111100101001001100011111011100111001100010000001001100110100101000010000101100100110001001110100101111101001;
#1 $display("%b", po);
# 1  pi=207'b001101100100011111011110001001011111000110110111100101011001001100011011110000100001001111011010111110101110010110101100111011110010000111011011101001110001110000110000110001001010111101011011011010000000111;
#1 $display("%b", po);
# 1  pi=207'b100111010010010000101100010101111001101111110011111011001101101000010111000010010110000110101101100001100011010010101101111011110010000000010000010111101111011100101111011110000110111101001010110010100100101;
#1 $display("%b", po);
# 1  pi=207'b100100001010000000101111000011011000100001110111011011110100000101101011000110110100110110100101001101011001100111111000001111101111000011010010100101001110100100011011111010101001000101101100011000011001011;
#1 $display("%b", po);
# 1  pi=207'b101101101111111111110111001000011110001110101111010000111011000000110001001001010100100010110101100110001110111110001010010001100100111100110000011110000010111010110101000001110101000001010000000001101000000;
#1 $display("%b", po);
# 1  pi=207'b011110000011010000101111010010001110110011011111111010011100000010000111101111001000011101011010010111110101010001000100010100111011100010110100001110010101000010110110011110100101100100111111111001011110110;
#1 $display("%b", po);
# 1  pi=207'b111110100001100110001110101110110001100111101110001111111111110011110101010010000000101100101001001011111110111101101001111101101100111100100000110011011110000100001000001011110000000111100100110100110100001;
#1 $display("%b", po);
# 1  pi=207'b110101010000101010010110100110110101101101110110001010010000000101101111011010011011010101111011010101010010000100100111110000001110001010110011001011111111101000011001111010100110010111111001011000000111100;
#1 $display("%b", po);
# 1  pi=207'b011001100000110001011110010100101001100010100111101100000011101101101010111001101000011011110101001101111110010101001111001000011101110010010010111101110100101000111101111001100001110011010001011100011100110;
#1 $display("%b", po);
# 1  pi=207'b010100111101000111100010111011000100000111101100000010100001110000010100011110010110100011110101110010101011000000001000000011001101000001000000011010000010011110110101110100101100010011100001000100001011001;
#1 $display("%b", po);
# 1  pi=207'b001101000011101011011101111111011010000101011100010101111000001000011010000000001011000001100110110000101110001101101000001110010110010010011011110111001111110100000100001000101100110101000011010000110101001;
#1 $display("%b", po);
# 1  pi=207'b001111111110100000100010101111011000011100111111010110011000111100111001100111001111000001111000110111010001111001001010010010111000100010001111101000010001110100111111101011000110111000111011111011001110011;
#1 $display("%b", po);
# 1  pi=207'b000101000101001001000111010000000011110000101011110000000111001011011101000010101000010001001000111010100001100110100001111011011100101111111000011110101101101111101010110001010010101010000000010000010010010;
#1 $display("%b", po);
# 1  pi=207'b100001000100101001101000110010010110111000111000011010100011001000010111111000010011000101001000001011111110100110100101001011001010101110101101111110110001110000101011110001111000101100110111101010100100100;
#1 $display("%b", po);
# 1  pi=207'b011110011110010101100100101101111000111111000000010010110001111111110000100100101101100100110111011100010111110010011101111101011000100000010111111010110011100101110100000111111010100101101010000001110101011;
#1 $display("%b", po);
# 1  pi=207'b010010100111000111000100101001001110101101000000011010101011000010001110011111100101011010101110100111101000101001000010010101110011111010001110101010111101110111111111011010100111111110000001110001101011000;
#1 $display("%b", po);
# 1  pi=207'b101101111110110100011111111111001101101011001001000101100010100001001101111100010010110001000010101010010011010001111101000111010100010111001010001010110110000001110001100100011001101100111110101010010111100;
#1 $display("%b", po);
# 1  pi=207'b111101100011100001010110110001110100111010010010000001101100011010000001101011100001100010000111111100100101100001110010011101111010010000111101010010100010001011010111101001111010011011110001101100110100001;
#1 $display("%b", po);
# 1  pi=207'b000111001010001010111010100100110000000001000001000110110100010001010110011111110011001001111101001110111011110011000111110000011011100111101001110000000011011100111011100001011001100111110001101010001110011;
#1 $display("%b", po);
# 1  pi=207'b000101011110101111101001001101011011010110010011000100101101010111001111100001100001100110000101110101011101110100110111011111001001110010011011010111010110011110011110101110101001100110001010011111100111111;
#1 $display("%b", po);
# 1  pi=207'b101001110010101000011011001000000111100110110011100010011000110100111010101010000101010101111101111111001111001001010010111111110010101100100110100100100110011101011001100011101000111110111011010010000111011;
#1 $display("%b", po);
# 1  pi=207'b111101100100000001101100000011011101110001111111110111001100111010101100011011101010111001111010101101111001111011110110100101100101111111111001100100111011110100000000011110111111111100011100010010000000110;
#1 $display("%b", po);
# 1  pi=207'b101011110001000110011000001011111111010111100011101101010000000100111110011011001001001111000100100010101100010111100100111010101110010000111110000000001011011000000000100111110001001010011110001000110011110;
#1 $display("%b", po);
# 1  pi=207'b000101011011110110010000100111001111011110011011010110101111110111001100111010001101010011101111111101101000001101111010011010000010010011011110011000010001100000011110011100000001000010010100110001011010001;
#1 $display("%b", po);
# 1  pi=207'b010110011011110111011001101001100010111111111110101111111000011101010011001111011100111011110111110101010010110111100001010100111111100110001100011011101011101001100100001100111110001011011101000010010111100;
#1 $display("%b", po);
# 1  pi=207'b010001001100100101100001010111100011110111111110010011101110100011101101110100110101011000000011011111111001010000001101010101110100010100001011110100110001010000101011101001101001001100000111110101111110010;
#1 $display("%b", po);
# 1  pi=207'b011100110100100000111110110010000011101001100001101100000001010101111010111100000000010000011011001000010000001001110101111101001000110010111000101000100011011000001011111110010000011001011110000011001011000;
#1 $display("%b", po);
# 1  pi=207'b110100101011000111110011100000101000101010101010001001011001010110100110110110011010011010011100011000110100010110001000011011010000101011100111110001111110000100100010001101100010111110011100100101010011010;
#1 $display("%b", po);
# 1  pi=207'b010001111101011110101111101110010000100111110110101010011000001011011011101010001010000100101101100010000100011000001011011111100011111100001110100111111101101101010110110001111000110101111100101110001101110;
#1 $display("%b", po);
# 1  pi=207'b010110111001100100011100110000111101001110000011010000010101001101010110001010011010000010110000110110011010000011000110010111000000101111000001111111101001100001011110110000000101101010010111001011001100010;
#1 $display("%b", po);
# 1  pi=207'b101010101111000011011000010110011000011001001111010111001010011111011011001110100000100110011101011011000100011011110011000011110000101100101000100101001100101010010101101011111101101111010001001101110100001;
#1 $display("%b", po);
# 1  pi=207'b111010010111110010101001101110000000000011010101110111110111001001101011011111001000001110011010111100000110110110100100110011101110110000100101000100100011110001011100111110001001100010000100001111000000010;
#1 $display("%b", po);
# 1  pi=207'b011111001110110000000001110100001000100101000100110110001111001110111110000001010110101001011111110000000111100000011110111001010100101100100111010010011010000010011101110001110011101110101000100111110011101;
#1 $display("%b", po);
# 1  pi=207'b000001100100100111010100000001111001011110100011100111011110010111110110110101001110100000111000101000111101110100101010100011011100110110101011110011000101010111011111000110010101011111110001100111111011111;
#1 $display("%b", po);
# 1  pi=207'b110101000010000111100111100111001001001101101010011100010000110100000011111011010010000100111011001001001100111001001010110101101010111111101100101101110111000001101001111100110000011111010111010110111010010;
#1 $display("%b", po);
# 1  pi=207'b110010101100111001111100110101110110011110011111110101010110101011001100000110100001111111001011011100010101100001011000001110101110111010001101111010011110101011010011010011000011100011101001000100111101111;
#1 $display("%b", po);
# 1  pi=207'b011010011001010111110001000000110101011001010100101111100100000001011100111001011011101100000111100011110111100100011100101011001100011100001010100111100010110001100011100010010011001100101011000010110010101;
#1 $display("%b", po);
# 1  pi=207'b001001000001001000101110110101101000010110001011111001101001011101000010101001011100010010010111011111010100100000011000100100110010101001011000111011000101100010000010001100010101110010011100010100111000110;
#1 $display("%b", po);
# 1  pi=207'b010010110001100001011111110111101100001000010101010011101111000101010100010001000001101101010000110001000101011000110110101110111011101011100010110110101001010011100010110111010111100000100001000111110011111;
#1 $display("%b", po);
# 1  pi=207'b011110100101101011011110111100100101110011100100000001100111100111101111110111100101001000110011101011110010011000111000011101000111001110001111010101000100100110010000111010011011000000111101010111001000010;
#1 $display("%b", po);
# 1  pi=207'b001110110011100110011110001110011000100000000010011000101001000101111101011100101101001001011001010111010010100111100100101011111011010001101000110101111111111101101110001010101111000011111100110010011110110;
#1 $display("%b", po);
# 1  pi=207'b010010100101101010010010010011000001110001011011100110100001011011100011101010001111111111111000110011000000000111010011101100010001011011001110011001111101101010000100110011100010111111111111110010110110110;
#1 $display("%b", po);
# 1  pi=207'b101100111000100000111101001001110001110101111100000000100011001001000110111010111101111011100100010011011011001101010010110011000010110010111010000001011001010110001001001010011110100001100010000000001110010;
#1 $display("%b", po);
# 1  pi=207'b000011011110001001111100010101110100000100001111001001000000001110100011101110000110011010011100000011011111100111001000110010011010010110100010000000110011110100011110101001110010111110110000101111011010001;
#1 $display("%b", po);
# 1  pi=207'b010000101011011011100100111111101010100111101111101111110001111000011110100110110101000001110011010110110001011011011000011001100110111101110101110101101011101000010100010010101010011001110100101111011100011;
#1 $display("%b", po);
# 1  pi=207'b000011100110000000010100111111001100100100100110110111101101001011001010110001010010011011110100111001111000100010011111000000100101110010110010110001100101111000101111001101100100111101101100000100011101110;
#1 $display("%b", po);
# 1  pi=207'b011110000001011111010010010101100000110100001001111011111100100101101100100100100010111000000000010011111101000110011100111000100110101001011011011111110100001110100100101001111110000110111000100110000111101;
#1 $display("%b", po);
# 1  pi=207'b001100010111000001111010101010000010010100101111101110101110010111110100011100100011011000110001111110110110111111100110000000000010111111110001111111001010110111100001001110110100101111000000000110000011111;
#1 $display("%b", po);
# 1  pi=207'b111000111010110001000000111001000000000011001000101110101100110010011100000000000010100110100111011010001101110111001110101100111011111100100100000001000111001111111010111111110000111000011101001110110001001;
#1 $display("%b", po);
# 1  pi=207'b100111110001011100110100001101111110010110111000000000010011010000001010100100100000101001011110110111111011011110001011100110010101111001111110011110000110001000010100000000001110110100010011010011101100010;
#1 $display("%b", po);
# 1  pi=207'b001100001000100001111011110101010100111001000111101110100001111111001100000010110111001011100010010111001001100101110101111110111011011011100000110001001100100011000001000100111011111011110001010111100010101;
#1 $display("%b", po);
# 1  pi=207'b111110001110000000001111110001011101000101000111011110001100000101110001101100001001000001001011001111111100111101001000110110110001011101011000101100010110100001110011100110001011001110100111101101100010100;
#1 $display("%b", po);
# 1  pi=207'b011101111011000111111101111000011010001100100011001101010110111100110101110111110011000100000100000001000000100111101110000000011101100101111100010010101000000101011101100111110110000001001110100000000101000;
#1 $display("%b", po);
# 1  pi=207'b111111011011010110100101000000100111000110001011000001011000000011010111111110111111000000011000000011011101000011000111110110011011111011100110100010100101010111010010110101111111001111000100000000101110111;
#1 $display("%b", po);
# 1  pi=207'b000000000001010001111101001101001110010110001111100111011011001000101101110110011001100011110101011011001001010100101000001101010100100101000100010001100100110110010001110010001101011100011101001001011001010;
#1 $display("%b", po);
# 1  pi=207'b001001010110110011100011111010011000000010111010101000001110010010111011000001100001010010001010111110110000010101000010011000100110011010001011100110010111001101110101010101110011110011000110110010011000000;
#1 $display("%b", po);
# 1  pi=207'b111101111101000010100100011110010111101100011111100100000101010110001000110010101001010001010111001011010011101100111001010101110111011111010100000100010001110000101011001000000011001000001001101110111000010;
#1 $display("%b", po);
# 1  pi=207'b101111101101101111011111001110100110101111110101011100110011100000100100110011111000011110000000101111001100100111100110010001101110101101001111110111110010110011010001101000011011000001010110101000010000000;
#1 $display("%b", po);
# 1  pi=207'b001001010010010100001001010100101101011001001000110011100110100000010011110001110011100101101100000010110011011001100001010001110110000100111100010110000110011011110001110110100100010011111000010000011110101;
#1 $display("%b", po);
# 1  pi=207'b101101110001011001000011000001100110000000110101100110101010010001000010000011101010111010001000011001101110101000001001100000101111000100101000011101111010001110000010010111111111011110101010010011000010110;
#1 $display("%b", po);
# 1  pi=207'b010001011011011000110100011000001111000101100010001100101101101111011001110100101101010111010110010011110001110000011001111100111111000010110010001100100100111011111000010010111011001000000010101110111001000;
#1 $display("%b", po);
# 1  pi=207'b011101011000001111000010001100110000001010110001101011011000110110010100110010001101110000110100110001011011011001100101111100001001010000111001101001111011000101111001011000111110110000000101111100000100100;
#1 $display("%b", po);
# 1  pi=207'b000111010000100100001001000111100000011011000000000110001000000101111011101111001010100011101000100001001000001101110111001111111111100111111100101010001110110100010010101011011011011001000011100111111001011;
#1 $display("%b", po);
# 1  pi=207'b011011011111001000101000011111010000011011000110011111010111101100010010011101000010110111000101100001010011110000010010000011110011100101000101101100100100110000100101111001010110001110010011101101010001011;
#1 $display("%b", po);
# 1  pi=207'b111000111011000100101010011110111000110111011011001111001111000101010010001100110010000100010101010111111110001000110101110111111111100110010111010000110000000010101000111111101011100010111100100001010000101;
#1 $display("%b", po);
# 1  pi=207'b101110000110101000110011100011001100101101000101110011001001000010101100100010110110101010001000000101101110111001010110101000001110110000100100100111100000110101110111000000001100101111110110010010001010101;
#1 $display("%b", po);
# 1  pi=207'b111101000111000000110001100110101010001101101111010011111011100010011110000111110101000110000110101110011100010010111000010100010001011001011101111011111100001010111011011110111010110100110011111011011011100;
#1 $display("%b", po);
# 1  pi=207'b101110010110111111111001001010111111010110101111010110111010011100110111011010111110000010110100001011110000000100101001011100010010101111100100111001101100001101100111010110010101001110010101101001101000000;
#1 $display("%b", po);
# 1  pi=207'b100011110100011010110101100111111001101110011111111001011101001111110100110000011010010000101000110010100111000011000101111111111011011101101010101111110001101100111011010100011000010101000011100100010000100;
#1 $display("%b", po);
# 1  pi=207'b001010111000000000110101001110100001001100001110111010101001010111000110010010001101101111000010101011000101111011011010011111011100110101000100100001011000100100101001111101100110011000011111010101000100000;
#1 $display("%b", po);
# 1  pi=207'b000001110001001100101111100110001001000010100101100000111000101101111101110100100011101000100001001100011110111111000110110101010011001101000000101101100011101000101110010001011100000111111011011010011011011;
#1 $display("%b", po);
# 1  pi=207'b000011011001001000111010011010000111000001100101011000111110110110000010011110101110001011110001100000111111001111101001001111000110101001111100010001011101100100001011111111001100100111011001001111111000100;
#1 $display("%b", po);
# 1  pi=207'b000010000001001000100001010001001100000001100001110001100010111100101000101011100001000111101010110111111001111100111110100110101000110011101111101111000111111001100110010001000010001110100111011101100100011;
#1 $display("%b", po);
# 1  pi=207'b101101011101101011010010111010000010110110111101110011100111001110110110101000011111100111000010110000010010101111010001011111101001100001111010111001000100110100100001101110010101110111000111010111001000111;
#1 $display("%b", po);
# 1  pi=207'b101011110110111010111100011000101110101001001000011011101101100000111010101011011101001100000111010010101000100111101101101011111001101000000010110000011010010110011001101010010110100011100000100101101111010;
#1 $display("%b", po);
# 1  pi=207'b010001000100101101101110011110001100111110001011010110010110011011110010001000101101000111100111110011110111110111110101000011101010000111001100001100001110011100110101101110110101010001001110100101010110111;
#1 $display("%b", po);
# 1  pi=207'b100101010000011000111000000101111110010010111110111001010010000111111101011000011010111101100101011100100000111101010000000011111100110100111011010000100000010111010001001011110001011010000011101100111011010;
#1 $display("%b", po);
# 1  pi=207'b000000011000001000001001101011111000110101000010000101100110010000001100100000001101111011101111110100111010100100000110000111001100000100100101110100101100000101110101000111101100010000111101111101100110010;
#1 $display("%b", po);
# 1  pi=207'b111110010111001010101001001001101100011100100010110000101001001110011100000000101010010011011001011001000110100111111000010011010011101010100101101010011100000011110000001010010111011010011110101011011110100;
#1 $display("%b", po);
# 1  pi=207'b111001100010110110000100011000110010011100111010111101101011011100011010000101110100110000110011000010001110001110001010010111011001010000111101011100010100111100100100100101011011011101010011100011000010110;
#1 $display("%b", po);
# 1  pi=207'b101111101010001001101011010110110011100011100101111000011000111011000110011000111000110110011110001011000100101111110010110111010101110111000001100001010011001001011001000010100011000001011100110101101011111;
#1 $display("%b", po);
# 1  pi=207'b011000111111111111001100010000000001011111011101101111001101011110110000101011101101101011100000001010101100010110010111000011001001010111010000000100111101100110111010000110010010110000101000110001111011001;
#1 $display("%b", po);
# 1  pi=207'b001110000101001111010110000110011111111001011111100000000100000011000011111110010110001011000010010110101000011011111110010001110100010000101111100010010110010101000100011000011011110100011001100101110011100;
#1 $display("%b", po);
# 1  pi=207'b000001111110101101110100010010000111111110001101010000100000100100111101111101111111111011010011110101000010001110011100011010001010111110000110001111000010011001111000100110010011101110100100001100000000010;
#1 $display("%b", po);
# 1  pi=207'b101101100000111110111011001100101101110101000011111011101000001101010010010010111000010001110000010111111110101001001111000101001001000001110111011110001000010001110000110110100111001011110111001011010101001;
#1 $display("%b", po);
# 1  pi=207'b001010011011011001000000001101000000001100010110110101001100000110000010100000010111000110110000110101010101111111001111000010111110101011001001000001100111011000100000000110000101111110001011111100010111010;
#1 $display("%b", po);
# 1  pi=207'b000100010111010001011110000010011110100111010001011111011000001000100001111010010011011011000011101001011010111001001001011001011010010011110001100110111101011101010101011011110000000001011010101010110101100;
#1 $display("%b", po);
# 1  pi=207'b001011000100100011100100001111010111001001001010000100010100011101101001011101110011100011100001110111011000011011001101010000101001010011100011010010000111000111111010110101001011110100111101000100011110000;
#1 $display("%b", po);
# 1  pi=207'b110110111111110101011001111010001000110101011100001011010101101011011100111000100100000110111110100101100000110011110010000011011100111110100101101011110111010110000110101011000000101000110010000101110001100;
#1 $display("%b", po);
# 1  pi=207'b101110011001110110111111111011001110010100011000111101101101001110101110001101000011100000001001011101110100110011111000011101101000100110111100000010111110111110000111001110001001101011000010001011110110010;
#1 $display("%b", po);
# 1  pi=207'b110001111010110101010011100001000010001001001101001111101110000110010000111100110100000101010001101111110000110000101110100100010101001010000110000100001000000110011010011100010000010010101111010010011010100;
#1 $display("%b", po);
# 1  pi=207'b010011010011101110001100001011110001001000110110110010001111010101010011001101000001100100100010010011010101111010011101100000101000011010110100100001101010100101000110110001101011101011100011001101111110000;
#1 $display("%b", po);
# 1  pi=207'b111011000100000001101111000110001011101001101101110101010100001001111011111101101101110001011101110011000001100101000000110011001010001001101001100111001010110000001010010001001001111010010110010110110010000;
#1 $display("%b", po);
# 1  pi=207'b100100111001010010100111100111100010110010101000010111100101010001111000001111011010001000000010111111101010110101001101010111011001000100000001100011101111000100000001011001000100111110010110101111000100101;
#1 $display("%b", po);
# 1  pi=207'b110110011110010000111011010011100111100100000000000110110110011110000000001101111111000010101000010000100011110001010100001101101000010000110010001010001001010011101101011010011011011100011011100101100110010;
#1 $display("%b", po);
# 1  pi=207'b100101101001100011111110011010001110111001010101000101001011000101110111110011011101101100000000010001011101010100011010110100001110000110000101011011001001110000111010011000011111100000011101111110101100111;
#1 $display("%b", po);
# 1  pi=207'b010011000111010001000010111001001111100001000011011000000110010101111011011000010111100101001001010001001000110000111011100110011011110101100100011100101010111110101111111001100010001000000010000001000000001;
#1 $display("%b", po);
# 1  pi=207'b001110100100010010001110000111100010110111111100011000100011101010101100100101010000101000101010011010101110010110110010100010101001101101110101001110100000101100011011011101001011000101011110011001010010011;
#1 $display("%b", po);
# 1  pi=207'b101010101011000001111101000111000101001011101000010000101111111101100101000011111001110100001011011100101101000010101011011111000011000101111000011111011001111010101100110101110101101101011100011111100000100;
#1 $display("%b", po);
# 1  pi=207'b101100010101001001110011101001111010000010000111000100110010110100101100101101100111111100101100011010111011101000100100110011001001011000100110110111101011000000011111001010100001000100110101000001101100011;
#1 $display("%b", po);
# 1  pi=207'b000100011111100100100110111100110110010110001111011010001110110101100101000111000010110011110100110110000111111000110000000101000110011000111000111101011011100110111101100000000011110110111011100010000100101;
#1 $display("%b", po);
# 1  pi=207'b001111101100111000001110011000111110110101010010100110100100111101001001110010110100110011101110011101011110011010011111001010000000100000100010001111100011111000110011110011000101001010010011110010011011101;
#1 $display("%b", po);
# 1  pi=207'b110110110000101101100100111111101111101110011011100111000000011001011000111100110010000000100100100111011111110011000010101110011101001110101001111010010110001100110011010111101101001100010000110111110001000;
#1 $display("%b", po);
# 1  pi=207'b110101010011010101001100001111100011110110101011010110001000010010100111110111011101111100110010101010000110100000111110111111100100111101011111000010000001011101110101110110001100111100110101101010001100110;
#1 $display("%b", po);
# 1  pi=207'b011100010001011111110111010101111101110110110010011011011111110100011000000100110110011001010000000101000100011001000111110111010111101001101000010011001100011001100010100011110001001100001111101110011111000;
#1 $display("%b", po);
# 1  pi=207'b110110111110001101010010101010011010010010101101111100011101010001010000110101011011011000110111000110110010001001000111110100111010010000111000110110011010111000011100001101011010110011111111101010001011101;
#1 $display("%b", po);
# 1  pi=207'b000111111111001000011110010110010101101000101111010001000000111101101111011000100011100000011011100101000111111111001100111111111100010001101111000101111111100011110110000111111000101100001011110111000110100;
#1 $display("%b", po);
# 1  pi=207'b100000111111100101100101011110011010010100110100101011100101100011111100011001110011110110100010000111111111001111011100100111000100001010110010010001001011000101000100001101111010001101111111100110011000110;
#1 $display("%b", po);
# 1  pi=207'b101101000000111100010011101101011100101101101101101010001101001010001011011010001110110101101110001100111001111111000101000000010001010110011110111100001011001101111100101001110000100000110100011111011101010;
#1 $display("%b", po);
# 1  pi=207'b111001001011010110111110101111010000010100001100101101000111110010101011111011110010010101000100101100000100111101000011100010111110010000101110111110111001111010100111111011111000101001100010110111111000010;
#1 $display("%b", po);
# 1  pi=207'b011010010111101110001001010110010111111100111100100111101110100101000010110000011011111010100100100100110011100011110001010001111000011010101110010101101110110100000100010010100001110110001111110001011010010;
#1 $display("%b", po);
# 1  pi=207'b100000001100110101111110010111001000111010100010100000000110000000010011001011011110111001100000100011011100100000100100100001000001000110111000100000010000001011100110001101111011100101000000011100100110001;
#1 $display("%b", po);
# 1  pi=207'b110101110010101101110100011110010010001101101001011011000101101011111011110100011111110111000101010101111011010011000101011011100010011110001100001001010111001101010101001111011010011000111111100100110000010;
#1 $display("%b", po);
# 1  pi=207'b011000100100111001011111001011111010110010110100011011010111110011010110101110001100011110100101011100001010011110001000000110111111100100101000000010101110001100001010011100011100010110001110111000100111010;
#1 $display("%b", po);
# 1  pi=207'b101000011001011110000000011000110001101010000100111111110010111100100101111010101000110100100111000001001100100000110000000100011111111010001101010001000101110001010111110000101001000110011100111101010101010;
#1 $display("%b", po);
# 1  pi=207'b010011111010001011000000011001001011101111110100101100110000100001101101001010010100100001111100100000100110101001110100101010101101000110110100111010100110111001010010100010111000110110001100010110000110111;
#1 $display("%b", po);
# 1  pi=207'b110101101000001010100011111011101011100000100101000111100100100011110110010001111100001111110011010101100010101010110111001101010011001110111010010111000111010011100101001001000100101111100101110000101000100;
#1 $display("%b", po);
# 1  pi=207'b001010111010001111010111110010100000011110100110001111000111110000001100001110001111010010101000010110100001111111110011011111010101000010100110000011110010001011000110101001001000111010011001010010101110100;
#1 $display("%b", po);
# 1  pi=207'b100000010001010010100001111000010000011000010100101110100000111101001111011010110100101001100101100000000000010111111010110100100001110010010111111110110000001110010010110101000100000001011111100001101001100;
#1 $display("%b", po);
# 1  pi=207'b010001101101010101000110010111111100011100000011011001111100101011010001011010101111100100011111110111011000011110110110100011011011111010101001001111000101110000001111100011011100111111110001000011111101101;
#1 $display("%b", po);
# 1  pi=207'b100111110110111101110111010100100011001011101101001100111101100010010010001000111100000010100011010101101101100001000010100101100000100100101000100110011100111000011111101111100010000110011001000101100010011;
#1 $display("%b", po);
# 1  pi=207'b000100010011000000001100010111111010101110111111101101110111101011000100011101111101001000011011011101010110000101010000101111100010111100110010111011111111111111011011111000110110001110110111000010100110001;
#1 $display("%b", po);
# 1  pi=207'b000010000110001000111101001100000101111110100011011110011010101000111001111001001011110001011010100011111100100000110010111101101001111001010000001101101100111001111010001111100110101010100001000000110011000;
#1 $display("%b", po);
# 1  pi=207'b100110110010100011001110010011001010100101000101110101001100100010110111110001110100100111001100111111110010000011110100000101000110000010001111100011001011110111101001010011000010001010110001011100111111101;
#1 $display("%b", po);
# 1  pi=207'b101111001100001000000110111000011011111110000000001011010111001001110111001011000101011010100111101001111111000000000000011000011000111000100111110100011000001011001010011001001111000000110101001101111111011;
#1 $display("%b", po);
# 1  pi=207'b000010000000010011111001101011000000010011111101001011100001010010000100100001110110000110100101011110001111100001101110111011111001111111011001010001111110000110011100011100110111110110100010010111000011010;
#1 $display("%b", po);
# 1  pi=207'b001111010011111101001010000110111110001000010101011000101001100010001000001001010000111111010000110001011010100111100110100100011000011101001001100101111101100110110011011010101111101111000111110111110011000;
#1 $display("%b", po);
# 1  pi=207'b101000011111010000101000001001110001011111101010101000001100001010011101110010011001100110101111101010111110111001101110001110100111011111100111011010111111100011101011001101111010010111100001011111110110001;
#1 $display("%b", po);
# 1  pi=207'b110011111110000000110000100111011110010001110010010110111110000101001110010001110011111111011100010001000110111111100101100010111111111100111000111000111000111100010011010001111111110000001100011100001000110;
#1 $display("%b", po);
# 1  pi=207'b001000110000101111011100110101010001001110111101100000000110110100011101001011011001010000101011000010011001101010110001010111011100011100110111100000011001001111110111111101000011110000000111011011110000101;
#1 $display("%b", po);
# 1  pi=207'b101111001000110000011101010111001011111000001101010101110101101011001111111100101101101111110001110000100100110111011110101101100001000001111111111001010100001110011000010100010110101001011111001010011100011;
#1 $display("%b", po);
# 1  pi=207'b001010000011011011011111010101111101101011011111000011100001110111010000010101101011110001100101001101101101101010101101011001000100110000100110110011100100000101001001111001000101001000111010011010010011000;
#1 $display("%b", po);
# 1  pi=207'b010011011010111110010110100011000110100011011001101011010000000000101100100001001010000111000001011110110001101101011001010010010001100101011010101101011001110011111010010100000111100011011110010000011011110;
#1 $display("%b", po);
# 1  pi=207'b101111100101010100011010010100111100010110001111110110010111011001010100001000101110100111001100011011110001001100111010101111100101001010001101001010111110000000100001111000011100000111011101001101001010110;
#1 $display("%b", po);
# 1  pi=207'b110110101000001111111001100100000010001001000010111000101001011100110101001010011011010111011001110110101000011101110010000001100010101000010111100110111000010110100100111011100011111101110010010111011111110;
#1 $display("%b", po);
# 1  pi=207'b000011111101000010111101110100111011111100000001000011100110010000100110010001101011110000000110010010110010100101011011000011110110010111011001001100000011001010111010110111111111100000001000101111101101010;
#1 $display("%b", po);
# 1  pi=207'b010110110100010100011111011001111101111011001100000110001010001100111000011010000000010101100110011001011010100010110011000010001111010001000111111011110110011001000010100001010011111001000111110110011100111;
#1 $display("%b", po);
# 1  pi=207'b110001111011101110000000100111010111111110001101001101110110111111010110000000010100011000001110110101010011110000111011110011001010111110110110011010101011000101001000011101100111101110011001001111101111100;
#1 $display("%b", po);
# 1  pi=207'b011110111111011110000111000001001000110010111010101001101110100000100011101000100011110000011011001101001110001110000110001111011100110000001100110010110111000110011100101100100101101111011011001101010101110;
#1 $display("%b", po);
# 1  pi=207'b101101101100011110001100110100101010101001101110001001010111110001001000101101110110101111111111110011011100101100101110100000100010111110111101100100101011000100000000110111001110100100010010011111110010110;
#1 $display("%b", po);
# 1  pi=207'b011001010101001001111011100111001010011001101000001011011111111100100101101010111010001010011101100110111101010100100010000011010110100101001111100100010010010010001111011000110011111100100000101001001111101;
#1 $display("%b", po);
# 1  pi=207'b000100100000100111111101010001011010001000111000100010001000011101111001111111110011111000001000101001110010001011011011010010001111110111011111100101000000000001111101000100011101101100011000100111100111001;
#1 $display("%b", po);
# 1  pi=207'b000100001001000011111101010000001001011100010110010010110100001010100101000010000001011010101101001010011001010001001001110000000001011101000110000001010110001000110011001100100110101100110000100010001010100;
#1 $display("%b", po);
# 1  pi=207'b110000011001011100011111101010101011001101101111100101000000000000000100010100010111000010110001010111110011100010001000110100101100001100110101100100100010011100011010011110011000010011110110001100010011110;
#1 $display("%b", po);
# 1  pi=207'b011011001000001100000010101000000000110101000011110101001000000001111110010111111101010011000001001001110101011000011110011101001100111001001101000000100000001001010001001100001110010000000101000101010000000;
#1 $display("%b", po);
# 1  pi=207'b111001001111110000110100001011110011110101011111101010011001101100100011011110011110001010100011010010011100111000010110100000010111001100001001011000110100001101010111111100001000100010011111011011111011100;
#1 $display("%b", po);
# 1  pi=207'b000101001101010101001011001100101101110110101110001111010110111101001000110110101010000001110110100101010001100011111011011011101101100101001101001000101010000100010100011110110110110111001111110010110011110;
#1 $display("%b", po);
# 1  pi=207'b100110001100001111101010010100011101100010011111111111000110000110101111110010010011001110110001010100011110001000101110011101100010100100001100011010100101010111010111111111001100111111011100101000101011101;
#1 $display("%b", po);
# 1  pi=207'b101101100011110011001111100011100010111011000010111101011010010100101010011111001100001010011011010000011100111100101111100010101000111001100010010111000100111100011000001100001101011000101100011000001001110;
#1 $display("%b", po);
# 1  pi=207'b100101111001010110001010001001000111001010011000110011101000111111100000111110000100010000011011101001100110111110001100111010010111111010111110000111111110101100011000100000010101011100001111010100110110100;
#1 $display("%b", po);
# 1  pi=207'b100111101101000000110110101111001100110011100011001110010001110111011110101000101111001011100001110000111011011000001111010111001101101010010010000100100000010010100000110100111110110101110011000010011101101;
#1 $display("%b", po);
# 1  pi=207'b010110110000101110011001011000111110100010111101010000111001100110101000110111010001101000100010010001000111010000101011111100001111000011100100110101110001110011011010110011010110000101100010000101000111100;
#1 $display("%b", po);
# 1  pi=207'b110110110010010000101001101010010101110101110100111010000010001010001100000111101011110110100110100100111000011011010001110100111100001110000101101001100111110101111000100101000001010000001111100010010101110;
#1 $display("%b", po);
# 1  pi=207'b010010000110000111000010001111101110110001101011001100001000111110001011011101100011001011101011011000001000101110011101111101001111000110111010100110011011000000100111011110000110110110001100100100011001000;
#1 $display("%b", po);
# 1  pi=207'b101000100101101101011110101010011111001010001011111001110101100000100100011010010111100000110000011100010101100100111000010111001100111100110100000101001111100010010000001100011100110000001011011000111000000;
#1 $display("%b", po);
# 1  pi=207'b011110010101011000100010100010000011010011010001111011100100010000100010110001111110001100101010010100111101101110011000000010101011100010111010101101100110011011111111101001011110011111100010000110100111100;
#1 $display("%b", po);
# 1  pi=207'b011111101011100101010111010111100111011001011000111001000101000011000111110000010010111011100100101111101010111111000010111001001010110110100101110011101100110001001110100011111010011110111000011110011111001;
#1 $display("%b", po);
# 1  pi=207'b011100010000010111001001011010100110011110011001001101011111000101100011010111100010010110110011010010010100010100111100101011010100001010011001000111010100011000111001101010001110101000000111100000110010101;
#1 $display("%b", po);
# 1  pi=207'b011110010110110001001110000000011011010110010101010100100100010110100111110101001010010001100101101110100000101010100000111111011101011001000110110010010010000110010001010110011001110001101101101010100010001;
#1 $display("%b", po);
# 1  pi=207'b000110110101001011000011011011000100111101110100000111100110111010110111010100001000100101110101010011010001011111010001100010111100000101000000111101000100110100111110101101110110000011110001001010001001101;
#1 $display("%b", po);
# 1  pi=207'b111111110010101111011011100101010111011111111001100011010100011000111110110000001010001000101001110110110000110011111100111010101001001111011000010101001001011100110101110001001101000100110101001011001101010;
#1 $display("%b", po);
# 1  pi=207'b101000101001001010010010011100100111001010001001100111101011011100111100110100101100100001111000100010111001011101011010101000000000111110111010010110111010011010100001101110000100101001111000011101001000000;
#1 $display("%b", po);
# 1  pi=207'b010101101001000101010011011101100111100001000110110000001110101001101000110010101111101001110001000101110111010010010110100010000011101000110101000010100010111011100000011001011110111111000011101001001101111;
#1 $display("%b", po);
# 1  pi=207'b111011000110010110111110000110100011011001101000100101111101111000110000101001011010111111110110000101000011010111100111100011010110011101001011001111110101100001101101010100101000101001111110100011101110111;
#1 $display("%b", po);
# 1  pi=207'b101100100001000110010101001000101110001010001010000111011010111101101000000001011111111001101101010101001000110011101101110110011010000100101101111101101100100110011110101000110010011000001111100111001000000;
#1 $display("%b", po);
# 1  pi=207'b101101110101001010000101111011110010101001100010110101000011000111100001111110000111001000110100101101001011111111000011011001101111000010110011110110111000111100010011001111111001001000101110111100110110010;
#1 $display("%b", po);
# 1  pi=207'b111111001001101011110111011011111011011000111101111011000110100010101000100010010111001001010011011000001110011011111000000011010010011100110110111101011011011110111011100111101010100011110000101000001011000;
#1 $display("%b", po);
# 1  pi=207'b001110000001010001100110001111011000011110100110101011000101010111001000001000110100000001110111100011110010001101100011110101111000001101100100000101111100010010100000010000011111101111110001110011101011000;
#1 $display("%b", po);
# 1  pi=207'b000001111110111101100001101111001000100111001100101011110101000010100001011111101001000000000011100000010110010011010110010111110111100010001101001000010010001010000110101101100101010000101010000101001111111;
#1 $display("%b", po);
# 1  pi=207'b100100011100000000100001001000010100000110001111100000101100101101110101000100000101111000110100010101000110011111110110001111111010000100010110010001110011000100110010000110011111110001010101001011101010111;
#1 $display("%b", po);
# 1  pi=207'b101010001011000001110110110111100000001101000101000100001010011011011010010100001101011100100000000001111100110100100100000111110011111000100111101100001001101101100001111101011100011110010010110111100000011;
#1 $display("%b", po);
# 1  pi=207'b101100010011110011110001101010111010110010010100010000001110110100111011000110000010100110100000011001110111000110110000010010101001010100010101001111111010000010010101111010001110001010011111101001110101101;
#1 $display("%b", po);
# 1  pi=207'b100100101011000011011000100001111011100110110001000111011010001001100111011001110011000110111111011111000001001101110100000000000001010101101111001100011010000111100100101100101110101110001010010101010110011;
#1 $display("%b", po);
# 1  pi=207'b011001111100011101111000011000000100001011100111111100010000101111101100011111000101111101000001001110010110101100011100001110110010001100010001101111011100000000001110110110101000001011101011010100001011111;
#1 $display("%b", po);
# 1  pi=207'b111111010000110111010011010000111001101000001011000011001111111100101100110001010101101110111111001001011110111010001011010110111000110111001010010011000011111000001101111010110111111001100101101000100110000;
#1 $display("%b", po);
# 1  pi=207'b010101111111010101011100001111111000111100001011100010001011110010000000000000100110100011100010010000010100000100111000000101011100100110100100101010110101011101101111000000001011000010010000100011111011110;
#1 $display("%b", po);
# 1  pi=207'b010000111101101111000011101111001010010011100101010010101101001000111111010111111000101011011100000101001011000011110110010111110001100000000000100000110101000011111100000011000000111000111001110000111000000;
#1 $display("%b", po);
# 1  pi=207'b001010101111000000100101000011011111001000110111111000010000111110100010110110011100010101100001101110001110000000101000110010111001100011100101001100001100101101001011100100110011001101010010000010100010000;
#1 $display("%b", po);
# 1  pi=207'b111000101010111001110111001011001100100110000100110111011001001111000110011000100010110110110111110100100101011000100111000010000111011100011001101110101100110010000001111111100001000101010010101001110101100;
#1 $display("%b", po);
# 1  pi=207'b010001010111110101001110110101000001011100010000101111111101001001011011001011110001100110100100000100001011010101100111000001000011110010011011000011101100101100010001000111100100110110010111000011010100111;
#1 $display("%b", po);
# 1  pi=207'b001011010111100011010100101100000001110111010110101000011001000001001110011011010010110100110001010101110100100000100011001010100101001000010111001000011001101100101011101001110001010101111101011011000000000;
#1 $display("%b", po);
# 1  pi=207'b110110001000101110001101111100100010101000001001000000100110101011001101111011101010111101110010110100100000111000110110010111110111010010000000011100010011010010110110010110001100110010011101101000000011101;
#1 $display("%b", po);
# 1  pi=207'b011010101101111011000011001100010011010100011001011010101101001011001101010110001111100101010001101010010100001100101000000101000000101001000001100100010001111110111100101111101101010111011101001111100111111;
#1 $display("%b", po);
# 1  pi=207'b111010010101011001100010011011111011010111011001111011010110111101110001101110000011111101001101110010100011000011101011000110000000011100101001001011011100100000111101101010000010001011011001010111110011111;
#1 $display("%b", po);
# 1  pi=207'b111011100110100010010001100011011111010011100000110110000000011100011001111011001001010000110000011010010100011001010101111101110110000000011100010000110101000001011110101010010000110010110010111110000101101;
#1 $display("%b", po);
# 1  pi=207'b111010110001000011000001110111100011100110111001111011101110101001100111100010110100000000110100101100000011000000110000101100000101100100011001011111001010010001011010101110010001100010110000101011111111101;
#1 $display("%b", po);
# 1  pi=207'b000000110010000101001100011100001100110011110001101100100000001011111110100010010000011101000001010010001101001011110101010111001000010001011010110011101110101110110010000101110011111000101001111101000011110;
#1 $display("%b", po);
# 1  pi=207'b010000000101101100000111000110001111000110011111001000110101011100111111011100011111110000011111011000111110111010111100010111000011011110011000110010110111001101001110101100101101101001001000100001100110101;
#1 $display("%b", po);
# 1  pi=207'b110100011100101010101111110001011010010101100001010000101101010000001010101111010101101111010001011110110000100010000100111101110010101111010100001101110010100110101001110011111001111110100111101000000111011;
#1 $display("%b", po);
# 1  pi=207'b101101111101101100011000110001110000010111010000101100101010010010011001010001111101100001101011011101110001011111001000100110101010010010100011001101011110110100111110100111010110100000000101011111010101110;
#1 $display("%b", po);
# 1  pi=207'b100000011110000011101011000010011000100010001110010111100111100111101111100100000110101010010100000101010110000101100011010111111100011110110010101100110101101111111010000001000001010000100100111001001011001;
#1 $display("%b", po);
# 1  pi=207'b101110101000011111010101010011011011000011010011011000011001110010111101000100001100101110110010111011110101101010100101110101100100010101010100110110100110110111100110001010111001010010110010100011101000111;
#1 $display("%b", po);
# 1  pi=207'b101110111000101010010101101010100110100001100100100100100100011111111100101101011100011110010101000001100110100010101001000010011100010001111111110100010101010111110001110001110010100000011101100110110011111;
#1 $display("%b", po);
# 1  pi=207'b100100000010010101001010001010011110110001101111111001000111000000111110001110001000101010000001101011110010111101010011001011110000100001100101110011000100101000010110101110010001011101101110111000111100100;
#1 $display("%b", po);
# 1  pi=207'b100101011100011000101000010100100100010001101101010110101011111010011100000101001110110011011001111010001100110110011111010101111111010001110111001100111100110001111100011111100100010011101001110010000111000;
#1 $display("%b", po);
# 1  pi=207'b100100101100101101110111011110101101101010111101010101001100110101010000010101000000111100010010101101001000010001001110101011100110010100111001100101101100010101111101111111001011110001110111011010000010010;
#1 $display("%b", po);
# 1  pi=207'b010010000111101010010111010011000011011010111000010000000011001101010110111001101111111000110010111111000111100110101000000110101111001100100010010100110111111100000010000001001100011001010001011001011100110;
#1 $display("%b", po);
# 1  pi=207'b010110100110110001001110010011101110101100110000000011101110111011011000101011011000110010011000110011010011110001011000101110010111111001111001010001100101001100010011011001000101101001001111011111101100110;
#1 $display("%b", po);
# 1  pi=207'b010100011011011010011101110011111011010001101100011100010101011001001000000010100111101101010110110011110101000001111001100101101100101011011111110101001101111011100001110001101110101001010011111000011011101;
#1 $display("%b", po);
# 1  pi=207'b101010111010001000110110011111011000101011100100111010101101101111101011001010001010110001011000000101010100010010000001000100100011000100110111101100111100101100110011010000111000100100000100011001100010000;
#1 $display("%b", po);
# 1  pi=207'b101110110100110111001101100011111111011011111001100011000000111011001111000011101010100111111011110000100101111000100110110110110010100101010010001100011001010111101010100100000010000001100001010110000110101;
#1 $display("%b", po);
# 1  pi=207'b000110000101110111100100111101111110010011110011110010010101110110111001110011111101101100101011011010011001100100011101110101010011100001101101001111001011110110110010010111001011101101001011001011101110111;
#1 $display("%b", po);
# 1  pi=207'b000110100110101010010001000010100001100000000110101111010111001101100010110101010110001011111100010010000011111000110010101000000011011000110100001011001011011001001010101100111101011110001110110100110011011;
#1 $display("%b", po);
# 1  pi=207'b000011101001101011101110001111001001111010001010110010010101011000011001011101110001111000111000001000111111100111001010011110000111010100011001100011010110000100001000111101100001101100011111100000101000101;
#1 $display("%b", po);
# 1  pi=207'b110000101101100000010000001001100010000010110010001100000100010111101110111011000110001011000101011010110101110011110011101011110101100100010011101001110011000111111011000010101101101001011001100010011111110;
#1 $display("%b", po);
# 1  pi=207'b111110000000001100101110101011001100011110000001101100010100110111000011111100100110101000111110010011011110101101100000010101000100100101000100001001111111001111101100111000001101101010110001101100001001101;
#1 $display("%b", po);
# 1  pi=207'b011000011101100011101100110111110111110001000000100001010100111010100110110011101111001110100100100111111111000100110100010000111100011011101011110100100010001010100010010100011100101100111110101111101110001;
#1 $display("%b", po);
# 1  pi=207'b100010010011111001110011101000111100010101111000010000001010001111101011000000010101111001000001000111011110110111000100000010111101100010011111011010001000110011111111000000010111111111100101010101111111101;
#1 $display("%b", po);
# 1  pi=207'b100010001110101001110110100111010110011111001011000000110100101000000100110100011101001111110100100011010101100010111011000100101001010111110011011001101000011101100011101001010011011001001010110000100100011;
#1 $display("%b", po);
# 1  pi=207'b011111000101001000001001010101111010010100101001001011111001100011010010110111010110000000111001100110111000111100010011110001000100011111000101001010011001101010010001010100000111101101110001011000001001101;
#1 $display("%b", po);
# 1  pi=207'b111111000010010100011111011101100110100101000000000100111111100100111100110101100010010100101000101000110110101100000010100100100100011011011110111110011100011100000010101111111000000100000111000110111010001;
#1 $display("%b", po);
# 1  pi=207'b101000111010111000100001011001111000001110011111010001001011110010111011010011000000111010110100100110000100000010000011011011110001110011000101000011111100101011111000000000100111101010101011100000111110011;
#1 $display("%b", po);
# 1  pi=207'b000000111000011001001101111100111111000110011011011101111001110000110010101011100001000010101001010001011000000001000001110010010100000101101011101100001101011001001010111110001010110010001001001001000100010;
#1 $display("%b", po);
# 1  pi=207'b110000001111010111100110111000010001001000011110111101110010011100000101110100011100111100001010000110011111000110010111101010110000101101010001111010100001110010011011111000111100100000100111001001101100111;
#1 $display("%b", po);
# 1  pi=207'b010101011010101010110001101000111011010100000011100111010111000100111110110100101001100000111010110000111000110101000111001001110110010101011001110000110111110000011001011100101111001010011001100100100001010;
#1 $display("%b", po);
# 1  pi=207'b000010101100101110101110101000111000011000101011010001110010101101000011100110100111001000110110010001010011011110111101110010001000100010001110100110011001100110100111000111011011110111101110101111100000100;
#1 $display("%b", po);
# 1  pi=207'b001010000101111101010100001111000001100101110010010100101000111001100001000111111000111110001001010100110010001101110111010010100000100000100100010110011111100101111100011011110010011111011000100101101100101;
#1 $display("%b", po);
# 1  pi=207'b000010001101100000100101000111000011100011101010101111000101011111111111101101011000110111011101010010110101011100010111101010001101001100010100111111000101001111011110101110011100101110010000001010000011000;
#1 $display("%b", po);
# 1  pi=207'b111101001111011011101111010101000001101011011001101001011111001000000110001111110010000110101000111100101001011100100000110110110011010111110011000110011010001111101011110010100001100111100111010100111110010;
#1 $display("%b", po);
# 1  pi=207'b011010110001110001100101011110000000000100100000001110101100110010101101011010111010000101010100100010010101100111100001010101001110010100010011000011111101100011010011010011000110011000000001110111001010011;
#1 $display("%b", po);
# 1  pi=207'b100101101000010110111101100010101001111011011001111001001100101000111101011110111000010110101010010010110110100010000100010000111010000011000101100000000001101011000001000111000000110001001111010110110100011;
#1 $display("%b", po);
# 1  pi=207'b010011100101010101000101110100100011111001110110110001110000011010000101001100110011101101110101000001111100010010000110000110010010001110010010101110110010110010000111100110100101110011010010000101011000011;
#1 $display("%b", po);
# 1  pi=207'b101111101101110000110011110001101011011010010111011011101011111010111110101010011101001111010110001111000100010011100110111000101011101010001111001101101010111011001100111001011011111101011101100111010111011;
#1 $display("%b", po);
# 1  pi=207'b000001110101101010110110111100100011000111110011011011001111010100001100111011101111110111101001000001000000101011001111100100110000100000101100110110000101100010001110111011101100000100010100010100011010111;
#1 $display("%b", po);
# 1  pi=207'b000100101010010010010011010110111001010001101111001000000011111100010101000010100001101000111110100101011011010101000111011000010000110101001011111010011010100000000011111010110110011011111111000100111000110;
#1 $display("%b", po);
# 1  pi=207'b101111001011110111000101111101101010110100010000110010000001011101100110101000010101101100110111001001011001000100001011011010000111001101011001010010010001101111110110110111101110011111111001100001010110100;
#1 $display("%b", po);
# 1  pi=207'b110100111111111100011110100000011001011101010100010000001101111100110110000101100011010100011111000111110111001001101100000101000010001101111110000001101000110011111011011010000001001101010110100001011111110;
#1 $display("%b", po);
# 1  pi=207'b111101001100010111011000110010100100011101101000010110011001101001000110001100110000100000001110001000111100110011001011100011011000110000010000001110001000111100100101110100101011111111011000010011011001010;
#1 $display("%b", po);
# 1  pi=207'b100101000010101011111111010111011010000111010000011111101101001000000000011110011101111111110100100111001100100101011000110111101000011010010010110101010010110000000101000011010101100110001110001001100011110;
#1 $display("%b", po);
# 1  pi=207'b111110011011001000000111010101011101101111001000000100000101101011111110011010100001000111101001000101000110000011101110111011111011110100111111110000000010100111010110110110110000011011100100000111110111100;
#1 $display("%b", po);
# 1  pi=207'b001100111101110000101000001000001101111101100111010001001100000001000110000101110000001101001010011110100100000001011100001010111100011001101011011111111111001000101101111010100001010000100101110010101010001;
#1 $display("%b", po);
# 1  pi=207'b111110110010101001000011010100011101001101100111110010011000100101011100101100001011110101101001011001010100110011001010001101110111011000110000010110001010100010111100000000001100010001100110011000010000011;
#1 $display("%b", po);
# 1  pi=207'b111010110000011100110001010111010011100010011011111000001101001101000100100001110001100000110000011010100000000001000101001001010110101111001110101011010001011111111101011010000000100111100001011110011111100;
#1 $display("%b", po);
# 1  pi=207'b100010010111010101110101110010101001010001011111110110011110101100111110001011110000011110011000111101101100101101111011011010110110001011000010011000100101111101000110101001001000010010010000110100010000111;
#1 $display("%b", po);
# 1  pi=207'b100000000111000101001010100101010010101110000001010110111110011000011011010010001010001001111100010010110111110111010111011111000000000110100011111010001000100100001010001001010110011000110001101011101111110;
#1 $display("%b", po);
# 1  pi=207'b101001101001001110011100010101010000101001011110101111100010100100101000100101110011010100010100001011001101111111010101101001110110100000000101110000100101010100110000001010001000000010101001100100011101000;
#1 $display("%b", po);
# 1  pi=207'b001111110011011010010110001011001101101011111110100000000000001111100000000001000000101001011000100110011110010001001011111100111011101100110100100001101001011000011100101111110100100101010001011111011011011;
#1 $display("%b", po);
# 1  pi=207'b100110011000011000011001101101111001010001000110110011100011110000000000010100101100100010011011010010011100100111010101111011011001111110010010111000010011010011011100100000111100110011110110000110000100100;
#1 $display("%b", po);
# 1  pi=207'b010010101001100111100010010111010001100101001101111110011101101101001001111001100011010011010000101110110110010101111110110101101001110100101111101111100110100110101001110010101010111111010001000100011011100;
#1 $display("%b", po);
# 1  pi=207'b111011001010001101101000011101110010010110000000110101001111011110000011000001001011000100111011001111101110110010111010011110101100011110011001001011101101111111011110000101011100011010110110101111011111101;
#1 $display("%b", po);
# 1  pi=207'b000111011110110100111111100100011101110010111100110110110101101111010111000000000011000000100001101110011110110110010011001110100010001000110011001100011100110011010110001101100010110010001011000110000000101;
#1 $display("%b", po);
# 1  pi=207'b000110110111110001010001111111100001010110100001010101011011001110101111110110010101111100000001010000101010110100101011111110101000010110111100111000111101001110001000010001110100101001011100001100000100110;
#1 $display("%b", po);
# 1  pi=207'b011111100110000010000100000111101010100101001111011001100010100101000001101010111011001000011001101011011011000000100110111011111100010101000100100100111101000111101101110010101011011100111101100011101000010;
#1 $display("%b", po);
# 1  pi=207'b100111010010111000000100100100101001000110000111111011001000110101000011001010010001101011000001110111001011000011000110000001001000110000001101100111000101010010100111100011010011101111001010010011110101111;
#1 $display("%b", po);
# 1  pi=207'b011001000100000011011000111111010011111111101110100000000110111110001010010001000100011000101100000000000101100001111011011101100011000111001100000100100100111011100010110011000100000100011101001101110000110;
#1 $display("%b", po);
# 1  pi=207'b100011100001011110010110110110000000111000000011100000010101010111011011100100101110110110010111010100111000001010110100000111111110100100101100001010001110000101000011000000100011110001100111111000100111011;
#1 $display("%b", po);
# 1  pi=207'b101000001110100100001000111001011101100110110101110000001011101101011001000110110001100100111101110111111110010000111010010110010100010110001010101010000101001011101110001101000011101111011101001001101010001;
#1 $display("%b", po);
# 1  pi=207'b001011001100010111100110011010110101010001111111111000011101100000111111111011100011100011110100000100001000110101101111110100010011000111001011011000011011110111101010011010101000100111010011011111100010101;
#1 $display("%b", po);
# 1  pi=207'b110101010010011011101000010101111000111111100110000010010011110001101001010011100000110001001111110000001010010011111100001000010010011010011110000110101111011001011010100010011111001110110111010011001101010;
#1 $display("%b", po);
# 1  pi=207'b111100010010101011001000000110111110000011101001101100101010011110011111111000111000110110101000101110100111111110010101010100001100001101100010010100011101010100100111100101010001101000110011100101100100100;
#1 $display("%b", po);
# 1  pi=207'b010110010100111000110000001011110001100010100101010111000111101011010100100101011011001101001111101010111111110101100010111110111110111101010110101100000100111101011010001101011100001110010001010110001111001;
#1 $display("%b", po);
# 1  pi=207'b000011010100010110010101101101010011100010011101100111010011011111001101110101011000001000101000001010100001010001010101011010101001100001001111110010001000111111110110001000000110000110011001101101111111110;
#1 $display("%b", po);
# 1  pi=207'b100011000011011110001100000111110101000001111100011101100011011000000100100101111110001011110001111000011101001000110011111111100011010001111010010000110000110001001111111010110100111000001110011100001010110;
#1 $display("%b", po);
# 1  pi=207'b100111001010011010111110001111110001100111100011101100110011010001011010001001001001000100101101111111101110000101101000000111010001110100010101101111100101101000010111110001100100110110001110001101100010011;
#1 $display("%b", po);
# 1  pi=207'b001010001111111110111110000100001011110100011010110100111001000000101110111010000000100111000111010100010010011111001110110111101100111110110010100001010110000111111000001101111111101111001110101000110001011;
#1 $display("%b", po);
# 1  pi=207'b100010000011011111101011111101010011010001111010010011010001111100111101000101101011010101101100110110110001110000100000101001101110111111101100011011111111011000110001110001100000011011111100101001110011011;
#1 $display("%b", po);
# 1  pi=207'b100011111010011010000110000100110001010101000010011000000110011110101111100001100010011011100100000111001101100011000010001001010111111001100001010011001110110010000010001011110111011011000011001011001100000;
#1 $display("%b", po);
# 1  pi=207'b001100101111000000100000011011110110110110001110100100101110100110011110000110011011010110111011110010111010000111111111000110001001101011100100000110011001101110001011001011111001110001101111100101000001101;
#1 $display("%b", po);
# 1  pi=207'b000100000010111110010110010000011111010011000001100011100101110101001111101110100001100000100011100010100000110011001111001100000100001001000111011111001110011110010010110111011111110010011011001010100101010;
#1 $display("%b", po);
# 1  pi=207'b110101011110101111011010011011001011110001011110100110100101100011010100100101100010100000100101001111101111000101010011001010000110001000000111000111111101011110100111010010100101111001010001001100111100001;
#1 $display("%b", po);
# 1  pi=207'b111000000110100000111100001100000000111010111010110000000110000101010110011001000101110110001010100111011010011000011100101110010000011101010010010001111110101011110011011110100001010001001011001011000101000;
#1 $display("%b", po);
# 1  pi=207'b111100000111111011010010000101001101000101100001110001011001001101100111100100010011000101000011000101011101100001110001011100001011101101010001101101010110000011100111100001010110001011011010101010010000101;
#1 $display("%b", po);
# 1  pi=207'b100100111011101101011101001111010001101011001010101001111001111000011101101110110001010111110011010100010111011001001110101100100111110101110100001100000101001100001011001100101111111001111111010101001010110;
#1 $display("%b", po);
# 1  pi=207'b010001101010100101100100011000101010111000101000101101000100011001000010001101101000110101000000111110111001110100011110000101111000001111111010111010001001100001101110111011001100111101101000001110001000110;
#1 $display("%b", po);
# 1  pi=207'b011010001100000101010011011100100011011100111000010101000110111001011011100101001011110111111101011111010010000100011000011000111000010110100011010001010111001011110101010100100000111001111001100111010000101;
#1 $display("%b", po);
# 1  pi=207'b001010010111110001101001110010111100110101111101100111000010001011010010001101011011110001100000011011011011101010000010011011011010000001010010000101001111101110001011001101111111111000101011001101000010101;
#1 $display("%b", po);
# 1  pi=207'b110101000001100110011001001101011100110100000010111111000011101010000011100001000010111111010000000001100110001000111010100100011001000110110000001101110100100110111101011011010010010000100010001111010001010;
#1 $display("%b", po);
# 1  pi=207'b100110100101010010010000010011000001001100011100000001010110011101000110110011000101100101001111111110001101001001111100001111100011001111000101010000000011110110110011100110111011110000101111001101101110101;
#1 $display("%b", po);
# 1  pi=207'b110110001101011110101110100010011011010011110101010101111000101010001011101110100111001110000001100001101011011010101101010001101101000000111110110001111100001010010011100101011111110100010010100000001111111;
#1 $display("%b", po);
# 1  pi=207'b000111111101011110101010100011101101100010000000010110000010100100010100001011111110110010100111110011101010010101111010001101010000100010010010100101110110111000011110101101101110010111001001111111111100111;
#1 $display("%b", po);
# 1  pi=207'b001110111101010000011110011110000010001010011001001111100111111100001010000011101100100011011111100010011011011011011110011011100101011110101000001110011101110010100011001000001111001101000111111010010001000;
#1 $display("%b", po);
# 1  pi=207'b001011111011100001010110100011011010010000000001100101101001010001001000001100000111100000100011110011010000011001011110000011100001010001100010000110011101001100101110011001001001000000000000110001110101100;
#1 $display("%b", po);
# 1  pi=207'b011010110110101110111101100101100111111010101110100010110111110001110010001001110101001110000000000000010011101110011001000001010010100111001001000110000111010101011011100110101110011101101011011000001101010;
#1 $display("%b", po);
# 1  pi=207'b011001011100101100101110001000101110111100011010010000101011010100001100101101000110010001111001011100000100001111000110001101100111011011011000100100110101111100111100110011000000111100101111100110101101111;
#1 $display("%b", po);
# 1  pi=207'b100100000101101000100001101110101111111000100101111001011001111011111101010101101000010101010011101100010110001110010010000010101001010100101110010111001001000011111000111001000000100000101101001001011010101;
#1 $display("%b", po);
# 1  pi=207'b001110001111110000001001000111101010011101001011010111111010011100000101111110011110000000001011000101110010001100111110110001010000010100110100000111101110000111110110100110001001101000101100110001110000111;
#1 $display("%b", po);
# 1  pi=207'b010110000101010010111001010001011100000101010110110001111111000110010110001011011111011101101111100100101000000000011000000000111001100111100100001110010111110010110100000101010101101101110011101000101001010;
#1 $display("%b", po);
# 1  pi=207'b001011011000010111111110101101001100101000001000111100001011001101011101000101100010110011000100100101000010111001011100100101011010000101100110001111010101101001010000000000011111100011110001011101011100110;
#1 $display("%b", po);
# 1  pi=207'b001100101100110111101111101100001100011100111100001110001110000001101001011101111100001011010111110101010101010101110111001100110101011000001110010000010100100011101000001010101010011100111011110111011000010;
#1 $display("%b", po);
# 1  pi=207'b000110111110011100111100011001110101010011000110101011100101101011011101010011111010001001100101010011101110111000011110101011000101011111010001100010010010100111100100000011101011111110111111100011011001011;
#1 $display("%b", po);
# 1  pi=207'b011101011011000111110110111001101011010111101100011111010111000111000010011100110000000001011011010001010000010011011010000011011001000110001000001111110111101001000101000101111010011101010011101001000111101;
#1 $display("%b", po);
# 1  pi=207'b000111001010000111110001101101111000001101111101111101101001000111110000010000100101011000101011100110000000010000110001111000110110000000000110001110000011001100010000011100101010100111000101100000010101101;
#1 $display("%b", po);
# 1  pi=207'b111010101100101111001010110101010000000000011101101110001100100111100110101110111001000111101011000111000100011001011010101101110001111101010111101110011011011011000001111001000110001111000110101000101010011;
#1 $display("%b", po);
# 1  pi=207'b000101110100000111110000110000100110101101111001101100001001110101001110000001001000001101101000000000110000110100100000001011111001000111110010001011100111100110000100010011110000011000011010000100110011000;
#1 $display("%b", po);
# 1  pi=207'b101001111100101001000001100001101011001111001111010001111110011001001000010000111010000101001010000111000101100101110001011011101111001110000111011111001101111101011000000100001010100011110101001000100101000;
#1 $display("%b", po);
# 1  pi=207'b000000011000100110101000110010111111100010010001100010011111001101001100000010001000001101100000010110110111001000001011000010001001010000011100110111001111001110001000010100010011000111111101111001000010011;
#1 $display("%b", po);
# 1  pi=207'b001001111001111100000101011011110100101000110010011101011100110111001111011001010011101010000010010011000011110011011101111101010110010000100011011000111000111101111111010010011111001111111000100011010110001;
#1 $display("%b", po);
# 1  pi=207'b111011010111010010100010010000110110011110111111101100100010000010110000011011000100101111001111011011101111001111010111101101000100110111010110101000110110011010100100100011010001111011101010100000101111111;
#1 $display("%b", po);
# 1  pi=207'b101010010110100110110011101101101111011011111011000011100011000101000000111001101000010110110100101110011000011101001110001100100110011110110111111101010001010010011100100101101001111001011010111001100101000;
#1 $display("%b", po);
# 1  pi=207'b111001001101101010100100010100110101111010001001001110000010001001001001101111100010110010010111111110011101000011101010110010110010111111000010101001000001101110100100101100101110101100000010011101101111111;
#1 $display("%b", po);
# 1  pi=207'b111101001100011100101011100000000000101011010110111100010001111101000111010101101001101111010110000110001110101111011100001110100100000011100000010111011110000000001011111111000000001001101010110001011111101;
#1 $display("%b", po);
# 1  pi=207'b001101011001110110010001001011000010000000110010110100010011100101000100011010100100111010110001101100110101101111110110001111100011110110000010110011010000110111111101111100110111000000111011001001101010001;
#1 $display("%b", po);
# 1  pi=207'b110000000111000100010000100111111111100100100111110000001111101011110101100011101110110011101011100000001111111001000110011011111111000100010000000000010011100001011110011001100001111101000111000100100010011;
#1 $display("%b", po);
# 1  pi=207'b101001000011000011010010010101001000000101000001110010110111000111011100011101000100001110010100100111010100011001010001000100000001010111100110011110101111111000101110111001010011110110101110110010000111001;
#1 $display("%b", po);
# 1  pi=207'b011111011111101111000001010000111111111111101101001111011010010001000101100111111001000011100000111010010101000000010001001000000011101110101110000100001011111010000011101100000010011111101010110100010011100;
#1 $display("%b", po);
# 1  pi=207'b000100000010011011101001010010110010010110011001000011110111110011110110000000010010000011101100100111010111000011011111101011100010001101011101101011010101100100000110101100001101010111000100001110010111010;
#1 $display("%b", po);
# 1  pi=207'b101101000001100110100001111110100101001001101100000011011101110111010000100111110010000011111000010011011101011101100000111111001100001100101011000100000110100110101100001000100010011101110110110011001111011;
#1 $display("%b", po);
# 1  pi=207'b001101001101110110001010100001001011010000100001111110001010000100001010110000101110100100000111111111100110010101110110011001011001110111100111000011111011100111100100000011101110110111111110101000100011001;
#1 $display("%b", po);
# 1  pi=207'b111110110101111010001101110001111101011011111101100100001000001101100000111100010110111111100101101011101001101100101011011110011101001000011000100111010010000100000001001011100001110110000110100001111010111;
#1 $display("%b", po);
# 1  pi=207'b000000001101101011111001010110111010011000110010111110100010111000111001100010010011010000101001110011010100000110000101000110001101001000001000110011001110000111100001100000111001110101011001001001000010100;
#1 $display("%b", po);
# 1  pi=207'b100110010110000100101100100100100111011110110001111111000111000000101111010111010100110001000110011001001010000100000100110000010011101010000000111010001110011010111010100001101100110101000101110010100011000;
#1 $display("%b", po);
# 1  pi=207'b000111011000111000001101001011001101101111001010101000010001100101100110101001001001110101101110001101111000000111101001101000000101111010110000111100011000110100000101110001111101000111111100000010111011000;
#1 $display("%b", po);
# 1  pi=207'b010100111111011110000011011111100101101100101011010101011111110011100111011100011100000100101111001001111011110000011101100000011101101101001001111100001111011101100100110010001010000100010110000100111000001;
#1 $display("%b", po);
# 1  pi=207'b001001101110101011110010000100100110000111010101001101111011111111001101001101101000100001101001101111001010000101111000100100111010100001110100100000110000101111110110010100000111111101000100100110110001100;
#1 $display("%b", po);
# 1  pi=207'b010010000010101110011010100100000110110100101111101111101010001000011110000100111010001010101110001001111100010101000010000000101010111001001101111101101111011110111100011001000110100001010011000011100111000;
#1 $display("%b", po);
# 1  pi=207'b111000000101000010111110010111100111011000011110100101011110001001011010111101100110101001100000010010001010100000100111001001100001001100100010010000110111000001111100101101011010110000100110111011010110000;
#1 $display("%b", po);
# 1  pi=207'b010111011110000111110100110111100000110111011011100111101111111010000001110111101010110100100010010010110101100001100000110100111010111001101011011001110110100110011000000010101101011000001111100110010111000;
#1 $display("%b", po);
# 1  pi=207'b101111001001010110111100111010011010100111101000010110011000100101001110111110000100110000101001110101110111100110110111001100001001010111010000101000000000001101010010001111101111111001000000101100011111000;
#1 $display("%b", po);
# 1  pi=207'b111010110001110000000101100010001011100111000001110000100010001000001001100110010000000010111010000010000010010001001001010101010110111101000001100000000000111001100100110110001101100010100010011101100011100;
#1 $display("%b", po);
# 1  pi=207'b101001011101101000100110000111000011100001101001000001011000000000101001000101001000110010010001011101110101100011011010010000001100010011100100100000100000000100100101111010111001011110011001110000100000111;
#1 $display("%b", po);
# 1  pi=207'b011101001110011011111001100010010110011110100011011010111111010101111101000010110101101010000011000001100000010001111000000100001110101111111111001001010011010100111111100010101000001001111010111101110101000;
#1 $display("%b", po);
# 1  pi=207'b010000111001101100001101011100110101111010110000001100110111111101111001000100110001111100011000101001010011100101101101011010110001111110110100110110111111010001001100011111101010100001000011011110100011111;
#1 $display("%b", po);
# 1  pi=207'b100010101100011101000101010001000001110100010010111100111000010100111110001110010000101001110101011101011100111010001100011000001000010001011000110011111011101111101011011011101110111101100111100000100110010;
#1 $display("%b", po);
# 1  pi=207'b011010000101101000001110010001001010000000101001110111111001111011001111101111000111011100101111100011110100000101101001000110101011111100001111000011110101000100011110100000110001100000110111001111011110110;
#1 $display("%b", po);
# 1  pi=207'b000001001010010001100011100010010110101001011101100101100101010001000100111001101000111001010001010001000110111111000011101111010101100010010010010000000001001110011010111001010001011110010101001001001110000;
#1 $display("%b", po);
# 1  pi=207'b001010100001010100110011110100100101111001001010111110010010110011011111011100001111110010010010111000000111101010011110000001000010101011000000011110011010100001111010111101100111010010101001111010100101010;
#1 $display("%b", po);
# 1  pi=207'b001101110111001010001010101101101100010100001000101101110001011111101011100011111111010001101110110111001010100001101100100101111110100101110010000101011101101000110001011101110101110001101011111101101001011;
#1 $display("%b", po);
# 1  pi=207'b000100111000110111110010100101101101111011110010001001111101100101011101000010110100010100010110110100111110011011011100100110100000001010011010101100110000100000010011111100010101001000000110101100110011001;
#1 $display("%b", po);
# 1  pi=207'b011111011011100111100110101101111000001011100100010111111101001111000101011010110101110101000111010000011110000101100100101010001111010000010010100101111110111001111011101011000010011010101011000111111011100;
#1 $display("%b", po);
# 1  pi=207'b010111001101101011110110010110100000101101001000111111010110010001110110111101010000101000101011000101100110101101101101001001001101000001000010001110011010000111001100100110011111000000101000011011000000000;
#1 $display("%b", po);
# 1  pi=207'b100100011010010000111011100111011000010100011001001001100010100100101100001010101011111011110001101001011110110011000001001011100000110111011111110100110011100001101110100100111000101111000010100101110010000;
#1 $display("%b", po);
# 1  pi=207'b100111110110010000011101100010100101100101001100011100010000101100111100010010010001110111110110011111101001000001110100000000000110111001100111010100111010111110101101011011110101010111110101010110100010000;
#1 $display("%b", po);
# 1  pi=207'b000010111000010101111110100000011010001001101101101001110010110110111010000001011100000101100101001110010110000100110001011111110111001111101100111000100100011101010011100010100111000110100111000010111100110;
#1 $display("%b", po);
# 1  pi=207'b011101100100010111000001111001011111001101011111101101000110110111011100001101100100100000010011010001111000100010000110011010111011101110000011101100000000111011011101111110100011111111101110011110010100010;
#1 $display("%b", po);
# 1  pi=207'b111010100110100001011101011100000100100100110111011000001010101111010101100011010001111101001011100010110110000011101011000101011001010011010110001001011001001011111111011001011001000111010100100111110111011;
#1 $display("%b", po);
# 1  pi=207'b000001110001000000100001000011101111001011011011110000111101111100100011110011100100000101101011101111000100111010101000111100010010001000000001000100000111000101001111011010110000101110010101001011101101001;
#1 $display("%b", po);
# 1  pi=207'b011001001011010101001010001001000110101110100110101111000110100000101100010010010000001000011101000011101100001110010101010000101111010001000101010011010000110111110110101010001100011100100101100010001001111;
#1 $display("%b", po);
# 1  pi=207'b000110101111010001000011101111010001001101100111101001010010011100111010101010110001001100010010111101001100100011000010110000111101010010101111011110111110111111100001001110101111000111011000111001100010010;
#1 $display("%b", po);
# 1  pi=207'b100010011011101010110101010000111000000011111110000100110101100001101111011100000110110111011011011101001111101010100011100010100000010001100101111011001110000011110000110000010000110101001000000001100010111;
#1 $display("%b", po);
# 1  pi=207'b000000110110011001101011101000011101001011101111001100000010111100010011111001011000010110000001000100001000010001001010011100011100001011000110011010010011000101100110111001111101001000100011001011110111000;
#1 $display("%b", po);
# 1  pi=207'b100011111111110110101001101101101000111110011110000010010110111011000111011100100110001001001010001011001010101000010111100101100110101011111100011101101011011001010101000000000101001101110101010000001100110;
#1 $display("%b", po);
# 1  pi=207'b110010001000100101100110011100110100100001100110100110111011101000110000001111000001111010001010000001100111001111111001010000000000111010110111111100001000011100011111101000111001001010111011001100010010100;
#1 $display("%b", po);
# 1  pi=207'b101001101000100011010111010101011001101010011100110111001010110110100010110110011100011011110000111100101001110110011010011110010000000010110011011101000101011110111101000011001100000111111111001111110111001;
#1 $display("%b", po);
# 1  pi=207'b000101000110110100100001010010010101000101110101000110010111111110110111011010111111111011111111110001111101110001101101110011111110100010110110110011100011110101111100000000000001111000010111001111101010100;
#1 $display("%b", po);
# 1  pi=207'b111001111001100110010111000011011100001110011001101100011011101011000010010001001010101010101110111011100110111101000100111001101010001010000000100100110111100111010001000001001110000111110101000100000101101;
#1 $display("%b", po);
# 1  pi=207'b011110011001100100101001101111001100001101101111000111011000111110111000100110110111101001010111001001010000101001001111110011110011111011000101100100001011101100001100110111110101110000100110001011010010101;
#1 $display("%b", po);
# 1  pi=207'b100011000010011010011100001001001011111010111000100000111010000010010101100111010111111000100011100011110010101000110110101100000110101010010111011101110111011001101010011110000000010110101001000110111101110;
#1 $display("%b", po);
# 1  pi=207'b110100111110101100010001010101001000111111011010010011110001110001101111001100010011110101100010110111011010110101110001000101100010011001001011110111101010011001000101111101001100000100100110011010000101001;
#1 $display("%b", po);
# 1  pi=207'b101001000100100111110110101001001010000111111011001101011110000100001010111000101101010101110001001110111011010100110010011111001111111100101011010001101000110000110110100010100111110000000110101001011110011;
#1 $display("%b", po);
# 1  pi=207'b001101010110111110010011011010011101010011110110011001111110001110101000011001011100010110110000111000010000000110101010101010101001111111001011011001010001111110111000111111011111111111011110100100111000001;
#1 $display("%b", po);
# 1  pi=207'b110100000001000111100010010011000001111101100011100011110110110101000101000010001101110101000100011011000001010101101010100100110100010111000100111100111101111010011000101100111101111011110110110000011110111;
#1 $display("%b", po);
# 1  pi=207'b101001100000010001111000100001100010100110100000101110011100000011111010110011011101101111101101010011101111001101110010000011101011000000001001111101011000011111111000001011010011111111001100001010111001011;
#1 $display("%b", po);
# 1  pi=207'b010111101110111011100001111101100000101101111110110101101001000111001100100110101001111010001000110001000000000000000000101101010000101111110111001100001111110110110100110001000110011111111111011011101101000;
#1 $display("%b", po);
# 1  pi=207'b011010001110001101100011101001100001111001000111110001101010101011001011001010001101101100111100011111001101111001101000001001000101011001100101110110111111001101110000111011100001000101111011100010101010010;
#1 $display("%b", po);
# 1  pi=207'b110100111100100110111011111100000101001100000110010100111001001010011011110011010100110101011001001001110000111111000111000001000011001011011000100011000110101111111100011110011001001010110111001110110111100;
#1 $display("%b", po);
# 1  pi=207'b011101011001100101100101111000000110111011011111110011001001100000000110011010001001101000010001011001010000111000000101101011001001000101110001100110111110000010111101000000001011011100011111001001101111100;
#1 $display("%b", po);
# 1  pi=207'b111010111010110011001010001101111001100001101001000101011110100010001111001101111101100010011100101001110111001011011111111010001011011110100110000000100001111000110010001011101111000001010101011101001011100;
#1 $display("%b", po);
# 1  pi=207'b010010011011010111111011011110111101010101001101100111011000011011110111101011011110101100010000000100001001110000000101011001000011011111100111111001100010111101110001010001011000100101111010001110110101110;
#1 $display("%b", po);
# 1  pi=207'b101000011000001010011010011001100010010011111111110001101011010011001100111011111111110100110101100011010110100001011111101110101101011100001011001000000110101011010111101111001000101110101111111101010010101;
#1 $display("%b", po);
# 1  pi=207'b011001111010011001101010101001011101101001010001110000101110011101110001011000010111100001001010010000001110100100010001010011100001011101000101010001001111000110001101111100010111011001100010010001010100011;
#1 $display("%b", po);
# 1  pi=207'b110111101000101001010101010010001011011010101110100001111101001011110100111000011001001000110011011110001110001010011110101100001011111011100111111101010100001000110111111111101111110110111000101011000111111;
#1 $display("%b", po);
# 1  pi=207'b001101101101100010100110010001011100001111110010010001011111001101001100111111110110110110010101111101111010001010000110110101010001010110111011110010110100100111001010110100110110101010011010100111010111101;
#1 $display("%b", po);
# 1  pi=207'b011001101101000101110011110101001100111010000111000000000101111010100010110101010101000110010111111111111011101010110110111011100100001110000100011110000100010101011010101011010010101101110101110101000000010;
#1 $display("%b", po);
# 1  pi=207'b000111011110101010010100111101100110110100111110001111011001101010101011101000111001001111011001111000110101001000111011111100100101111100010100011110010000110101101010100011011011000000111110001111001010111;
#1 $display("%b", po);
# 1  pi=207'b000100111110001000111100111110111000100000000110000011101100111101001011111001110110001001110100110100011000111010100010000011000011001010000110110001100010011000000100010101110011100010011001010110000000110;
#1 $display("%b", po);
# 1  pi=207'b000010010001111001100001111101010011101000010001110010011101011001111111101111010000001111110000100110110011101111000000110101010100111011111011001111100001000010001010111111101110000001101110111000001000110;
#1 $display("%b", po);
# 1  pi=207'b011010001110001001011100001000001110101001000100000110110010000010101101110011001010111010001100010110110101001001111000011001010110100000010101001100000110100010011101010110000000000101001000010101001011111;
#1 $display("%b", po);
# 1  pi=207'b100000011001111011111110110110110100101111100001110111101111100111110010101000011100111010010110101110000010011011011010001011010110100000111010010111000101101011101001011101000010011010010011000111100111001;
#1 $display("%b", po);
# 1  pi=207'b001101001010000000001010011010011011100100101001110001010111110101111001011001100001101101011000010011111000011010100011010101110010110000111001100110001110100111000100010101010101110011011110100101111001011;
#1 $display("%b", po);
# 1  pi=207'b010101111100111000011101001000101001001100111101101110101000000111000000101111001001100010111110101011111011110110010101000111001111111111001010110000100100010111101000010100000111000010001110111011001111001;
#1 $display("%b", po);
# 1  pi=207'b111110000000011010100011101110010001100010011010101101110000111010001010100111100111000000110000100100011010110011110001011101011111001101010001001110110110111101010111000010101011000011110010100010101100010;
#1 $display("%b", po);
# 1  pi=207'b000000100001100001100000101011101111110110100010011111010001010001101000000100010101000011101101010011110011101111000011011010000101101110001001111100110110000101110011010011100001010010100001110100011100010;
#1 $display("%b", po);
# 1  pi=207'b000100011011011111000001111101101000001010010111111000110101001011011110110000100011101101011100000111000011111000101111011110110111100010111011101011100010101010011010011011101000110000001000111110010100001;
#1 $display("%b", po);
# 1  pi=207'b000011110101111110110001000100100100111110111000110001110110010111010110001110010010000010111001010111011110000100100101101101111001010010110110001000100101110001000000000000010001111101000010001111000100000;
#1 $display("%b", po);
# 1  pi=207'b100011111001101101001110100111000101011100110000111100011101011111100010100010011000001111110000000010011100110110110000100011101110011110001100000111010101001111011110000100101111111001000110011110010001110;
#1 $display("%b", po);
# 1  pi=207'b010111100100010010010111100110110100100111011011011100111010100101000011000011101111001001011101111011000100010001111001110111111011100001001101010101110110010100001101010111101001000001001000100010100011111;
#1 $display("%b", po);
# 1  pi=207'b010101010010100000111111100100111100101101110000011101010100000011101100011110000001101010100010111100110001110111000010000010101101110111101011101110111110000000101001011010110011011011100001101110100001010;
#1 $display("%b", po);
# 1  pi=207'b001010001111000001010000110101010000110110001000010010010010111111000011100000101100011010010111100000101011001010111100100011100100101101000001000001101111101010111011110010010000011001011101101010111000110;
#1 $display("%b", po);
# 1  pi=207'b100101000011010010001001100111011111010101100110011100100101011110010001010111010110101110000011111110011001010011010001000110111011111000010111111111000101100000010111010100010100010001110011000100010111111;
#1 $display("%b", po);
# 1  pi=207'b001000000110100001000001001111100001001111001010001011010101001000111110000010001000010000110011111111111011011010010010010011110110111100011111101000110100011010000001101001111000000010100000011110001011100;
#1 $display("%b", po);
# 1  pi=207'b110000010101110110100110000001001101111101000111000100111111001110111110111010101110010111011011001000101100111001010100101001101101111101111100101001111001000111000001111111111001011000010000111110001110111;
#1 $display("%b", po);
# 1  pi=207'b011000011000010001011011111100111101001110010011111010000100010110111010111011100010111110000011010101111001100001100111100100011111011101100010010100011101100000111111000011111001000010011101000110011011110;
#1 $display("%b", po);
# 1  pi=207'b000111001101101111110010111001000000100011111110010011111010100001010001000111001110101101000100101101100010111001101100011011100100011001100001011110101001111011010101101010011100001010110101100001000110110;
#1 $display("%b", po);
# 1  pi=207'b100111010111000111011011100100110101001101011000110010001110010101111011111001000000101011111101110111111110001010001001001010111011100100010001010111101100011101000100001001110111101111011000110001100010011;
#1 $display("%b", po);
# 1  pi=207'b000000101001101011011101010111100111001111101001010100000110111000001011010010001101110000001110000111100110011110001101100001011111001001010100010111001010110101110100111001011010010000100100100000010101101;
#1 $display("%b", po);
# 1  pi=207'b001111110011111100011010000100010110000010001011111010110100010101110101010110011111100000000110010110111100011011011100110100101101011111111110110110010101000110111100000000100000010001111000001011001010100;
#1 $display("%b", po);
# 1  pi=207'b011101000110010111001110001000000110011111011010100000000010010111010110011010000001000001001100001100111011011110010000111100001101100110011100011110111010110001111000100000111100101101111110110000001000011;
#1 $display("%b", po);
# 1  pi=207'b100111100101101001100010100011001001011101000001101011001001110100110001011101000111100010000011100101011011010011100011000011001010100010100101011101111110111100001011010111110111001001010101101000100111100;
#1 $display("%b", po);
# 1  pi=207'b101001110101011011110010010010000111101110100000001111010100001110011011110001101101000000110110011100000110010011101001010010000010100110111111111001101101011101001101011000111000110000001011111111001011100;
#1 $display("%b", po);
# 1  pi=207'b100111001100101101100101010101000110000101011001110100100000011010000110111100000010010100000011100000010111010111010000110110011001101100111011011010010111110000011010010101110101100011101001111100010000011;
#1 $display("%b", po);
# 1  pi=207'b110111011011110100001111001010110011111100100101000111111001011100000110100101110010101000010101101100001000100011110011000010001110100110000001011100011101110111000101111011000001011011000100010001111011110;
#1 $display("%b", po);
# 1  pi=207'b111010111010001000101000111001110011010100100101100011111000111011101110101001011001101110011111111100100100101001010101011011100010001001100000100111101011101010100000001101101101010000111001010100000000000;
#1 $display("%b", po);
# 1  pi=207'b001000010001100011101001001001011011010110110001101101100110101100001011000101000110111110101010110000101001111001100010110001101000001001001101011001000010001010000110000001011010011001000001011110000001010;
#1 $display("%b", po);
# 1  pi=207'b010000101000001010111110111010100000110100111000010100100111111100011110001000001001100111100001110101001000011000110100001001000000111011001000100110001010110010000010011111000010110000001101111000100001000;
#1 $display("%b", po);
# 1  pi=207'b000000010110011001001111010001100101010101011000001110110010001000101000001001110000010001000011101000000100110011111000010100110011010101001001010111110100111001001000110000010100011111100101001101011001000;
#1 $display("%b", po);
# 1  pi=207'b110111000001011010011101011010110110010101111101010100101011001001000101111100111010000000010101100111101011000110111111000000110101100010010100010101110010110110100000111101100101101010010011000001110011011;
#1 $display("%b", po);
# 1  pi=207'b000100101010100000111000111011000110111001001011000110111010011101101110010110011100100110101000111011100111111010100111001111101011111111110000010111001111111111001110010001100001001001011010111111101111110;
#1 $display("%b", po);
# 1  pi=207'b000110011100011011110100110110011101101101001100011010010011110000000000010010111011101100100100111100101110000101010001111111000101100010001101001101010001110000100101110000101000110110111010000011100101011;
#1 $display("%b", po);
# 1  pi=207'b000000110010001010100101100000110010001101111011110110001101111000001000001110010110011111111001111101000000000110100100011110110101110001101101101000010011001001100001101111010101001010111110101000001010000;
#1 $display("%b", po);
# 1  pi=207'b011100100010011010110110111001011100000101000000001010011010010000110010101010111100100101000000011111010001011100000110110011110001010000010010000101010010101011010010011000010000001110001111101101101111001;
#1 $display("%b", po);
# 1  pi=207'b010111011111100111110110110100101110001001100100011110101110000000110111110101101101110100110000010001110101110000011110011111001001000011000000000001110000100011000101100001100011101111101010110011010000001;
#1 $display("%b", po);
# 1  pi=207'b110111000100111010101101100101011110100011100111010100001001111101001000010000000000011011100111100100101101111110111010101111001110111111001100110000000110000111000001110110001010110110111101010011110100000;
#1 $display("%b", po);
# 1  pi=207'b011101010010000100100001101001010001110001010010100110010011101110000010111101100111110000110100100011111100110001011101000111110111001010000111010110000111111010110001001000100010101110100101010001010010000;
#1 $display("%b", po);
# 1  pi=207'b010110100101101010000010101111001010001011010000011011110010110110001111010101101101000111110000111100010110101000000001100011010101000100110001011010001010010100110101111001010000100010000101111001001110100;
#1 $display("%b", po);
# 1  pi=207'b111111001101111111111101011100111100111111100110010000111101000000110011000001010010010100110110101011001100100100000010110000010100000011001000000101111010010000000010000110001010100111110111010011111010100;
#1 $display("%b", po);
# 1  pi=207'b011111111011110010111011001111011001100000011111100110001001100110100101001000100100100010111100101111100111001111100010000010011101101000100000001111110110011101100010011101111101010000011111010010100001011;
#1 $display("%b", po);
# 1  pi=207'b000001110110101010101000110100100100001000101010100001010101101110011010100101100100000110011101100010111011100000111010111111100011111101011011000010010110110010100100000111110100111000000111111100110001101;
#1 $display("%b", po);
# 1  pi=207'b001111001011001011010011101011011000011011101100111010011010001100001000011011100010001000001111001110110011101111011010101011011001101101111010010110010000011000000111111100000011111011000001000101111001010;
#1 $display("%b", po);
# 1  pi=207'b011000011000000000110110100110001010010000000010100100010010010101101101000111010110100110110001010110100101100100010010100001110010110100100101100111000100100101100001000010011000011110011111101111101011111;
#1 $display("%b", po);
# 1  pi=207'b011011010101011101100011000001011100110000001011110101001111101100000011111000001011101011010000011111111001011010010100101110111111100101001010101111000110110100110110000011011001101111010011001001010101011;
#1 $display("%b", po);
# 1  pi=207'b000101100011011100101001100001011011000011100101101011001000101011110110111011100011111010011001011111000101101110100010011110110000110011001111100010111010110100111000111110101111110010111001101111101101011;
#1 $display("%b", po);
# 1  pi=207'b000101001000111101110110101010001011010010011010011101101110000011000000100011000001111000100001001001101010111110001111001101100101101100001011110111001111001000101001010111000101111010000010110101011011000;
#1 $display("%b", po);
# 1  pi=207'b000100101010001110010101000110110110010101111000100001101000010000001001110111010101110000110001000011001011010010111011101000101001001000000001110101001011000001110110000011011011101010110010101011001100111;
#1 $display("%b", po);
# 1  pi=207'b110111101010111101000011010100011011111100001111010100011111100110010100100111100110010001111011010011111010111101111000101100010010011000101111010001101000001101000100111000110001001110000001110001010001010;
#1 $display("%b", po);
# 1  pi=207'b011010000111011011000001001101011010111000010110001111110011001101100011101000000000000101000010001110110110111110010001011110111000000111101110111011111011000000001111010110100111110100001101010111010111000;
#1 $display("%b", po);
# 1  pi=207'b111010111010001010000100001111011111011110011010011011011000010010000111011000001100000100011100011010111000010010111010010101001100000000110101010000111100111000010000111000010011011010101100111101100000010;
#1 $display("%b", po);
# 1  pi=207'b101000111001000111011011111010101110100001000001000100100000011101000010101110000000010101101111011110001000000100010001001100010100111000010011001010000111111101001101101110001011011101011001010000000010010;
#1 $display("%b", po);
# 1  pi=207'b100011111100001000000101001101010110010001100101001110110010110000110000011110111001001000101100011001101001000110010101100111110011101011100110111100100001100100010101111001110001110101110010011111101010111;
#1 $display("%b", po);
# 1  pi=207'b000111010111111000011111100011110100100011101100101101110111001110100011100100110101010101110100111000110111010011010011111101111011110010000101110110100100010000101011101010100010001100001111100110100101000;
#1 $display("%b", po);
# 1  pi=207'b101100100110101100110100110110000111100110101110110101100111110111011110110011111111111001111101110010001101101001101010011001001111101111111010110011010000111011011111001110101000101001110111000110110000010;
#1 $display("%b", po);
# 1  pi=207'b011011001010111000110011010000000000000001011010111100010110100010000000010010011011010000111011001100011101010110000111000111100100101010011001110111111010111110011110110000111101101010001000101011011110000;
#1 $display("%b", po);
# 1  pi=207'b111111000001111110011111000001011111111101100001001000000000011110100100100000111101001101011111000001001111101111111001010011000101011110011000000011100110100010110011110001001111100101101001010000100010000;
#1 $display("%b", po);
# 1  pi=207'b010010011110101100111011100000000011000100101001100011000001001001000110010101101111111110000000010101110111010100010000000000111101111000010111100111100101110110001110101001100000111010011000010111100111001;
#1 $display("%b", po);
# 1  pi=207'b100010001001000001010100001010101010011111001101100000101000111010111111000001011100001100101111110111111100110011111101000110010100000110010001100101011111111011101100110010000000000001101100111110101000011;
#1 $display("%b", po);
# 1  pi=207'b101101101000010110011000101100001110001010100100011110111011100001110011100100010000101000000101100101111011111000011111010010100111000010111101100100110100100010010101001111101000100100011101111100000010010;
#1 $display("%b", po);
# 1  pi=207'b111101001110101101011101110110101001100110110010101101010111011111100000001010100110001101010000011011101101000101000000111111001111101010111101100001010000101000100100100111001000110001001111011110000111100;
#1 $display("%b", po);
# 1  pi=207'b000101111000000000010000110000010111110000101011011010001110111011010110011111111110000111000110100010011100110010111010011101001010010111001111010111110100000011101010010111101001111100011110100000101010101;
#1 $display("%b", po);
# 1  pi=207'b011100101110100001101010011000000010110101000110011111001000110100100100001110111010101000000000001110100100110001000100100011000111111100111100000111110011001010010000101111001000100110100110011101111100101;
#1 $display("%b", po);
# 1  pi=207'b001100010010000001001100000011111000100110101001001010110010011110110011111001111010011111100100100011110111111101101000000110010000010001001000101000010100111100101010000101101011010000010010101110110100011;
#1 $display("%b", po);
# 1  pi=207'b111010110011010111111110001111001110100111101110111110111111101000110110000111011011111110011111010011110110110100011110011111101010011101001001011111010100100110000010010001001100000000101000000001001111110;
#1 $display("%b", po);
# 1  pi=207'b111111110110100110010100100001100001110001011101011001100011010001001001111000101110111110111100101001000101001110111001111001100101011101101100011101111101100100100001111110110010001100110101100100101011100;
#1 $display("%b", po);
# 1  pi=207'b101000011000000001110010010100110001000000100100000010001111001000100100111101010111001110111110000111000101010110111110101010100110010110101001010110010001101011111000101011101001101101110110111010101001110;
#1 $display("%b", po);
# 1  pi=207'b100010010100001101010111011100101011011111111101101111101111110101110001010001000101010110000101101111110010100100101011010101001001101010101011000100010110000010101111100010100100011101010000010010010000000;
#1 $display("%b", po);
# 1  pi=207'b001001100011000111011000011101001111010110010100001100100100110111001100011010100010000010010100111100110001100000011001000100011101100100010000010110010100100001101110011101001111011000011110101100010111100;
#1 $display("%b", po);
# 1  pi=207'b011101011101001011100101000011001010000100101001101110001110010100010111000100010000111001111010000000000101111000101010001001111011111110000001110011101110001101001001010101111000001000110010010001011110000;
#1 $display("%b", po);
# 1  pi=207'b101011010011000001001011001100011010101011010100010001010000001010010011110011010100001111010000101001101101000100011010000000111000111001010100000000110111111100111101001010100011100001100101100011010011111;
#1 $display("%b", po);
# 1  pi=207'b001001011110100110011111110011100001001010011001100101010010000110101110011110101000010111110011001010001111010111100110001011000110010101011010100010010100010011101100100101101100001110001111100110101111000;
#1 $display("%b", po);
# 1  pi=207'b110100001101000111000000011110101111010110001011001001111000000011010001011001000100000000101110111001101101011110100010011011110001010110001100110111101111001100101100001101000010100010000010011100000001010;
#1 $display("%b", po);
# 1  pi=207'b111001101000011100111000010110000011111011010101001110100111100111011111110100100111001101110110001011000000111011111100010011100110101000100001110011110010100010101010101010110000100001110011110000111110100;
#1 $display("%b", po);
# 1  pi=207'b101101001111100001001110111111111110010101111011011010101011010000000100011000101000110110001000000011100001111100011010101000000011101001001110111010001111001110111001110000100110101001100011011100111100111;
#1 $display("%b", po);
# 1  pi=207'b000111110110100011101011111010001001010011000111100111001110011110001100101110101101000000001101110011011001101101100101111001110001100110001001000111100101101011000001000001101111100011000111000001111110010;
#1 $display("%b", po);
# 1  pi=207'b010101011001111111100011000111000000100100111010111000111100000101101000011010100110011001111100001110001110101100101010011110111011111010001110110101101001101100011110010101100110011000001100101001010110001;
#1 $display("%b", po);
# 1  pi=207'b000000011111111011101100101100000011111000101110100101000101011010110010111001000001110010000011010010000010110001101100100010111011010100000001001100000001001000001111011001101100000100111111100110111101001;
#1 $display("%b", po);
# 1  pi=207'b110101010111111100011101000110101111110000111111011000100001001100101001110001100001000111000010111010100011010011111001110010110111110110010001110101101010000001010001100011110011001100101100100000110011101;
#1 $display("%b", po);
# 1  pi=207'b000001001010100011001001011010010100011000101010011100110100010001010011111010110111100101001000110101011111100101110101101011100001000001111000110010111111000010111111001100010011001111001000101110110000001;
#1 $display("%b", po);
# 1  pi=207'b001110110000011110001101001101001011111010100101110111001001111011100101110111110100111101010101110001110000100011110111010011000110010000011000001011001110100001010100001000000100001001100001001001110001101;
#1 $display("%b", po);
# 1  pi=207'b101001100001110010000100111010110000001011010011110110010001000110101101010111001100111011001000101011001111001101010110000111000001000000000101001000011001000100011100001100110001101001111001110000111111101;
#1 $display("%b", po);
# 1  pi=207'b010010010110111101111001110001100010010011010000101011010101001100010111000110000010110010011000001100101110100110110001000111000101001111010101001010000001100101011110000101100111101010101001010010101101110;
#1 $display("%b", po);
# 1  pi=207'b111001010010110101101111011111111001010111111001001000000011111000001001101010100110011111110011101001111100011000011010111100101011001010001010000101101100001111110011000100110011001011000000001101111001000;
#1 $display("%b", po);
# 1  pi=207'b001010010010000111000100100110111110011110111001011010000001011101111110111100100011010110010010101100001011000100010110100110010010110000011110011110110011100101001101000101000111011100100101110100101001111;
#1 $display("%b", po);
# 1  pi=207'b110110110001111010111010000110010110100001110100111011110011110101101000101111110101110110111010011001011000111010101110001001010111110101011000000000100001110110110000100110001111001110001110111110011110001;
#1 $display("%b", po);
# 1  pi=207'b000101010010100110001011100110000111000000100010000010101010110000110111000100101110001001011010101110110101011000100100101010101011001101011000100110000001111000011111101011011001011101010110100100110101000;
#1 $display("%b", po);
# 1  pi=207'b001111001000011111010110011111001010100111001001000111011110101010010011011100001111010111100100000110111000011111110100101000111101110110001110100111011001110100100010010011110100000101111000110100100110111;
#1 $display("%b", po);
# 1  pi=207'b001011100111111000000011110011110010100101010110001111000000010011100001111110011000000000010111100110011011001101101111001000100000010100101100111001110011110000100001100100100011001000100001100010110011000;
#1 $display("%b", po);
# 1  pi=207'b011110000011100110000101110010101001100111010101001101101101110001011100111101000011001100111010111111011100110101110111000111110101100000010001011110100110011011001101000100000110011010100111011110011001101;
#1 $display("%b", po);
# 1  pi=207'b101001011000110011000100100101100110011000111011000100111011001111111111011011100011101110111110001000001000001010111100101101011011001100011001001110001011011010010000001000001001110110000100110111100011001;
#1 $display("%b", po);
# 1  pi=207'b001101001110100111101011101110001100011100110000101110001001100001010010011001001000001111101111100100110001111011101011011010100011101101010100100101011100011101010110111001010110111111100101000100011000010;
#1 $display("%b", po);
# 1  pi=207'b000111100110010111001010010000001001000110000011011000110001011010100011001011011110001010011011100101001010011101111011100111001011001110111010001000100011101001111100000110101000001000110001101111110100101;
#1 $display("%b", po);
# 1  pi=207'b011000001001110000100010110111001000001100100000000010100100100111010100011111101000001001010100100111110001101100000000010001001111101001010001011101110001110101101000011100011000000100110111111100101010111;
#1 $display("%b", po);
# 1  pi=207'b001000111001100000000111000011100100110100001010000100001111100110100000011100001001011110001001011011001101000000110110000101010010011001000001110000110111100001101010000101110001101101111011000100110110111;
#1 $display("%b", po);
# 1  pi=207'b111111101011011110011000011100011001001101011011101001100010010010101111011000000000101100111001111100011010010110100110010110111000001011101000000111101001000101111000111100000111110010101000100101011101100;
#1 $display("%b", po);
# 1  pi=207'b010101000111001001110110011111000101101010110000100011001100011011000010000001111110000010011111101111100001011101001101011010000011110011011001101001100110110101110001111000110010010001110111010010101001010;
#1 $display("%b", po);
# 1  pi=207'b010111100000111010010000110001010110000101001110001111011111001110110011101000111011101111010110100100001110111100110001000100111000001000110010001010110110011010111100101100111000111001000010010000110011101;
#1 $display("%b", po);
# 1  pi=207'b010011110010011111110011011010110001111110101111100000000100011110100101100000110001010100100110110101010111010000001111001100101010100001011101000110000010001011110101001101110011111000011101011001001100100;
#1 $display("%b", po);
# 1  pi=207'b001111011100100000001011000111101110110000101001000010100011110110001110111001001100000011100000101001101001101101111100110011011000111000110110110110100010100110000001110001001110011110110011001000110110011;
#1 $display("%b", po);
# 1  pi=207'b000110010000101100110010000010001010010000111001001000000100101100010011000110111101100011111001100001000010100110000100011011110111111001111101101101111111011000111100000001011000101100110001011111010100010;
#1 $display("%b", po);
# 1  pi=207'b011010110111110100011011111100000111111001000100011101010100101010100101110011000101100001100011100001010011001111110000001000001101010010000001110001100100110111011101000110111000111110000010100100110000001;
#1 $display("%b", po);
# 1  pi=207'b011111000000110010110010011111111000011001110001010011001000110100011100000010000101010100010100000010010101011011000111010000010101110110011011011000001111100011100011100010101100100010110000000011011010100;
#1 $display("%b", po);
# 1  pi=207'b111011110111111100001101010100110010000101011101101001010111111001001010000101100000110011110011001101110110100100010110011011110100010010011001101100111001000111010001011000001111000111011000010000100101100;
#1 $display("%b", po);
# 1  pi=207'b001111111110110111111011011011101011110011011100101001100011110011110110010001010000101111011110100100101111000011100111001111111001101100101100010110010101011010010111011000110000100101010001110011000010110;
#1 $display("%b", po);
# 1  pi=207'b010010000010101000100011111101010111111011000101100101111011010100011101001011011101101001111101000111110001101000011110010110000111011111110001101001101111111000011101001011101010111001011001110111001111111;
#1 $display("%b", po);
# 1  pi=207'b110000110011110100010010011100110010000001110011101110010010110011101110110100010110011110100101000010000100010001000110101010101111110011100101001111010100011110110001101000000000100001100100111111001111000;
#1 $display("%b", po);
# 1  pi=207'b010110010101000000101011000100000011001101000001000001110001010001111011010110101100000011111011111110000110100101010010101111111001101100111101111000100110010111111101011100010010001011111010000010110110000;
#1 $display("%b", po);
# 1  pi=207'b101010011111001111001110101000010000011011111001100001001000111100101101001111101011001010100101001110010110011001011001111001001001001000110100110010111001010010001100001100111111101011011000111101101111110;
#1 $display("%b", po);
# 1  pi=207'b101111111011001011011010011101100000100111001011000110000100001011011010101111001011110000111000001111101010101000010101100100011101011101001100100111010000000100110010010010001011010111100011110001000001000;
#1 $display("%b", po);
# 1  pi=207'b110100001011100010111010000110100100001011011100010111011010010110101110001100101001011000100000110111011110001101111010111110100001011111111000111010110011110100100010000110000001110101001011011010011111101;
#1 $display("%b", po);
# 1  pi=207'b001100010100111110011101001110001110011100110110010011011010000110111101010011100000100100000101010011001101101110111100110001110011000111010101111111001000100011001010111111010101110111010111010111011101001;
#1 $display("%b", po);
# 1  pi=207'b101101110101001000000110101100100011110010001001011101011110100010000011001000110010110000100010010101000001011001010010110110001000001001011110011101011100111100000000100001101111010001010101110010011101001;
#1 $display("%b", po);
# 1  pi=207'b010010110100010110011010100001100101001011111001000010010101101000000111110001111111101011100011100001100100010101011011010000101111100100110010101100001110001011100011011100100100111010011101011011100100011;
#1 $display("%b", po);
# 1  pi=207'b101110000101011101100010101011101001011011100111110110110101101111000000011101100001100010110111011000101011100110001101101100001011010111101001001110000111111101100000111010110100110000001111000110001011011;
#1 $display("%b", po);
# 1  pi=207'b001010111010010001100100110001011101111111101100001100111110100101001100111011001111110001100110011110101100010000000100111101011001111111001001101010110101111110001110110100011000101111110110100001101000100;
#1 $display("%b", po);
# 1  pi=207'b110000011111101001110010000010100000010111010110111000010010010111011110111101101101001101011010010011001010000010110011011111001011101110010000011110110100011011100110101011111110110000101000101011010000011;
#1 $display("%b", po);
# 1  pi=207'b111110101110101001001110111101000100010111011011011110010101101011000011110100110100000100111101011000011000100010101101100011101100100100010111100000011000010011110110110100010110100111010011100100010010011;
#1 $display("%b", po);
# 1  pi=207'b010010101110000110000001111001001101101000100110100111010010001101011011010010010011001000101110000001000001101110100110101000110001100000010110011010100100000111110101111100000100110010011010000110100011110;
#1 $display("%b", po);
# 1  pi=207'b010010010011001000111110100001111000100101010110011010111001010011110111111001111111000111111101010000000110110100100011000111101010001101010010100110110101100010010110011011001011111001001100111011011110001;
#1 $display("%b", po);
# 1  pi=207'b100010100011100010111111110010011000010110010001011100001101000100111110101011011000011101101110001111110110001011101001010000001111010000110001110111000110101010000011101110010110110100010010111001101110000;
#1 $display("%b", po);
# 1  pi=207'b110100001000101010111001000010000101010100000111111110011001010010101001000010011000011000000000111000100110101110010111101101000000000111111000010010001010000011101010010010101001010111000010011100110000101;
#1 $display("%b", po);
# 1  pi=207'b011101001011110001000101001100011100011001011000010111000101000110010010011001001000111000111010010111111101101101111101011000010000110111001110100000110010110000000010111010010111100001010111010001101111001;
#1 $display("%b", po);
# 1  pi=207'b111010000100001010110011100110110000110100000111001101110110001000010100110011111111001101110001110110100101001001001100100000101100011111001111100011011011000011100111000001111101000000110000001011101011001;
#1 $display("%b", po);
# 1  pi=207'b100100010001101110100000100011100001001110101011011010011000011111100011011000110000111001101000010101110001110110001001110011001110001001100001100111101011111110000101011011101110100100000011000101111100011;
#1 $display("%b", po);
# 1  pi=207'b100000101001011101011001011001100000100001000111000101001010010001000111000011001110111010001100011111001100010000001000001001010111110110101100000100001010101000011100101001011001000100100111010010101100110;
#1 $display("%b", po);
# 1  pi=207'b010001110011010110111011010001010111110010000100000110110001011110111110101110011000000001111010010101101100111010110010111111000000011111110111111011101010101111011100101011011011011111001000101110111111111;
#1 $display("%b", po);
# 1  pi=207'b000010011110010100011110010100100100111011111001000100001001101101010110111110110011001000100100011001111101001111110010010010110000100111011010010000010010101101100000010011001111001010000101001111100111111;
#1 $display("%b", po);
# 1  pi=207'b100110100100111101110000101010110101110110100101100000011011111101010010010100101111011111001111101010100011010010111101011110000101011100111010000101101000001110011000110100111001001011001100010000010011111;
#1 $display("%b", po);
# 1  pi=207'b101100010011110000101110110010100110001100011011001000110111001011011110111100111101101110100111000000100101010111011100010011100111011101111101011111101010100011100001111101100011100001010000101110011001100;
#1 $display("%b", po);
# 1  pi=207'b011111111110001011110010011010101111010100110011100111110011100010110110000101010110001100110011111100010111110011011000011011010101001001001011001110100000111111001000110000011000110000100000000001001110000;
#1 $display("%b", po);
# 1  pi=207'b101100101011000110101011000001010111101011001011000101000011001100111110100100110001110110111100100111110000000010100001100000011001010100010111000011100010111101011100011011110101101010011001100001001111101;
#1 $display("%b", po);
# 1  pi=207'b000100111101110110001111101100000100110010110111101001100111011101110001100001010001111001011101011111101111101100101011111101001111100111100101100101101011000011101110010101111010001110101000001000111110111;
#1 $display("%b", po);
# 1  pi=207'b001010000011100011010011000011011011111000011000111000000100011100100111000000001110011111100100011010100101110100100010001000010011111111010111001001000110001101110100011011000000000111001101101011101100010;
#1 $display("%b", po);
# 1  pi=207'b000101111101010110011111111111111000101001100000111011110110100100101000100011001101011110000100111100100010101001001101101110001101100010111000000010111110110001000010000000011101100011000110001011101000010;
#1 $display("%b", po);
# 1  pi=207'b101010100100001001100011111010010000100101010011111111011011000101001010001000100111010001000001010000101100111101001001010101001010001000011000000100101001011110111001110000001011101001010000010011101010000;
#1 $display("%b", po);
# 1  pi=207'b110010000110101101100001010010011010101110101101001010100100110011000010010010110110010010101010010111001010100100111101001101111100010110100011111110011101110110110011110101000111101011101011011010101110001;
#1 $display("%b", po);
# 1  pi=207'b001010010101110110011111111101000010100110000101010010101010101010101100101110101111001010111001101001101010010101100010011010011110111111111110111001110010000110011000101111110101010011100100101110111011000;
#1 $display("%b", po);
# 1  pi=207'b001011001011111100101111110111000011101100001001010100011011011011110011010010000001111011010001011100111110100110010011001010011101001101001111011001110011101110101101111010111101001100011011001000111001100;
#1 $display("%b", po);
# 1  pi=207'b101111101101100111000000110011100010010110110101001011100000100001111111111011110111111000110111001001011011000011010101011010100001111010111000111011111111010010110110011101111100101111011000001001001000111;
#1 $display("%b", po);
# 1  pi=207'b111101100100100011111000100111110101010111001011010000111101101001010010000001110011000000010011111010000101100011011011100111100110101100000111110011111111100010001011101110100101000000011000110101001100111;
#1 $display("%b", po);
# 1  pi=207'b110100010000000001110110000010101010010111100000000100110111011100101000010001100000011101110011001000010011011101100010101011101110100100001110001001001110110001010000010010100011011000000011111110000000101;
#1 $display("%b", po);
# 1  pi=207'b100100100110110100011010100101011100011000010011101111101010101010011101101011100100101010101101010101011011100100101010001001000111111111010010010010000101100010010110111110000010110110010001011011101001010;
#1 $display("%b", po);
# 1  pi=207'b001010010110000101101010000001110100010111001000010101110110111101100011011111000010110011101001100100101001100001100001111000101001001010111011100001000000101011010001001110100101111011111101001110101110010;
#1 $display("%b", po);
# 1  pi=207'b111110111001010101110110110110110100011110110010011100000101011111110111110111111000000101101101000001011110001001000100110011111110101101110000000000000011001011111011110110010010110000101110001100110010001;
#1 $display("%b", po);
# 1  pi=207'b011100000101011010000100010010110101010101101001011111101010101001110110110101010000100101111010111101010001101000110001001101001010100011111101110000100010111100010010101000010110000111100001011111000001001;
#1 $display("%b", po);
# 1  pi=207'b000010101101111010001010010010101001111110011000110100001111110111110010100010101100111000010100001100111101001100010111000001010100000010100100001100100000000011011110011010101000001001110101110111000110111;
#1 $display("%b", po);
# 1  pi=207'b101010011101011111110111100000100101100100100011110101010100110110110111110101010100110100001110010101100011001100111110101101011110101000101001010100011010110110011111001110000110111001100100100011110000000;
#1 $display("%b", po);
# 1  pi=207'b110111100001001111111001011101100011100010011110100010001000001100100111000001111010001101001001001001100111010110000011011010110001010111111100011011100101010111110010000010101110110110111001110001111001110;
#1 $display("%b", po);
# 1  pi=207'b100111011111001101000110111101111010101011100101110010110101001001111110110111000100001100010100110000011010100001111011100110111100001010011001000010111000011011001110010101001111111011110000111110100010000;
#1 $display("%b", po);
# 1  pi=207'b111110110111111110001111100010111010110000011111111000000000010100000101000100010001010010100111111110001111100111110101100010110100110100101011001110101001110100100001011001001010001011011101011100111100011;
#1 $display("%b", po);
# 1  pi=207'b010001000000100110100101001101111001000011111001110111110100011101100010111101010101000011101100001100011100101100110100010100110111111001111101010101010100110010010011010010011101001010011000110001000100001;
#1 $display("%b", po);
# 1  pi=207'b100010110100010000100000100000000000110000010101010010001101100101010101001001101110000100000110111101000011101110001100000011000001011110011000000010011000011010100001100000110000110111010110101101111110100;
#1 $display("%b", po);
# 1  pi=207'b010111101111001111001101110111111111001000111001010101110100001101101000000110111101110000111100001110111011000011110101111011010110001000110000000110010001111010010110010011011010110010011001011011010100110;
#1 $display("%b", po);
# 1  pi=207'b011100101101010001000000110010100110001101000111011100101011000000110110000111011000000000011011010100010100110010111010011111110101000101011101011000111001011001010000001001001101100010010111001000000111010;
#1 $display("%b", po);
# 1  pi=207'b010010111010011010011010110111000100111101010011010000111010110100100110011000000100111100110011001000011111100000011010000000000101011110110101010100001101101100100011000001100001111000110101101111111010001;
#1 $display("%b", po);
# 1  pi=207'b001010010110111011001011101001000010111101001110001100010000011011101000001101000111010000100110100100011100000110010111110101001100111011000111010110110111110000101101011000011001001010010011100000101101101;
#1 $display("%b", po);
# 1  pi=207'b111011011001100111101101010101111100101110001110110101110101101110110011101101110100110100100001010101110111110001000111000000001011001111111100010101100011111110011000101001010001000110001000010010010101110;
#1 $display("%b", po);
# 1  pi=207'b111100001101111100101010110101111001111011011010001100000110000100010111010111001110001101100101101001010111100011001000000110111111001111100011111011011001000001100010101111010111010010100000000011001000101;
#1 $display("%b", po);
# 1  pi=207'b110010100000101001101111111000100111000000000111010110010111110000001101010101110100010100110101101111101110101001010000110101011011111100000011111000000100011001010011010010110110001110100010110001011011111;
#1 $display("%b", po);
# 1  pi=207'b000010111001111000100011100111010100011001110111011110100100001111010010001111101010101100001000100110101011110011011101101111000101100000000010101111101110110001100111101111011100000000111001011011001111011;
#1 $display("%b", po);
# 1  pi=207'b001110011100111110110101011010010010010110001111110011011011100111001100101101110101101001010111000110101000001100110101001110110010110101100010011010011101000110101000111011101111000010001001111011000000010;
#1 $display("%b", po);
# 1  pi=207'b001001100100000001011101001101000010101110100110101110111001010111111100010110011111001001110101000000110111010111101110011011111110010110110000000010010101100111000011111011011100111011111100101110001001111;
#1 $display("%b", po);
# 1  pi=207'b110001000110000011110010101101010011111001110100100110011010000000111101000101111101110011110111111100000000001011101101010000011001001110000110011010111111010010001110010010110010101111100101111111011011010;
#1 $display("%b", po);
# 1  pi=207'b000111010101000001110010110011101010001001111100111110111000111000011001001101010010010110010011000111000110110110010110100100011011001000101101101111000000100011010010000101110000011001000110001111010001101;
#1 $display("%b", po);
# 1  pi=207'b111100011011010100110001010001001001011000101111111011011101010010010111110001100000100100010101010011000100001110110100101101110010111011110101110110111011000101111111011001111010101011000101110000101000101;
#1 $display("%b", po);
# 1  pi=207'b010011010000100101101110000100001110001001001010111101011111110101011001011101110101101100101101001011001011101011010010000111100110001111001001100000111011101001010000101100111000000001100110010000001001011;
#1 $display("%b", po);
# 1  pi=207'b111010100000010000101001000000101101101001000011010110111110111100111100010000111111011110001010010111010111001010011011000100011000100101010110100111000000011011010001110100010101111010000101101100010000111;
#1 $display("%b", po);
# 1  pi=207'b001110000011010001011001010100100000001000011000011011110010101010101100101101101001001000000101110100100010101001111001111100000011101100001010011010001011111010100110101010101111001111110100100011010011111;
#1 $display("%b", po);
# 1  pi=207'b001101101100010100100101111000011101011011011011101000010100001000010011110001010000010101010001110100010110010000010100101000110010111111110001100101010101000010011000011100111011111110101110010000010100001;
#1 $display("%b", po);
# 1  pi=207'b001010110100111011001011110110100101111010011100101000111001010100110101011000000010111110111101000001001001000010110111100100100111110010101110000001011011111001010011100010001000110111101100101010011000000;
#1 $display("%b", po);
# 1  pi=207'b011001000010111011011101100011011010110011100010100111101110011101101101110001000110011010010100001100011110101100000000001011001111101001101001010110100110011011111000110000110100100001110111000011001011000;
#1 $display("%b", po);
# 1  pi=207'b001011101101001101110010010101111110011000001110110110001100101011110100011011111000111110010000000000100111111010111101101101011100001100111100110001100111000000100100101101110011001011001010110001100100001;
#1 $display("%b", po);
# 1  pi=207'b110010111100001011101010001001101011000011011111110101001010001100111111001101000000011001011000110010101111101100110100011001000100001100100001110110111000011100010010100011111010000001010100010001101011010;
#1 $display("%b", po);
# 1  pi=207'b010000111101111110010110100110001001010000111110111010110101110010010111111001000000110101101011000000101110001001001110101010100000010000010101000001011101000101111001111011111001100000101111001010111011101;
#1 $display("%b", po);
# 1  pi=207'b001111011110101001001011111000110111000110001101110101010001111100000100101100011100111110001110101001110000111000011110111110011100101101100000001010110010000100000000101000001000100011001101010101101010101;
#1 $display("%b", po);
# 1  pi=207'b100110101000010001000001011111101101111001110010011011111111010111011000011011000111010110101011100101001101100111111001111001011111110101110111011010001101001010000001111011000011001110111010100110100000000;
#1 $display("%b", po);
# 1  pi=207'b010010100001110100001110110010110011100110011101001000010011110010111100110001100011100000110000001000010110111001000101100101100111101000100011100010101010001000101010001010101001111111011100010100100100100;
#1 $display("%b", po);
# 1  pi=207'b001101000010110100111000010110110010100001001001111011101001101011111111111110001011101110110010010001010001011000110111010100100010011001001010100100010010100100000010010001000110100111011011100110111100011;
#1 $display("%b", po);
# 1  pi=207'b100000011010000101000010111101001011000001110100100110100010111100000010100111100011000010001000111110111000011001110110000001010111011000101010110110100010011010000110111101110111110111001100011101100101111;
#1 $display("%b", po);
# 1  pi=207'b110100101000011110010010110000101010111101111010001001011111000001111101010101101000110001111011111111100000001001000000011111101011011110111010110110011110001100111010000100111011001101001110001110010100101;
#1 $display("%b", po);
# 1  pi=207'b011100011101110101010010011010001000101000110010110110100110101010110110000000001010011010001010111010011111000001110110010010001110010001000101010111110101011100111110111001100000101000111010111110110100011;
#1 $display("%b", po);
# 1  pi=207'b110111011110000010111110100111000000110111011001010100010010011000101011011101101101010101100001100000000000100011111110100100010001001101100111111011110100101000001011000111011101111001100111111000000111010;
#1 $display("%b", po);
# 1  pi=207'b100111000100111010001001100101010111111011111101110011100011110100100100000101011011110110011010010101010110100100011101101010111011110010100000110111001111010100111111100000011110100001100011101001111011111;
#1 $display("%b", po);
# 1  pi=207'b101111100001011010100110100101100110010001011111110000100110100110100010110000001001010000110100001001101110011001100011101111010001110010011011010000101110100000100000110100110000000010110001001001101101101;
#1 $display("%b", po);
# 1  pi=207'b111111011111011111100100100111011110111011000001001110010100010111111101001111100100000100001001100010110100000110001010001111110111011100110111000000000111000100110011000100011001011111000011111110001000111;
#1 $display("%b", po);
# 1  pi=207'b010111011001001101111111001110000100110111100001000000001101000000100111111110100101111100001010010011111100101001111011111100100110000011000011000010101000111101001111100011001000000000111011001100011101110;
#1 $display("%b", po);
# 1  pi=207'b111101110010001011001011000111100000111101110111011010000001110010111001010101101010010000001011001100101101110000000000000000001101000101011011111101010011110100011010010111101001000100100101101100001110111;
#1 $display("%b", po);
# 1  pi=207'b000110010010100010001000001011001011000001011101100000011011000010000100000110000011001101111010001100010000011101100111100001100010111000110011010101001000010010110100100011101100101001000000000100001000000;
#1 $display("%b", po);
# 1  pi=207'b101101100100111101110010100001110100111110001110101101100111111000000110111011101001100000000000101010110011100100111111011001011110000010110100001100110111101101011010001100001100010000110001101000101101111;
#1 $display("%b", po);
# 1  pi=207'b111100011010011001111110111000110101000011010101100001111110001110010010110110001100010010001101111000111100110101100100111101011101110000000111001101110101110001111000011110101001010101110100001110111011101;
#1 $display("%b", po);
# 1  pi=207'b110100101011100101000111111110111010111011001100111000010011010011010010101000010011010001010111001101010101111010100011101111110001001101101101101001011110110100101111010110010000111000011010101010100000000;
#1 $display("%b", po);
# 1  pi=207'b101110011001101000110100101110111111100110000101101111011101101110100000000101110001110101101100100011011001111110000110111101010111010011011100101001000011000011001101001101110000010101100010010101001110100;
#1 $display("%b", po);
# 1  pi=207'b101010011100101001111101101001000111011001110111011011101100011100111100110011010001101100001010101010110011011000111011110010100101110111111011001101001010111001111010011010111100111010000110100101010001001;
#1 $display("%b", po);
# 1  pi=207'b001101010101101001000101001101000001110001101100110000000001000001000101110011010111100110110101000011001110110110101111000110010101001010101001110010011111000001101011000111011111111100000000111111010111000;
#1 $display("%b", po);
# 1  pi=207'b101100100000100111000100101001000101011100101010010110101010110001101010110111111111111011100000000110111101001011010000001111110011100000110100000100101111001000100011010000010001100101111101010011000100100;
#1 $display("%b", po);
# 1  pi=207'b010001011101011110011010111100010000100111011101001011101100100101011000100111110010111100111010111010010110010001000100001101000111011011111011000010001110101101000011111000011000001100100101101111110101001;
#1 $display("%b", po);
# 1  pi=207'b100011110111100100011000110110000100111001111000000110101100001101111001001100010000100000001101110010011001000000010000010100101110000110111110100111010001101101001000011101111100010110101110101101000000000;
#1 $display("%b", po);
# 1  pi=207'b111010011101111010111100011000101110001010011001010100100100001101000010000111011100101011101001100100101101100101011111000000110110101110110011010110011010100001111100000111111011011000010000000101001100010;
#1 $display("%b", po);
# 1  pi=207'b000100100100011011111010101000001110110000100110011001010001001001011101011011111010101010000100010110110011000110110110111110000111001110010110100101000100011100101000010001101111111101100011010100110000100;
#1 $display("%b", po);
# 1  pi=207'b111111011101000101111110110010110101101101011010010101100011101001000001100001111110001101010111011000010101010100001010111111010010011110110011100000111011100001110000100110101110111100101001101011001011001;
#1 $display("%b", po);
# 1  pi=207'b111100100010010011011010000111011001011101000100110011110101000110000010100111100111100010000000001010001000011010011010110010011101010010111111100011011001100001000110000000111101001101110111111101011011100;
#1 $display("%b", po);
# 1  pi=207'b100100101011011101001100100110000101111110000101110110001110001000110001111001001000000000110000010111010110011011011010111111111110011010101001001011110100111010101010010011001011101101101110000110010110100;
#1 $display("%b", po);
# 1  pi=207'b111011101011101100010111001010011111011111000011011011010111111000000111010001000000011000111110111111010110001110000101100101001100100011100000000010100110100111010110011011110010101011100010110101010111110;
#1 $display("%b", po);
# 1  pi=207'b001001101111110110111101100011000000010111101110000010100010010101011100110011010110000101111000101001101100110101111111111111010111101010101100010001001011101100101111110000000010100001111010001001100011111;
#1 $display("%b", po);
# 1  pi=207'b000100100000100110100010001100000110111011111010101100111001001110111110101110110000100111000101101101001110100000111101010000111011101100110000011010100011110110111110100000101101101111111000000011010100001;
#1 $display("%b", po);
# 1  pi=207'b110101000111100010001011101011010011011000011111111010101010110100000001101101001100000111101111000100110111110100110111111011000011010111100101100111100010110011001001000101100001111111100011101011000100011;
#1 $display("%b", po);
# 1  pi=207'b010100101100001000010011101001100000100101010011010100110101100010001111000111010000000011101011000010110111110010111101110101101100001111010110100101000110101110011110110110111111000101111001000001100110110;
#1 $display("%b", po);
# 1  pi=207'b010100101100000001100010010110111000101110101101111110010001001101001101011111001000000000100101000010101100111101000100011010011101110111111011010001110110100001010001110010001101000011000000010100110011010;
#1 $display("%b", po);
# 1  pi=207'b011000110011111100110011111111010111111101111111100010111101010111100110001010001101010101010011111101110010010110011111110110001111010001111011000000111010000110011001000111110100101101001000000101010000110;
#1 $display("%b", po);
# 1  pi=207'b010110000101001111101111000011010000010001001011010001010101111110011101100000001100010110000110000110111011011110001000100111100101110100111101101010011111001101011001101100101010001001111110100010000101110;
#1 $display("%b", po);
# 1  pi=207'b100100011010000011110011011110001101111100111011001100001110000100000010000110110001011110111110101111111111001101111000101100110111011011011011000001111010010101110010100010111110001000010011110010101000001;
#1 $display("%b", po);
# 1  pi=207'b010111000011000101011101101001110101101100110000101100101010011110100111100001001100110111000100011011011101110000000111101100110010110001110100001111000001101101101110111000101100110101011100001010000011101;
#1 $display("%b", po);
# 1  pi=207'b010110110101101101101001111111011101110101100110100011000010001111111101100010010111101110111010010010001011011110110100000110111110011011001111100100001011110001100000111010011011111110001111110011000000101;
#1 $display("%b", po);
# 1  pi=207'b110110010011000011100001101010101011100000011001101100010101011100101111001110111111011011101101010100100101010110111110010010110100110111110011011110100110100011110111000111100010111011100010001011101001111;
#1 $display("%b", po);
# 1  pi=207'b000001011001001000110111110001000001110001011010101011001001001111111010100010100010000110101000111000101111001010010101101011101010011000111110110110110101111100100000001111001100001010110101011111001001010;
#1 $display("%b", po);
# 1  pi=207'b010010011001001011101111000010010100100100001000110100100111101110001111100001010101110101110001110111001011100010010100101101111101101100110011011010110101011110111110110011100111100001001010100100101001011;
#1 $display("%b", po);
# 1  pi=207'b110011011001010111110110010001100110010101000100011101010000000111101100000001111111010001000000010011010001101000001111101111010100110010100110010101100111101111101100011010011010100000011011010000101000100;
#1 $display("%b", po);
# 1  pi=207'b111100010011001011011100100011000010011000100011000110001010100101111101000111111011011001000111100111100100100001011010001100001101011011011001000110001100000010100111000111110110101000100110100101010100110;
#1 $display("%b", po);
# 1  pi=207'b110111000110011000000001100000101011001110010001010001100001001110001000101111001000101101000001101001100101110011000100100111111101101111110110010111100000100110011110110010100000001001011100010001100001010;
#1 $display("%b", po);
# 1  pi=207'b100110001101100001101000010110000000101101111001111000101000011111000001101110101001110011100110100001011111011101001101011110101001100010011101111001010011000101010110001000011001110111011011001010001011110;
#1 $display("%b", po);
# 1  pi=207'b011101010010101100000010011011011100011011010011001001000011100100001101001010011111000111111001001101110100101010101011000110001100001111010010001010001110011110011100001001111001100111011001001111010101000;
#1 $display("%b", po);
# 1  pi=207'b001011000010000000110110110101100011100000110000100010011000101011111000100010100101100011101110010100100111111110110110100010010100010110001100000010010001010100100010000101110011111011110010010111101111011;
#1 $display("%b", po);
# 1  pi=207'b100111000010100010010011100110001001100110101000010100100101111001000010101001011001101100001111110101101110011111010111101101100100101001001001111100011111011010001010111111010010111000101010001001110000000;
#1 $display("%b", po);
# 1  pi=207'b101100111000000100010101101110000100110101000110111000011011000100110001001101001111011101111101111011010101111101100111100011100000110110101110011010000101000101010111110110010001010001100101111001100110100;
#1 $display("%b", po);
# 1  pi=207'b110011000011011110011110100111110011011110101001101011010011100001100111011101010000111110001110100001110101011011011101011110001111010011001000111111010011110000011101001100000110101110000000111011011010100;
#1 $display("%b", po);
# 1  pi=207'b001010011000000011111100101001010011110000001011001000001000111100011110101111100101000001000101010101111011101100000101110110010010111111101001000111110010001111010000110111000101110111100001100111101101101;
#1 $display("%b", po);
# 1  pi=207'b110001101100101011100010010111001011100101001101100111110010011111101001100000010101001000111001111100100011111100111110000111101011101010001100101001100111100101011110011001010111010010000010111110011001100;
#1 $display("%b", po);
# 1  pi=207'b001100001101001011101110101101011100110011000011100000001111110010010101110110001111110011011010111100011000111101011010011011001101001110011000011001011011100011000100011001011001001110110011111010011100100;
#1 $display("%b", po);
# 1  pi=207'b000011011110100011001010000000001110011111001100111101010010000101111001110100111111111010010011101001111010010110010011101011011110110000010101001100011001111100011011001011010100111100110110011101111100110;
#1 $display("%b", po);
# 1  pi=207'b000110011110110100010100001101111110110011011101110100100100000010111110101000101011000010100010101101100010110110000000000110001101001101111001011011110000110101100001010101110011010010101011101001010011001;
#1 $display("%b", po);
# 1  pi=207'b000001001111011100100100011011100010000001111111000110001001001010101101010110010001100011101100100001100100101011110111101100000100111010101101000001001110010010010110111110110111001000111101100101001001010;
#1 $display("%b", po);
# 1  pi=207'b011111010100101111110011110011100011001011000010011111111111000100000111000111101011000000100111100011001110110010111000110001001110011001111111111111111111010000000001011101110011111010101010011111000011100;
#1 $display("%b", po);
# 1  pi=207'b001111100111101001001011101001100110111001100100011110100110010101110110010101010100000101000001110100111110011111110101111110001100110100010001010010010000011001111011100010111011001110101001011101010001110;
#1 $display("%b", po);
# 1  pi=207'b000101110111001001100111110001001000001010100101011001001011101101111000111010001101111111110000011100010000010110001101001011000110001111101111101000001110100110001111111110101010100000101000101011000110100;
#1 $display("%b", po);
# 1  pi=207'b000001001100111110011100110011000000011001011110010010000001101111010010101111001010111100101100001000011100100010001100110001111111111100010010011101101100100101110001000101001001000111000010100000010011100;
#1 $display("%b", po);
# 1  pi=207'b010101000101111110100101111111101100100010010111101001101001111110101011001010000001101011000110000111110110011001001000110011010001011100000111011001111110101111010011111000010110100010001110000101011100011;
#1 $display("%b", po);
# 1  pi=207'b110110000101001010011101010101000011000110010001001001101111110111010010011110111101110011101110100001001000000001110101101000001110000110111010111100110011010110001110110111000110011111110011001010010011001;
#1 $display("%b", po);
# 1  pi=207'b010111101101011110001110110011001011011000100100010110100000011100010010110010000111000011100111000010010111111111101110010101000101110011101111101010010110010100101100101011101011101110100010000111011001110;
#1 $display("%b", po);
# 1  pi=207'b100010100010110100000100010001000100000101011110000100001111110000000100111000011000001110110000110101110000101010011110100101101000111110011000011111111111100111100000001011001011100110110111111000100010001;
#1 $display("%b", po);
# 1  pi=207'b000111111110010000000011110011001110000010111000110100011010011010011101100111101111110100001011110101100110011010001000000110011010010000010011000101010001011101110110001011101010011010011100010010011110100;
#1 $display("%b", po);
# 1  pi=207'b110000001101001101101000011101110001010100100001111010001101110101110011010110011110000011100110110100010000111000110000100001011111110010010010101100010000010110111110101111111001111010010101100001101000000;
#1 $display("%b", po);
# 1  pi=207'b100000001111101001101110110001010001111111101001110100001110001101110101001000011010000011000000000001101010111001001010101000001001101011011101011100010000001000001110111100001111001010010001011011011010100;
#1 $display("%b", po);
# 1  pi=207'b010010110011101101001111100000011101110110011001111000101001000111011010111110001001100011111110010110101110000011110010000010100101010010101111001110010011011110011011101110110000111110110001001000101111000;
#1 $display("%b", po);
# 1  pi=207'b000001110001110010101101000000011011010110011101000000100101010110110001101111010000000101011110100111001100011101010111001110111001100111000110101011111111100001010110101100100111111111001001010100011011100;
#1 $display("%b", po);
# 1  pi=207'b101111001110111110001001010101001100010011111000100110000001011100010010010010100110111111001010111000000000001011110100011110111111111001000101110110011001000011011010111010001010011010010010010101101101011;
#1 $display("%b", po);
# 1  pi=207'b101111011100010111111100000010100011110000000011000110000000101100010110011101101101010100101101010101001001010001110110100110100010101101111110100110010001000011100100000111101101100110010111000001110100001;
#1 $display("%b", po);
# 1  pi=207'b111110011100101001010001010111001100001111100101100110001010000000101100100101001110010101111111101110101011011111110100101010100011010010110000001100101001010111110000101001111000100110010100111110010000010;
#1 $display("%b", po);
# 1  pi=207'b110101000110110001101000110011011111110001110000011000100010111111101101100010011110011001100011101001000011111011100010000101111100101101000111111101110110101010111000111100100100010010001101100010001011100;
#1 $display("%b", po);
# 1  pi=207'b001110000000011011011011101000011110101100000011011110110100101110001100011111100000111111101010001101000111001010011001110111110100001100110100110101011001111111000000000000000110001100100000010011010010111;
#1 $display("%b", po);
# 1  pi=207'b010100010001010011100010100100000010111010100011100011101011100101101101111010010001000001111111110000001011001101101001100111010001110010100001100011110011110000001100100001111110100000111000001010001010101;
#1 $display("%b", po);
# 1  pi=207'b011010100111001111111000000000001000010111000001000100100100001011011010100110101010111001010010001000001011111011100000100001001111001111110000111100010010001100101101111111010111011011011011101001010111001;
#1 $display("%b", po);
# 1  pi=207'b110001001100010111110110011101001110111100001100011010110011110111010001100101110111001010110011110011011011110111001011011101101010011111110100111010011100011101001111000000010000000101100011010100000111001;
#1 $display("%b", po);
# 1  pi=207'b111111010011100010110110011101011101001100100000101100110010010111100111111010110010010101111111001000110110010011011011001000111101000010100101100100101001010010001001111110111111001100001011101111110110011;
#1 $display("%b", po);
# 1  pi=207'b011101000111011001101100001101100000100000111011001100011111101101010000110110001001011111001000101101101011110001110000101100100111000110100110110001100101101011110001001100001011100010101111110011111011001;
#1 $display("%b", po);
# 1  pi=207'b111000110101110011100000101101111100011011100101110000101101010000100010001010010110110101110111010110101111001001100100001110110111111010110010011001100010001100010001111100000001100001010100101001111101101;
#1 $display("%b", po);
# 1  pi=207'b111100100001011000010111110011111101101001111000000100111100101101010100110000110110000100111010010100001101000100010110100000010100100011001000001010100010101101010100100010001011110010000100001000100011101;
#1 $display("%b", po);
# 1  pi=207'b001110100100001010100010101110001101011011101110100000011011101000000110010000101101001000100100010001110011010010101011100011010111010011001110001101110011101100111111101001100101001100111111011111010001101;
#1 $display("%b", po);
# 1  pi=207'b011000001100011110011110100111010000101001010011001100110010101110010011100100010000001101100101111110001101001001111100110100010011010110100010111111110011101000011001000001001011010000010011000000111110101;
#1 $display("%b", po);
# 1  pi=207'b001011001000111001100101100101111100011100101101100101111110011101101101100010001101111000100001111110110011101111110111011101100001011011001011001100001010001000000001111101011010101111011110000101111011011;
#1 $display("%b", po);
# 1  pi=207'b111010010100101000101110000010100001001100101010000000101011100100111101000100000011101010010000111110100001001110001110101000110100001110010001011010100111011001001011011000100001101011001100100110100010010;
#1 $display("%b", po);
# 1  pi=207'b101110000100000001110010001000100001101101010000000000000011100010101010110100000101010011110100110010111000101111001000001011001010010001111110000111100001100010001001111000000001000011010111010000001000110;
#1 $display("%b", po);
# 1  pi=207'b101011001011001101100000111101100001110001010000111101100110100010000111101100111001011011011011100111001111001101001011101000110111111111100011010011011101100010111010101100011001001111000010011000000011110;
#1 $display("%b", po);
# 1  pi=207'b101101010000110000100101110010101111001011100001011101000001100010010100001111000010000011110001100101110001110001111000101100101011001000010011001100100100101010011110001011001000010111000101010111110111111;
#1 $display("%b", po);
# 1  pi=207'b010011100110100111010001010001110000111001101111010010000100001101010001111100110011101001000110001100111010101000100010010110011100101110011001101110111110110110001111001010011100110011101000000011101000000;
#1 $display("%b", po);
# 1  pi=207'b111111010101001111011111100001001110010110101011111110001100100010001101110011111001010100101010001111110001010000100101101001010110010001110100111100000010000111111100001010001101110010000001100111011100110;
#1 $display("%b", po);
# 1  pi=207'b011000101111011011001100111011110111111011010000101111000011010110010011000000100011000101101011111000111001100100001101000110011100000110111110100010110101110110000001111011110010011100101011001100100110111;
#1 $display("%b", po);
# 1  pi=207'b101010100111111110000111010100000101101000101000010101010000011000111111011101111000111010010101000001010010100100111101100110111001000100011101110010101011001011000000111100011010110100001011110110100000100;
#1 $display("%b", po);
# 1  pi=207'b111011101111100110101101110101001111001001110101010010101100110010001100100110110001000110000101100111011001011011111110111010000101111000000101001011111000010011110100110100001011001001110000110000101101111;
#1 $display("%b", po);
# 1  pi=207'b001100010110001101110110111110000111000011001011010100001011101001110101110110101100010100111001101110101100100110100100111111101101011101111110100111000101001010011100100100001110110011001111110010100011111;
#1 $display("%b", po);
# 1  pi=207'b100000110111101011100010100010011000111101011100110100110010010110111101001100101111111101101011010100011111101010100011100001101010000100011101001111011100001000011101111011010011010000101000100100100000010;
#1 $display("%b", po);
# 1  pi=207'b001001001000100110011011010100100100011100001000010111100011010110001011001011011100000010001110010010100001100000010010010000111100111001010010011011100001111010100001001011110100010101101111000011011101000;
#1 $display("%b", po);
# 1  pi=207'b111110000101001111100100101011100111000111001011111000001010100111111100011011110000110111001010110010101001101101101100000010010010000011110001010001100111101000010000010111110001100111101010011010101101001;
#1 $display("%b", po);
# 1  pi=207'b000001100101010011010110001001111101011110010110011011011000001010110101100001111110100110101111001011100111101010000001010010111111111111001000000101100100111111111101011010100111001111001000111100001111010;
#1 $display("%b", po);
# 1  pi=207'b001001011001010110100100001011110010001110101000000000101100001010000000100001001111110011100111010011100010010000011101001001010010010100010100101100010111100110011001111000111101100110111001001111110011100;
#1 $display("%b", po);
# 1  pi=207'b100010110111100001001100000101011011010001111111010011100001111111001001010101100001100000101101011100010010000110010010000110011000100011100110100101001100100000101000100100001010010100110000100101011110001;
#1 $display("%b", po);
# 1  pi=207'b010100110111010001011000101100100011101000001011100111111001010100011000011110101001100010110110101100110100111111110001111101011011100010100111011001000010101011000001101001100000111110000000110001110101011;
#1 $display("%b", po);
# 1  pi=207'b110001101100010110000101010111110010111100111110001011110101100001111011110110011010101001110000111010000111010110111000011111111110101010011001111101000011000011110111011101111011001101100100101001000010101;
#1 $display("%b", po);
# 1  pi=207'b011101011011010110001100100000110000110000101000100001000111010000100110000010100110101010011101001010110101000110110111010100101101001101011000101011001011111110100110001110011010010111001010000100010001100;
#1 $display("%b", po);
# 1  pi=207'b001101000000111111000101001000110100100000010101101000100010100100110101100011000000111011011000100011111011101101100111010100111000011111110001001111110001010010110111010101011010111011100010010101000110110;
#1 $display("%b", po);
# 1  pi=207'b011100100001110101101100000101101111000011000100000001010111000000100001110110111110100000010100100100111011100000111010100101111001001101010001000010100111011000111000111110001110101011111111011101000100101;
#1 $display("%b", po);
# 1  pi=207'b111000011111010110110001110111011101010001001011000111011101010011101110011000001101100101000111001000100000111000110100111100100011110000100000100011100011111000100111100111011111010011101100111000010101000;
#1 $display("%b", po);
# 1  pi=207'b001110100101001101101000000011000101001010101000111010001100111111111011111101110100100001001110111001011010011100011011101100011010111100010111100000100010111000111001001110110010010111010111101100110111111;
#1 $display("%b", po);
# 1  pi=207'b000101111001101010011011010101001010001101101111010011100011100011010110110011011001010111110000010001011011011101011000100100110111111001011011100110010011110111100011011100101110001000100010011011101111101;
#1 $display("%b", po);
# 1  pi=207'b111010100110111111111011111110000101001000011100100011011011000100111001011111101100001010110110110100100000100000101100101111000000000001011000011001001010110101000111111101011100000111011100110100101010011;
#1 $display("%b", po);
# 1  pi=207'b111101101101011010010100101100001110100111101010011111100011001110011110111010110000011010001011100100000001011100000110011100101111001101011011111110101110010000100111101100010000001011010100111000101111010;
#1 $display("%b", po);
# 1  pi=207'b000010001110111011010001010001111011100111000010111101101011111111100111001001001100110100010010110101011100001011101110000111111000100011010111111110111110010110001111000000001111011100100101110001111101101;
#1 $display("%b", po);
# 1  pi=207'b110100110100100110000111111100101001111011010111010100110101110000100110001100111100110001001001110100100100111110100000100000110011000011011010110100110000000000000111101000001001000100001001001111010101110;
#1 $display("%b", po);
# 1  pi=207'b011100101110011010000001100010110110110110010011010011111111011000100010100100010010110110100010101010111001110111000011101010100100111110010011101000010010000000110001100110010100100001101111110001011000111;
#1 $display("%b", po);
# 1  pi=207'b110110010100110110010110011001010111010111110011010101000000001101110011101111101101110001101110010111000011000111010010010000010001110001000011101011010100000111100001101010100100010111000010111010010110100;
#1 $display("%b", po);
# 1  pi=207'b000001110101001010011101011010011011010110110010010100010010011101111011001000011010001101000010011110101110111011000101010110000100101111100000011010110100011011110100111110100010000110001001011001100011110;
#1 $display("%b", po);
# 1  pi=207'b010001000011110110010111001110011001010001110101011100010110110101101100001110001001111011111010000001010111000110010111010010110000111111000100010110011000110100101000000110110101001100111110000011001100100;
#1 $display("%b", po);
# 1  pi=207'b000100101001101111111101010101101100011010111110001011010011000100010101011011100001100110011110100110100111100011000100100111011101110001000011111101111101001110010010110001011000111110000101110110101000111;
#1 $display("%b", po);
# 1  pi=207'b000011100101100110001100001011111110111100111011100000110100100100010010101001101110110010001110111101101011111000000001110101101001111011101101100010100100111000010010111110000110110000011111111100011001000;
#1 $display("%b", po);
# 1  pi=207'b000010101000011111101101101000100011001011010000011100100011110111101011100111001110001010010001100000001001010001111111101011000100101110011010110011101101000100110010010011111011110100001111101100000011010;
#1 $display("%b", po);
# 1  pi=207'b001011101111110001000001110010100111000001101010100000101101011110110100000110001001000111011101011111100001010100100110000100010110010111001100000110111010101100000011000010110011000001101111101010111101101;
#1 $display("%b", po);
# 1  pi=207'b100001000010100011110100011111010110001011000110110110101001011101001000111101010011111001111000000100100101100111111110011110000110011000100001010000100111001100100101110111101010010010001110101001110100001;
#1 $display("%b", po);
# 1  pi=207'b011100010011111000111011001001010101101001010100001101010110111011010110010110100010110101110111110000010010101011000101001111000000011101011011010100101111010001101001010001110001011100101001100000011010101;
#1 $display("%b", po);
# 1  pi=207'b111011011011101110001100000000010110000110011011111101100100000011001001101100011101001001111100011111010011010101010101100110101010000010111101101001111111111101110111100111111100111000010000100001101101101;
#1 $display("%b", po);
# 1  pi=207'b110110001011110011000011110100111101011101010111100110010000100110110111010101000010000011001001101000101110101110101001110011111011010001101010000101000011011100111100010110001110011100010100001110111011100;
#1 $display("%b", po);
# 1  pi=207'b011011100001110010000111000100001101001001111001000001010111101001111111001000010001000110100110001010000100111101100101011011011101110011001100011111101000010111111001011100110111001011011010011011111001011;
#1 $display("%b", po);
# 1  pi=207'b011001011101001010110101000111010111100101111000111010011000011110010111011101011111101001011010001110110111001101011110100010011111001101101101000111110001110101000010110111001101110011000111000100101011100;
#1 $display("%b", po);
# 1  pi=207'b010111000101100101011001000011101111001101101110101101010110010001101111000010110111110000100000100011000011010110000111101001010111011110001111101101010110000001101110111100111010010010110001101111010110110;
#1 $display("%b", po);
# 1  pi=207'b010010010010001001100001010101100110001100110001001111011011000010001011011001110110111001110111010001100010011110011110110100100000011110101010111001101010110101010101100100110011100101000100000101000110000;
#1 $display("%b", po);
# 1  pi=207'b010111000011001010000011011011001000100011110101111010011000001011111111101100111011011111011010010011100010000100000101010010100010001011100111000001101001101100110111110110010010001111011111000000011111010;
#1 $display("%b", po);
# 1  pi=207'b010000100110011011100100000000101100001110011111100111101000101001000101111000011011011010111101000001101000011011101010000000011111101011101011010100110111000111011101010101000111101101001010011001001000110;
#1 $display("%b", po);
# 1  pi=207'b100010110001110000101001111101011011010011110010001010010000001001000100010010011011011010001111111010010110011110110010101001011011010011100111011010000001111111001100110000101001101111110010011111001110000;
#1 $display("%b", po);
# 1  pi=207'b111111011001010010101001111101001011101100011101100100011011000100110111000101001000110100000100110001100100010111100100000111100000111101101100010000010100101011111011001010111110101100001000111010101100100;
#1 $display("%b", po);
# 1  pi=207'b100100110110000011110001101000111011111011110011000000011111011111101100110110000001001010001011010100000011000101010101100011000000010101000010010010000111111111000100010010010001010100110001111111110010001;
#1 $display("%b", po);
# 1  pi=207'b000100010010001101111100110110000110101011010001100000100111101011011110010111100101110100011010001100010101101011110100110011000011010110111101000001101100111101101110001001000000011100101101000100100101101;
#1 $display("%b", po);
# 1  pi=207'b011101010010000100101010101100111011101111101110111100001011000100000011011011100100110101100100010000111010000000101000101000111010000101111000111100101000011101011001111010001110100011101110101000100100000;
#1 $display("%b", po);
# 1  pi=207'b000100101111110100111110010111000011110001010011001101111101111100100100011110010110011111010001101000101111110100100100000011001101001100110010000011110111101000000110101000000101110100000101101111111010110;
#1 $display("%b", po);
# 1  pi=207'b100100010100000101001100111011001010100100011000010110111100011010100010001100111011101011010010000111111001111101000111100100010011001100111000011101010000111010111111101001101010111100110011000101001100011;
#1 $display("%b", po);
# 1  pi=207'b011100100111100000101010001101010000001000100111110001011101110010010101000111110011110010111111011010110110010010101111101001101110000000001000100010110001001001100000101101110110011000111101111110011110000;
#1 $display("%b", po);
# 1  pi=207'b001101011011100000011100100000101001100101011000100010000111001100101001000000110110011011101010011100100001110101111111011001101000010111001111011001111111110111010010000010100101010110000010100101101101111;
#1 $display("%b", po);
# 1  pi=207'b111001110100111110110100100111101100111000101000010011010001110010101000011001100100010000010000111111010100001101010100110111011100010111011111011111011110100010010101010101101110000011101001101000101011010;
#1 $display("%b", po);
# 1  pi=207'b010111011010011100000010111000101110111110000000000101001100001001110001110010001010001101011000010100111101011110101010000101100001011000000100010100001101110001001010000100111001111011111110010010001110101;
#1 $display("%b", po);
# 1  pi=207'b010001000101101100101111111000110100111011110001101110100110011000001000000011011100000100100010000100101110100111110100101010000101101000001110101100010010111010111111001001101001101111111110100000101110100;
#1 $display("%b", po);
# 1  pi=207'b101110010110110110010100101001111101100110010111110001111101011100101010101011111111111000000000101101101010101010101111100010001010111011011011101000001010110111000011000000101100100110100001110001100010101;
#1 $display("%b", po);
# 1  pi=207'b010111011100000101100111010001011111101100100010000001100001111000000111101100011101010011100010011100000011001010011100110110111111010101101100010001011010101110111011101110111110010110000000110001101100001;
#1 $display("%b", po);
# 1  pi=207'b100100100111100101111000101000010111001101100010101101111010000110101001011111000100100110100100000110011001011101100001111011001001010111010111111111001110110100100010001100111001110000101011011100001010010;
#1 $display("%b", po);
# 1  pi=207'b101111000110001000101110101110101011101100101000011001011010100111110111001110110011110100000100110001000110100111111100011001000000111010010010110100111001001100000001110010001100011111010000010010110000111;
#1 $display("%b", po);
# 1  pi=207'b100001100100010100110110111100110010011111100001010101010100100000011011010010000110110000110111011001010101001010000100001011101111100001110100110011111011111111011110111100100010010010111000001111110111110;
#1 $display("%b", po);
# 1  pi=207'b110100000101001100101011111100011101011001111110110100100111111001001101110110111101110101100001100100011110100111001010100011010101010110001001100011001111011011100110110110010100011100000100110010111000110;
#1 $display("%b", po);
# 1  pi=207'b010100011110111011110111010010101000001000111000001111011011000010011000000111011001110110010000011101001001001101011100100011001000001100111101000100001110111110000011101111101011100010110010000010010100010;
#1 $display("%b", po);
# 1  pi=207'b101101001111111101001001111101011100101110000101000011010101100110111101111010001010000001011101001111000110011111100001010001110100011100010110110100001010111101010000110100000000110100110001100010110111010;
#1 $display("%b", po);
# 1  pi=207'b111010110111001100101111110001110110011101101101010101001011111000001100000011101011110100010011011011111011011010111101101111000110101101111110010101110110101010100111000011101110110110001001100001000110101;
#1 $display("%b", po);
# 1  pi=207'b111110110011110101100101001010011101000111010011100110111011000100110000100101000101101000111111101101010011110001101101011101101010101100001000011001000100111011101011100111000110110001001101111100111010010;
#1 $display("%b", po);
# 1  pi=207'b101011011100111000010111011101101001100011001111001011101001111010000011110101101010111001000100111101000011101111111000000100011010000001111001010000000001101100110101011011001011011000011101110001111011011;
#1 $display("%b", po);
# 1  pi=207'b011000100100111000001111011010101001001101110001000010101101101000011110000001110010101100010111100011010100001000010101011110101001011011100011000010111010101000011000011111001010010010100011001100110000100;
#1 $display("%b", po);
# 1  pi=207'b111000010100110111000101011111011000101110110110101001001110001000010011010110001011100010001110011110110111111100101111011101111111011001111110111110100000101010001101001011011100010001001101011011011100000;
#1 $display("%b", po);
# 1  pi=207'b111100011011001010110011010010111010110110111001000010011010111100010001110101010000010100010111100100111010111000011101010010110000000000100010010000011111111110011001011111001010111000101001001110001100010;
#1 $display("%b", po);
# 1  pi=207'b011110101010010101010000011111010010001000101100001110111110000100111100010110010011010010100000110111110100110110011010011000110010101000111001110000111010011111000011000100100111101011110111111011111011011;
#1 $display("%b", po);
# 1  pi=207'b000001100101101011011111111001000000011101011110001100011100100110101011110011101000100110010111100010101110110111100110010111000111000111110100000001111010011100010101000000000010101111001110110101011110110;
#1 $display("%b", po);
# 1  pi=207'b101111000101010110101010011011100000010110110010000111101111001111000010101111101100101001010110011000111100100011010011001110110010000001001000011000000111000110001001000110100111101101101000011010110000000;
#1 $display("%b", po);
# 1  pi=207'b100001110101111001101100110110010101001111101001110001101100010110100110101111100001111011100100010011011010011010101000110111101000011000110110101101101111000101001010001111100001001101010101111011001011001;
#1 $display("%b", po);
# 1  pi=207'b011101100011000010110001111001110010101100010101010000110001001001010101101101100101000100001011100011110110110010000101101001011101100011100101000110100111100000101101001011110000101101110011001001110001001;
#1 $display("%b", po);
# 1  pi=207'b100110100011100111100110000101001100011001111101011001110110110001010010101000110011100010101001000010101001000010111000101010101101100011110000111010000100111111011111111100100000010011101110100011000100100;
#1 $display("%b", po);
# 1  pi=207'b011001000001011000011001101010110110111000101010111000000110001111001101001000011011111010101101001010001010011011110100000100011101110000101111011001110100010011100110101011110111001000111001001101111001010;
#1 $display("%b", po);
# 1  pi=207'b101000010000010111011011010111000001000011100000010100101001100100001000110101011010101010010010000000100000101100111000100110100111100011110000111011111001001111010111010011011011001001000110011011111000110;
#1 $display("%b", po);
# 1  pi=207'b011010100110101011111100100000000101110110101100110000011110011111101011111101100001100001011001111111010100001001010110000100011011011111000100101010110110001010111101000001111011100010100010100100000001001;
#1 $display("%b", po);
# 1  pi=207'b100011000010111000001101010110111010100011001100010100010010010001001011011100000010101100101110010010000110111011111100111111110011110100100111110000001001001011010000110011000111000011010110011101111111100;
#1 $display("%b", po);
# 1  pi=207'b110010000000110111110110110111010011010010011011001110111011101011101111011111010110101000100111110110001110111111001010100001001110010000000111100101011111000101000101011001101000101101111110111011010111111;
#1 $display("%b", po);
# 1  pi=207'b001111010111011000111001001000001010001010111110011100011101110010011011010111101100111110010111101000111101110110010101000111100001110000011000000011011100011010000111100010100101110010000000000101101101100;
#1 $display("%b", po);
# 1  pi=207'b110100000101010110101001010100010111100100001010011101000100111100011000100110100110101101111110000000010010000100011000000110010110010001100000011010110101110110110001111011100010000000111111010000011100010;
#1 $display("%b", po);
# 1  pi=207'b101111111000010000011110010010011010111100011101110011111001011100010100100010101011000111111101100100001111111111011101001001111000011011011110011001001110010001001110110111000101110101100100011100001101101;
#1 $display("%b", po);
# 1  pi=207'b011010000011111101000110111100001011010101111111100000111100000011101111110001010001110010011001011000001111111101010010101111000011100001000011111100010001101110100000110011001000001111011001010010111100011;
#1 $display("%b", po);
# 1  pi=207'b110011101000101101001111111110000101110010011010101111000011101111010111000010010000011000010011010110110000111100110000010001000110101000111001101100111010010000111101001110111111010010000111000101011100100;
#1 $display("%b", po);
# 1  pi=207'b100011101001001010111100001101111100101000110010010110100011011110100100001110000010111010101100101001010100011111101101000100001111100111011101101111000010010110100110001101111011101110101000101001111111111;
#1 $display("%b", po);
# 1  pi=207'b000110010011011000100010010101011111101100000011000101110111111110000100010111111111111100100111100000010001011010100001110111011101010111111000111100100111001101010101111100001000010010000010001010110100000;
#1 $display("%b", po);
# 1  pi=207'b001001011011110011000010011111101111101010111011000111011111001001100111101101101001000010111011010011000000111110011001100101110110000001111101000101001111010100010110110011011101101000010000010110111001001;
#1 $display("%b", po);
# 1  pi=207'b100101100110001101111011010110011111011110010010111001010010010100101101001011010100111100110010110000100011001100100111010100001110010010011010101001100111000111100010001101101011010100010011111110110110101;
#1 $display("%b", po);
# 1  pi=207'b100110001111101101110011110110001110101000110111011100111110010011110100000001101000110000011001000111000000110011010110010110111101001010101001011100110001000000100000000101100110011010010110001011111010011;
#1 $display("%b", po);
# 1  pi=207'b000101010010111011010011110110000000011101000101000110000010111000100010111101001001101111100101111011101101000001011111111000100001000010000000010001111101101011000101110111011111110010100100000001001010101;
#1 $display("%b", po);
# 1  pi=207'b100111110111111100011001011100011101100101100011011001101101001100001111010011000001001011101101111001000011111001000010010111110110111111010101110101011011110111101011110010000111100100010100010100110011101;
#1 $display("%b", po);
# 1  pi=207'b111110110011101110101100010110111000011111111011100011001001110001111011001000000000011101110101011111011111000100010111001101010000110100111000101111001001010110110101010110111101001101001000011100100111100;
#1 $display("%b", po);
# 1  pi=207'b010100001110000110100010010011100001001000001100111110100001000110011101110000011001011110000101101101001111001010011101101010010101100000001000011010010000110000111001011000111010000010011110011011111010111;
#1 $display("%b", po);
# 1  pi=207'b001101010010110000111100110100001100010100110110100010001101001001101010010101100000011111110000101110011110111010101101000011011101111110010000001010101010110100100011101000100010110111001010010111010000000;
#1 $display("%b", po);
# 1  pi=207'b010100111010111011001001100001100100010100000110110000111101110101010111010011011111111000010010011000001000101000101010000000100011000110000100111010010111010011010110011001100001000010100011001100111000000;
#1 $display("%b", po);
# 1  pi=207'b011011011011110001101011101100111111000001011010000101010100100001010110111011011000010110111010100001101111111001000011100001111100011100110101110100100110010011000100101111101001101101100100010000110000100;
#1 $display("%b", po);
# 1  pi=207'b010101110000110001100011111011010001100011100001111110000100001000001001010001010110111010010100000001101011101010110110010100101010101101111101000101100001011110001110100111000011111011100100010001101011011;
#1 $display("%b", po);
# 1  pi=207'b010011110001110001001100000110011010111011000111101011001100111111100111100000001011100000110010000001100000110001001100111011000111101100011100101100100111110001101101000101101010111000111011111011111110000;
#1 $display("%b", po);
# 1  pi=207'b011000010110110000000000110000001001111011101100011010001110001111010010000110101010010001010110010100100111101010000011111101011001000111110011010101110011110101101011001101000011111001101111001100100010001;
#1 $display("%b", po);
# 1  pi=207'b111110101100010110011010100011101110101011111101000011111100010111101100001011011111111011010000000011011110101110010010111010100001001010001101010100101110100100001010100100111001000101001011001010000010001;
#1 $display("%b", po);
# 1  pi=207'b110110101010010010010101001001110100010110100010100011001000010110110100101001011001100101011100000110001000011001001100111001100001001011011100010110110101111101011101000011010110111111100010000110011101000;
#1 $display("%b", po);
# 1  pi=207'b110001101010100101000000010100011100001110000010000100100110010000000100001100000010100100100100000010101111100000100001110110100111000010001101110110111010101010111000110011101101101111000110001110101101111;
#1 $display("%b", po);
# 1  pi=207'b011100000110010000111110111111111000101001100110000101111101010100011000011001110001001000111111011111001000001010111101111111111001111011101111001101101010100001010111101000010101100001101110111100100100100;
#1 $display("%b", po);
# 1  pi=207'b111011010111001001010001001010110111001000000001001001100010001011100100000011111010000011111011000101101001101110101010000010011011011001100010110001110000001011011101010110100010011010000000110101100111010;
#1 $display("%b", po);
# 1  pi=207'b111100110111111111001111011101111000101100100011111000110101111111000000111101010100101111000010101111101011100010100110100111100010001111111011000110001110111011001101000011100110001000110010111011010111111;
#1 $display("%b", po);
# 1  pi=207'b001110000011100110011101111110001100011001101111011000010000101011000011001101110110100001100100000100101000010100010111000001110001010110101011000101011010000110100100000001110110000101110001010000010111110;
#1 $display("%b", po);
# 1  pi=207'b000101010110000011001001001100100001101011010110001110100001010010101000100101000001101000001010011111001110110010101110000011000100110011110000000000011010111001010001110000011000010101000000111100111101011;
#1 $display("%b", po);
# 1  pi=207'b111110101100101001101111110010000011110101000101000110101110010110011101011011110001011000001110000110001010010110000011010111110100001011001110000111110110110111010110011000101100001001011110100010101101101;
#1 $display("%b", po);
# 1  pi=207'b111111011110001000001001010011110101001100011100001000010110011101010011011101111000000101001101000110100100101011111010101001110101111111111111111101011011010000011111001110000010100100111000111000111110010;
#1 $display("%b", po);
# 1  pi=207'b010010110001010110111011010110100000100001001101000010101110100011111000110100011110001001001010101010111000000111010011110110101000101101010000011111000000100010101010101000011110000010000010000010001000001;
#1 $display("%b", po);
# 1  pi=207'b110110001011011001000110000111111000001101100101011001000100110011100001101111110111100111011111100000010110001101000011101111011101101010101111110100101100010000100011011010011001111010011010001011000010000;
#1 $display("%b", po);
# 1  pi=207'b101001011001010001010001011010010110010100101110110100000110110100101011011111111101100101110111101000010111111110111010110110110100100001110000110001001110110111111011111000000110101101011010011010101110110;
#1 $display("%b", po);
# 1  pi=207'b100100101100011111101001100100101010101110011001011010010010010111000110101100111001111100011111001111100110100101000100001000010111100100101111000010010000111010101010100001111000101100111111010001011001010;
#1 $display("%b", po);
# 1  pi=207'b000001011011111010100100111000001011110111101001111001001101101000011101101101111111100010010010111001101101111001110110000011110111011000111000001100001010100111010100000001101101110100111011011001101001110;
#1 $display("%b", po);
# 1  pi=207'b010001101001100001101110110101010110011000011101010100110110111110110110110011010000001010101111000010010010001010100101100010010001000011000100100110010100000001011000100100000101011001010011111010000111010;
#1 $display("%b", po);
# 1  pi=207'b010101101001111100010011001010001001111001010101111111000001010100111100110110000110000011110110000110000000011000101010000010101101111100000001110001000010000101111111000011000110001101101110101100000110001;
#1 $display("%b", po);
# 1  pi=207'b111101110000111001001110101110111011100010101100101110001101010111001000110110101000000001100101101111101100100110011110000101100111110111111000111010011100001010111111000110100111001110100011010110000101011;
#1 $display("%b", po);
# 1  pi=207'b110100110000001111101000101000010001100110010000111110101010000110011100101000011111110100001000001000010011110011000111001001110011101011001011100001101110110011110000100001101001010001110101000111110111111;
#1 $display("%b", po);
# 1  pi=207'b001111111110110100001011010011011101101111001111010101001111000000001011111101111000101101110010111111011001000011000000000111011100100110010011100010000001010101101001110000100000000101010110000011101011110;
#1 $display("%b", po);
# 1  pi=207'b010011000001110010000010111001110101010010100101100110000101101011011001100110101111100101010111111010111000111001000110010010100101110010100010101001100111111010100101101101100100011010101000111100111011000;
#1 $display("%b", po);
# 1  pi=207'b010001100101000011111101111101001001111010110000111011100110001011010011010100100010001110000011101001110010111010010000110111110101011100001100010011011110010011001110101000111101101010110011101010010011110;
#1 $display("%b", po);
# 1  pi=207'b000100100101000101111100100000111001110001111111000101100100111000011110000000100001000011001100101000100001000110101010000111011110011011010110000111010000101110010101001011010101101000100001110100100010000;
#1 $display("%b", po);
# 1  pi=207'b001001110101001111100100101010000101111001010100000001111011010010101100110001111100000010000011110000010011001011001111111101010001100001011000110010101100010000000110111111111111101010011000101000101101011;
#1 $display("%b", po);
# 1  pi=207'b110111010100011000110011011001110101100111101001100010101000110110100011001101000010001000000101010101101111110000000100010000010010101111001100100000011110100111101000010100000101111000000010110100100001100;
#1 $display("%b", po);
# 1  pi=207'b101001101001011110000111100110101000011000011010000000110101001101111001000010010011001101000011001011010100011001101000000111100111000100001100110110110001011110111101100000000001001011110010011010110101011;
#1 $display("%b", po);
# 1  pi=207'b010110100000100101110100000110100110010100110111111100000100011101000001111010010010101001110010110011100111000011000101101110010010000111101001101100010001010001011010100011011100001101110000110111010111100;
#1 $display("%b", po);
# 1  pi=207'b100011101100000111011100010000100110100110001000010111100011001011010100000001101001011110010001011110011101011010000010101110111111010001110101101000101111100010101101011010101011011010110101110000001011000;
#1 $display("%b", po);
# 1  pi=207'b011001010011100101100101000010010000111010101110010100000001000111101011100111000000101001101011011001011010000111101110001010011000101000101000010110011001110100000010111010110010101111011101010111001000101;
#1 $display("%b", po);
# 1  pi=207'b010001011110101111011110001111110000011101100010011011101010101111100101010011001000011001010101001100100010001100011000111001010001101101001011111100000100000010000111111101111000001011100110100000010001111;
#1 $display("%b", po);
# 1  pi=207'b100100011111000010101011110000111000001000010111111100110010111000010001010101001010010001111000000101000010110001010111101011101000100101001000010100101011011011001111010110010100101101100000101001000001100;
#1 $display("%b", po);
# 1  pi=207'b100010010101010011011000010000000011000001101010111111000011101001111100000111000001110011011001111010110010010111101001111100011110111010100100010111100011001100011000111111101011111101111101001010001010100;
#1 $display("%b", po);
# 1  pi=207'b101100111101011001001100011101100101011010001110011011001000111101011101100111000101101010110100111010010011010101110111110000010101011111111011101101000110111011101101011110001010010011000110011111110111010;
#1 $display("%b", po);
# 1  pi=207'b100101101000101000101110101010100100010110010111000010101110010110101100000101000110111000001010010110110010110111001000110000001110111100000100010111111001011100111000100101110111011110100110001001101110100;
#1 $display("%b", po);
# 1  pi=207'b000111011001110100101010110001001100100110110101100101101000101110101110001111001001011000110100001001011001011010110000010011100000011101011100011111101100101100001110100100000000000100101101110010010111100;
#1 $display("%b", po);
# 1  pi=207'b101010010110011001011111000101100000011001001000100110110111110001010011110111100011010000111110101000101001100110110001001110101100000010010110001000010100100000011001101110101011010001100010001010101001000;
#1 $display("%b", po);
# 1  pi=207'b010010011101101111101011110000000111001111000101011100100010011101101110111100010101110001100111111010111001100000011100101101110010000111001111101101011101101011000011110000000100000101110010110100110101101;
#1 $display("%b", po);
# 1  pi=207'b000101010000010000010001000001011011111101110110111111100010110001000101111100111100010011100001100011010111101110001001011100011000010001011011010101101111101110111000011111010011010110111001110111001101010;
#1 $display("%b", po);
# 1  pi=207'b101000110111101111011110111000101100110001010011110110101000111010110100011110110001110000011111111001010011111101000011101010001100000011011000010100111101101010101111001111001101111100111010111111111010111;
#1 $display("%b", po);
# 1  pi=207'b001100001101011011010101111010010101010101000110111001111010101011011011011111011110111101100110011101100011101111101010111101001111001010010100001110001000011100000011100111011000010011011011100011101000111;
#1 $display("%b", po);
# 1  pi=207'b110011000100101100111000000100001100110100000100111101100000111110111000101110000100000100000111011100000101101011010000011001001110001111011010011010001001110110000001100001010011010001011100010010011101101;
#1 $display("%b", po);
# 1  pi=207'b001101100000000011110011011101111111110010011011100110110000000001000100000100001111111111000101011000011001111011011001101110011010111000010001111011101110100010000110010100001010101010111001100010011001111;
#1 $display("%b", po);
# 1  pi=207'b011111110110001101010001110100010111010110110011101101001100001100011000100101000011111001110001110001001001010101110011110011001011100111011111011001111110100000100000110110111101011101101010010101001100010;
#1 $display("%b", po);
# 1  pi=207'b010111001101110011101011100010101101011011100001011000111110010110001011110100100111110110001010010101000011101110000101101100000111001011101111000100101010001100001111001011000010100011110001001101111100000;
#1 $display("%b", po);
# 1  pi=207'b110110111110001001000101100101011011100111110101010100110101000100111000000101101011011110000011011111011100010110111111010000010011011100100110001010010111110010001101011001100010101010010101001111001000010;
#1 $display("%b", po);
# 1  pi=207'b000100001000111010010000111001101001001001011001100110011011000110000111011101100011111001101100000101111111110110101010110100000101111111010111110100100000001100011101110010100100110110001011011010011110011;
#1 $display("%b", po);
# 1  pi=207'b010010010110001111001100110010100000111101111100010001010111100001100010101100011111100100101101101001100000010101000100110110101110011001000111000001010101100110010110100100010111010001100111010101001101101;
#1 $display("%b", po);
# 1  pi=207'b010101100000110000100001110010001000100111101101010101110001100000110010101101100000110011101101110111010000011011100100011000000000111111101001011110011010111100100010100001001111100010101100111011011001000;
#1 $display("%b", po);
# 1  pi=207'b011001101100011001101011000101011100100001100111111000111001010101100001111100011001110100001111111010101001101001111010101110010011011000101101100100010000011110001100101111010000001100111100001110011111111;
#1 $display("%b", po);
# 1  pi=207'b110011000110110110000011100001110010111011110000100101111001000010100101110010010111000111110111011011110001110110000001001011010100001110000100001001100000011011110000000011001000010111110011010011100100001;
#1 $display("%b", po);
# 1  pi=207'b010101010101011110011111001100011011011001011001010111001110110111101100010010000110011110011100001011111101110000011001100001011011110011000100000110000000110010111011100111010010100111101001100111111010110;
#1 $display("%b", po);
# 1  pi=207'b011000011000010101001110000010110011011010001001110111111010000101011011110011011110001000110101011111010010100111100111100011111001100010100000101011000111001110010111100111111111000011100101011111001000100;
#1 $display("%b", po);
# 1  pi=207'b001111110011010111010010111110010101101000000010100011001101001001101111100010010100000101100101111101000100100010000001011101010100110110011100101110010110011111101011010010010011011010010111100111110110000;
#1 $display("%b", po);
# 1  pi=207'b000111110111101101000001000110001101001111000001111110111001100011001110010011010110111100100000001000110100100001000000111010000110101001010001000000101011110110011010001000011000111101000000000000001011000;
#1 $display("%b", po);
# 1  pi=207'b001001010100001110110010101001110100100101000001101110010111100101111110110000111010011010000110000111010110101110111101110001011110011000101000101111101011101110000101011111110011011110000100011001100011010;
#1 $display("%b", po);
# 1  pi=207'b011101000111101100011011010101010000010001101101101010010111011000010101101110111000011010111000110000010001110101000011111011110001111011011101111011010111001010000010011010110101010111100111110011011000010;
#1 $display("%b", po);
# 1  pi=207'b100011010111111111111111101000011001111110100010111100010101011010010110111010101100111110001100100101000110100010010010110000100110100100100101011001001110100010000111010000111000111100101000110100110010111;
#1 $display("%b", po);
# 1  pi=207'b100010000110001001001111110011111100100010110000010101101001100100100000111110011110110000001101101100111000001011011100011111011011010101111111000100101110100010100010000011100101010001010001001000001100111;
#1 $display("%b", po);
# 1  pi=207'b110101011000000000110101111111110000001111000111111110111110101000010110101011110100000000011110101101001100101000100001101101000110000011111000100110100100110010011110110110110111010010010101011100010010111;
#1 $display("%b", po);
# 1  pi=207'b100101111000101110010111100001110101110000000011000110001010011101100000010100001110011000001101110111100111010000001011011001101011010000000100101110000011100001000111101011011101111100001000101000101011111;
#1 $display("%b", po);
# 1  pi=207'b111010011101001110100001110111100110100000000100010000111010111101011110100111101100111100011000111100010101010001000101111111001010000101100101101000011111110000011100000001110101011011101100000111111000111;
#1 $display("%b", po);
# 1  pi=207'b111111000111010001110100000100110101011011000011110111111111110010001011000110101100111111111101001010010101001111110111110111001101001001101101111000011001011011010101101110111011110101101000101110100011101;
#1 $display("%b", po);
# 1  pi=207'b111100010010011000001100011110000111001000100111000101011000001001011101101000101100011011011001010000000101010110011110101000111100111000101101001001001010010010111011100110110001111111101001001011100010111;
#1 $display("%b", po);
# 1  pi=207'b100100100001111110011111100110010101000100010111111010000010010111100010000000111101110010000100000111111101111001010100010110011101101010110010111010100010111000100100100001111111011010110000001110000101010;
#1 $display("%b", po);
# 1  pi=207'b001101010100100100001101001011001001001110100111110101011001111011101100110001111001001100110001111100110011110011101110001100101000011011001000010001000000000000110010010001010100101111001010010100000010100;
#1 $display("%b", po);
# 1  pi=207'b111101011101101001110000000110111000100111111110100101110101100101110100000011010110110010100111010110110101110011111100110001101011001110100000101000100110001001000000010100101101011101111000001010010010011;
#1 $display("%b", po);
# 1  pi=207'b110101110001001101001010001111010101110101011011110100101111010110010101001011010010110110111010001011101010011001100110011011100101111111011100011100100110001000011000000110101110000010110111101100111100001;
#1 $display("%b", po);
# 1  pi=207'b111000010110100101000101110110000001010011111001101000111000111010101101011111110001101111100000001110010111101001000110000000100101110110101010101001100110000001111011011001011110011110101001110001100010001;
#1 $display("%b", po);
# 1  pi=207'b101100100011010001011011100101010110010010111001000010010111100010000001001000000001111110000100110000100000111011011111110111000110011111010100011011110111111010100010000011001000011111010101100100001100001;
#1 $display("%b", po);
# 1  pi=207'b111010100001001011111000010001100100011100001010000001101100011000111101011110111000000111010001110011001011000010110101100010111100010110111101000110100110111010111010110001000001101100111110111100001000011;
#1 $display("%b", po);
# 1  pi=207'b111111000111110110100011000010001000110101100001011010100100011111101101010010100111001010111010111010001001001001010100111110110010110100110001101101101100010010000101111111111010110010111110111000101010000;
#1 $display("%b", po);
# 1  pi=207'b101101110000011110000000000101100111111000110100011110001111110011100001010110000001110001111100110001010111100010100000100101000111101110010111110110111011000101011000100000011011001110001100010011100011010;
#1 $display("%b", po);
# 1  pi=207'b100100100000111001011110110001000111111110001011100110010111101000011100011011000110000000111110110000011001111000100000011111011111011111001101111000001001100000110001010000010101001111001010100011000001000;
#1 $display("%b", po);
# 1  pi=207'b010100101000110010000011100001111110001110110111001010000011101101001101100010101101000100010010001110000111101011101110100111100011100001110011101101110110111011011001011101111101011011110000100011100101111;
#1 $display("%b", po);
# 1  pi=207'b111111011011001000011010000100110000000111110101010110011001110101111110100100010011000000100011111111000010010110011110001000001011010100100011011000000011000000001000101100110101000111011110100100111101000;
#1 $display("%b", po);
# 1  pi=207'b110000110010000110001010011000011100100101000000110111000001000000000101000010011011110110100111100100100101010100110001011000011100100011000111001101011100111110010000101100010001001111010011000000010111001;
#1 $display("%b", po);
# 1  pi=207'b111000000111110000111010011010110110011100110010110110100010101101001100000111100110101001101111010111110100000100010100001110111010011010011100001011001100101111111001101101101101100101001100001100100110010;
#1 $display("%b", po);
# 1  pi=207'b000101001100011001010100001100000001101101000011011010100101110001110001100110110100000110011101101101101011010010011010110111001010001001010110111001100110101101011100001111100111011111000111100110111001100;
#1 $display("%b", po);
# 1  pi=207'b011010000001111001000011000011011000010011001010000010100001101100011110011011011001000011001111111011111100101110010000010111100100110010110111111111111110011011101000010101011100000100011111110001111101111;
#1 $display("%b", po);
# 1  pi=207'b111111000111010001001010010011001111011111000100111100101011110011010001110010010100100110101001011010001011010110111000110010110011011100101011011000001000010111100111110001000100001000110100101100110110000;
#1 $display("%b", po);
# 1  pi=207'b101011000000101010110010001010100111111011000110000000110010100100111011101001111001110011000011111011001001001110110000011101100110010011010111001110111111000111111110000101001001000100100101100011001010101;
#1 $display("%b", po);
# 1  pi=207'b000111001101001001001110010101110011111111001100010011111000000011110010000101011100110001110001111011010011001010110100111010111111011000100111111110101011011010100001110000001000001000111110110010010111101;
#1 $display("%b", po);
# 1  pi=207'b010011010011000001100010011101101110100000100111001110001101001011001100001010011010110100000011001010011011100001110011110010100110011111010010110110011011111000001101011101101101010000000111111001010101110;
#1 $display("%b", po);
# 1  pi=207'b011000011011111001010001110000110101011100100001000001100010011100101100001110100010000000001101101101111010001110000010010101001011011110001011111000100000100001101001100011010000000001001101001000101101100;
#1 $display("%b", po);
# 1  pi=207'b101001101000101000101001000100110011101110110100010111011111010110111100110111000010000011000111100111010110011101000001101100000000001001010111001101010110001110101100111101010001011001100111101000001001111;
#1 $display("%b", po);
# 1  pi=207'b110001010100110010001110110101011011011111000010100010010010111011100111011100000011100100101011000110010001000110101001101011001101101011111110010111100110011100100110110110011100011101100010101111111110001;
#1 $display("%b", po);
# 1  pi=207'b011100000111111011000100010010000011101001010111010000011110011110100100010101010110010101110000100001101111010101010011000010001100010010010001001111101010010000001011000000010000111100000001011000110100000;
#1 $display("%b", po);
# 1  pi=207'b101100110110000000100101011111010100100111000111010101100010110111000011110000111111000001000111010010000000100011111110010100111100111111110011111001000010101110110110110100110011000001110000101101100100011;
#1 $display("%b", po);
# 1  pi=207'b101111111100010100011111111001000010010100001100100100101110101111101000111100011001011011010101100101000011010101011110010111110011101111010110111001101100000001010111100010110101011001011101100100000001111;
#1 $display("%b", po);
# 1  pi=207'b110101111101101111100010100101111011000010111101100110100001110001000010110110100110000111100010111111001010000000010111001011110011111100001000011001011101100110100011001100001110100111011110001000101101100;
#1 $display("%b", po);
# 1  pi=207'b001101101101111101011001111001110100011110100111001011011101001001100000111111100111000010101101001011000101011010111101010011110111010111101000000101111101001001110110010001010010101000011011001010100100000;
#1 $display("%b", po);
# 1  pi=207'b001110111011001000000000000100100011001101011100010011011000111111111101011111011101100001100110111011101011110111001100111110100010011110100011000110010110111011110111111101100110111001001111101101000110110;
#1 $display("%b", po);
# 1  pi=207'b001011011000000010011101101111010111011000100000001110011010101110110011000001000100101101000100101001001001001101111111001000010100000111001111110010001110001000111000111110100000001100100100111110100101001;
#1 $display("%b", po);
# 1  pi=207'b110111010100100001001000100111000100111110111100111010000110000100001110110001001100000111100011011000000001001100100010000000111001010010011000000101010001101011111011111100100011101101100110100001011010010;
#1 $display("%b", po);
# 1  pi=207'b011111101001010001110011110011111100110010011001000101010001001101001011111111101101001010101001011001001101010000111110110101001001110100001111101001110010100101111000100111001111001001010100001100001110100;
#1 $display("%b", po);
# 1  pi=207'b000101100110000001110000110101111011010100000010100010111100100000011001011000100011101001111111001010011111010110000001011101101001110100001100010111101011100101101000111101011100011001100100011110000111011;
#1 $display("%b", po);
# 1  pi=207'b100010001100001010010110000100100110011110001100111000001010100000001001010100010100101101111001101000011110101001111100100010001011011100001000110100011011100000000100110110010001111010011110101010111011110;
#1 $display("%b", po);
# 1  pi=207'b111011110000111001010010111001101010111101001010111010011011100101111100000111001000000110100010001010100001000010110000101000110110000000101111111111100000000000010011011111011111100011111011110001001011110;
#1 $display("%b", po);
# 1  pi=207'b010100110111100100101010110101000010110111011001010001101111111101000010100100111010111011001000111111110111001001110001100011001110101000010011010111101011110101000110010111000101110100011101001100010101011;
#1 $display("%b", po);
# 1  pi=207'b000000001111010100110100001011000000000111100100001100100111001110010000101001101001101111101101010010100101010101010001111111110111110110001010010101101001111100101110010010001101011010100011000110001111111;
#1 $display("%b", po);
# 1  pi=207'b110111011100100000001010101000011010011010001011100101001001111100100101000010110010111111000101100001111111100010111100111101111100101010100010100011111011000101001110010111001011011000010011011110001111101;
#1 $display("%b", po);
# 1  pi=207'b010001101000010111100001100100100001101110111101110001011111101000001011000111101101010101110001100110110000110101101100110100111100101100011100000101100111001101111010100101001000010111011110000001100110111;
#1 $display("%b", po);
# 1  pi=207'b100101111000011111100101100100110010111011011010100100010101110011101011100110110101011100010101000011001100000110111100111110011100101111100111011101001000101110001011101000001011110100001001110001000110010;
#1 $display("%b", po);
# 1  pi=207'b011001001110111010100000100110010010111010110011100010110011000000100000101000011000100101011101110011000110111001101111110000011011101010111101001111111010111101110001110110000100000111001001110010111111000;
#1 $display("%b", po);
# 1  pi=207'b111111000101111101001000101101001011111101110100111110011111000011000110101000110011110001110000100110111111110001111100010000111110001100010100100110100110010110000100101011101101000001100011100100110100010;
#1 $display("%b", po);
# 1  pi=207'b010000001111001101001101101100101011101010111100001111000011000010100100111110101001010110100001100110011101100111101110010111000110101011111100010011000010011101111011011101010110010001011001110111110111111;
#1 $display("%b", po);
# 1  pi=207'b101111100000101001000111101011000001110011011101000000011010110101111011111111100110101010000101001010110000011010001110011001011111110011000001001100101001000000100001011001110110010010010100110110101001001;
#1 $display("%b", po);
# 1  pi=207'b010100000110100010000001010000010010101001101100101110110001100110010101011001101001110000111011110111010001000001011000101100001011011011111000010011100010101011111010110100000111001111011101001011111101010;
#1 $display("%b", po);
# 1  pi=207'b110100100100100101110100111010010011001100000011101001011000000100010011110001111100000010001011011000110000011011001010000001011011101110100011010001000111110011010001001000010010100111001000100011100110110;
#1 $display("%b", po);
# 1  pi=207'b101010111011000101011001001111011011010010110100000010011101001000111100111100000101110011101001000011101010100100011100011010100001010010001110111011001111010001110010111100001011111100101011001000001010001;
#1 $display("%b", po);
# 1  pi=207'b110011000000010011010111111101100001001010100010010011011001100010010010110110010100111010110011110011100101010101001111001001011101010001100001101100100011110000011000111011000101100100111110111011001111110;
#1 $display("%b", po);
# 1  pi=207'b010111011110111101100111010001110011000100001011111000101110011100000110101010001101000111010010011110111000001000001010011011010000100100001110000010101111010000000101101110110000111101101010000101011001000;
#1 $display("%b", po);
# 1  pi=207'b111011100011000111011110111111011000011011000110101011011100100001100010001011011010101011100001101111110010010110111100001011001100011101111110000010100000010100101100001000011011100000001100110101011110110;
#1 $display("%b", po);
# 1  pi=207'b110011111000111000011101000011110001110101101101111001011001111001010101000010111101111101000001100011010011101001010000000111001001010001110110010111111000100010001001010101100101111110101000110100000110001;
#1 $display("%b", po);
# 1  pi=207'b010010100010111110001100111010000110010111100100010011100011011110010111000110011011101110011000000100001110010011011000000000011111001000011110111101001001001000000001011101101110010010101101100100011011001;
#1 $display("%b", po);
# 1  pi=207'b101100110100001110100000111101101101111000101000111111101100100011100000000011000011001100100011001110110110111010001100101000111011011000100100011000001111000001001111010100101111011111111110010011011111101;
#1 $display("%b", po);
# 1  pi=207'b001110000101101011011011110001100001101001011011101110101011110111100110010110010101111001100010001010010101111001010001011101011000111101010100110111010010010101110000010100000110111101010000010000001010001;
#1 $display("%b", po);
# 1  pi=207'b010001001110011010101011001011000000000010101110100010101111001000010100000001110100101101000010111101001101001010100101110000010011101101001000000110101001111001000000101000111101100001101010111101110011101;
#1 $display("%b", po);
# 1  pi=207'b010011000011100111001001101000101001100111001000011010110010111110111111010011000011000110100010001101101000011101011101001000000110110111111100101001011110111111100111000001111001101001001001011001000011111;
#1 $display("%b", po);
# 1  pi=207'b010000010001100001011110000000000110000110100011100010110101011100110100011110100110100110010001001010000100000100000110100110000111000010110001111110111111001010001110110010100000110100101011110111001000111;
#1 $display("%b", po);
# 1  pi=207'b110001000110010001001111011010001010010011011100100010111101000010100010000111101011110011100011100110100011111000000100100111011010001100010110000111011001000001100011011100000000101110100111001001100000110;
#1 $display("%b", po);
# 1  pi=207'b010001000001110000111001100010101110111100101011010001111010101001100101100000000101011001101000011110111110011110011101111001000010000000011110001100110000010110111011110001110111101000101101100100001101010;
#1 $display("%b", po);
# 1  pi=207'b000011111010011100010100000001010001010011101110011010110010100101001101100011100001010100001011111101100101011111001110011001011011100011111011011101100111000110110111010001000111110010111011100011101110101;
#1 $display("%b", po);
# 1  pi=207'b101110010101010000001000011000110110110000010011000111001001110011100111111000110011111000101110100011010111101010100001001000011010000110001110000011101111101010111010110110011001010001101100001000000010101;
#1 $display("%b", po);
# 1  pi=207'b101100001111001100010010101010000001101101011010101011110010111111011110000110011101000111101111011010001101011100111000110100001001111100011101001000100000000001101101100111101010001100001011010010101001011;
#1 $display("%b", po);
# 1  pi=207'b100011111101010111110010010011011000011111000110110010100110110101100111100101010000010111101010000101100111000000101010111000001000000111101100011101000101101100010101111001101010100100000101101011101100010;
#1 $display("%b", po);
# 1  pi=207'b001110010010011010010110111101000100101001101110000100001100100001001001111001011100011001110110111011110011111111011100101000100111110011100110100010100100111000110000100010001000011100000010110111001010011;
#1 $display("%b", po);
# 1  pi=207'b010101010101101011001011101000101001001110101000111011111111101101100101110101101110001110010001110101000110100001010111101101111100100110000010011010110110100010011000110110110001110011001010010110001001000;
#1 $display("%b", po);
# 1  pi=207'b101100011100100100011100011010000000111101101101001011110100110111010111101011010100101011000001001111010001111111001001011110111000110000010000101011010101010010101101101011111011101111010001001001010011000;
#1 $display("%b", po);
# 1  pi=207'b001110101001100111111100010001001101010010010010111001100010100001011011010011111101111110011010001100101110111101000101001000100110110110010101011101100101110001110111101001000101010101101110101000101000100;
#1 $display("%b", po);
# 1  pi=207'b000011001111000100100100011111011110110111011100011010111001000011111010010100001110000010011101001110011010011001101111111011001001010010100101101011111000101001110011100001110001101011101011010001111001000;
#1 $display("%b", po);
# 1  pi=207'b101011011001011101110010011001011001011010111000010111111001000111100000001111000101100101100110011111101001001110001011010111010001101001000001101001011110101100000001101010100001111011010000010011110001101;
#1 $display("%b", po);
# 1  pi=207'b111000011111101111011110001110111000110100011011011011011010111110000111111101010100101011011011100011101110111111001010100010011000110100100110010011010010000001010001010101100011001001100110110001000011100;
#1 $display("%b", po);
# 1  pi=207'b010101111110110000011100001100000011011001100001010000010101100101110011011000110101011100100101000001110000100010001100100010101011101011110000100011101111001100101001110001100010110010010100001000010010001;
#1 $display("%b", po);
# 1  pi=207'b010010011001100110000010110000011011110010000110100000110111011010110110110100000011000001011110011110011010011001110111101101111010110110100111011011111001111010001100010011011010101111001011000001000010000;
#1 $display("%b", po);
# 1  pi=207'b101101001000010001110101100001011010001111010011101111110101111101100101000010111111101101111011011110010011111001110100101100100101100011100110001101001001111100010111011110100000011100000110000001000000110;
#1 $display("%b", po);
# 1  pi=207'b111100001111110100111000110000010111110100111001000111011110001001110010010111111001101010111110010101001000001101110111101111011110010111100001111010101101110110100100010111110111000000101011001011010010011;
#1 $display("%b", po);
# 1  pi=207'b110101000100111101100011000001001100101111100010111011010101010001000101111110100110011111110101110001011001011101101011000111000010100101000100111000001110100110110111100010111011000111011100101111100111011;
#1 $display("%b", po);
# 1  pi=207'b001000010010011000000101010000010100100011110110111000001001101000111010101110110000011111001100111010100000110101011110110001000101101011110000100101001010011101111000010011110100110101001011101010100001101;
#1 $display("%b", po);
# 1  pi=207'b101101010101101011001111001100111010110000111011010101100000110101111010000000001100100101000000000010100011100011101001101110010100101011111101101111111010111011111001000000111110011110100001101011001101000;
#1 $display("%b", po);
# 1  pi=207'b010011100111010101001011011001000001111011111011101000010010001010011101011111110101100101100101111100101111101010011101010010100100110110010010010100101110011011100001100011101010110101111101010100100001001;
#1 $display("%b", po);
# 1  pi=207'b010000101001110000110100101000110110001010011101101010001001111010010100011000010101101101100100011010011010111101011010101111001110111000100001001011110111001111001110101110100100100110000001000001010110011;
#1 $display("%b", po);
# 1  pi=207'b011101110010000001101100010001100101010001011000011010101111100100001110000110110111010000010111110011000010101001010101100110100100101011101111101100001011101110000110100101001101010101001101110111101101111;
#1 $display("%b", po);
# 1  pi=207'b100010001110011000010100100001011110011110100101010111101000010101110101110101101010101111110111000111110000001110000000001110001010011101010111000111110101110100110001101010110000111101010001111111000100000;
#1 $display("%b", po);
# 1  pi=207'b001000011000001111000101000110111000111100101010010011101010100111000000110000100001001100100000010010001010110000001101101110000000000101001111101011100000010010011100100111101110011110100111100011110100110;
#1 $display("%b", po);
# 1  pi=207'b000010000001111110110001111010100101101011101001010010101110100100100001101100001010111001100010001100001001100101101010100100001110110001001000001111001111011010101010100000111001001110011101011110110100100;
#1 $display("%b", po);
# 1  pi=207'b010010110101001110000010001111001001010000101111010001000001100100010010100000111010101111010001110011010101100111001000000001101011000001010110100101010100100010111100011000110100011010100111110010011110011;
#1 $display("%b", po);
# 1  pi=207'b110010110100111000011000000011011011100100011100001001000110111101101111111010000011001101000100010110110100011101100111001100011100000000000011110110011101011000101010011101111111111010100101110001111011001;
#1 $display("%b", po);
# 1  pi=207'b101100011100101001010101100101010111111010110110101111000010000110000000101010001001001001100111011100010011110100100110001101000010011111101101011111111001101011111000100000001000000110010001111100011000110;
#1 $display("%b", po);
# 1  pi=207'b111001011101110111010100101111001110100100011001010111101000011111001011100111000100111000011110010100111011101000001110100000011011110011101011011110011100110100100110101100001001001110001011001010101101111;
#1 $display("%b", po);
# 1  pi=207'b001011110010110011110001011111010101011000001000111110101011111001000110001100000000101101000100101001110000000011100100100101011111011111111100111011000000110011010000100100001111101101001110011001011110100;
#1 $display("%b", po);
# 1  pi=207'b101001011101111100110011000001011001101001001110110111010001011111111011111001000010011111010010110001000010110111010000111110111100110111100110100001100111000110110001101011100111011010011111011010001111111;
#1 $display("%b", po);
# 1  pi=207'b110101011001100110010011111001010000111100000111000110111001000110100011001011011111110100000000000011111000000110011000100000111001111100001101000101110101010000101001010110001000100010011010001100000001110;
#1 $display("%b", po);
# 1  pi=207'b110011101100101100101011101111001011100111001000011111010100011111100110100100010000000011101000010101111010101011010101010110000000011001110111010100010110110101101001011001100000110110011100010000001101100;
#1 $display("%b", po);
# 1  pi=207'b100111111001001100111100000001000111001000010011000101111110001100001111111000100101011100101111100001110100101110000001110111010110011111001001011101111111101100110010111011111110010110100000001011000111001;
#1 $display("%b", po);
# 1  pi=207'b011100100111001010111000101111110011000011011101011011001010000000111001111010010010001000001001001001111100110111011010011111001101101101111111101001101010011011111011110101000111110000110100111100010100010;
#1 $display("%b", po);
# 1  pi=207'b001010111000111111010100100101001010001100010001010111011110100100100001010111101101001111111110111010100110111100000001001100100000100110100101010000111110000000101010110101101110110011000011110101110001011;
#1 $display("%b", po);
# 1  pi=207'b001010101011101101000010001000011011000001010000000011100011111010101010011111000101011101100110101101000101100011000111001000011100110101011000110001111110011001000011101111100111001010000010101100101111010;
#1 $display("%b", po);
# 1  pi=207'b001101001001101101100011000011100101101110010011010100111011001101100001010001110101011100010100111010000100111100000101001111100110001101111110111001101000100011100001001101000100111100000011000000100111100;
#1 $display("%b", po);
# 1  pi=207'b001101000010001110100000000011011011010010000100001110101111101000100110011100111000110000010111110110010000100010010110001100011110010010001000110110111010000101101101011001011001011010011111101011101001000;
#1 $display("%b", po);
# 1  pi=207'b101110100010000111101110000111100101000100001110110101101110101011011101101000100101101110001010110011110111001101000111010101101011011110010100111110100111010100000000100000010100000111011001000001000001101;
#1 $display("%b", po);
# 1  pi=207'b001000101111000100000101111101011111000101111111111100010111001010010100001001111111011000011101101110001101100111001011111011110001010101111111010110111100011000001111110011001000110111110010001100111111100;
#1 $display("%b", po);
# 1  pi=207'b101101010110011011111000011100001111110000010010001000110011101110111000100110000000010110110110110010110101000001001010011101110010101011101100000100010111000010100001011110011101111101111001101111011101101;
#1 $display("%b", po);
# 1  pi=207'b011010000100011011010010010010011010011111101010100101111011111000001010101000111000000001111111001011000000000101010100111011011001001111010011010110001010110011010011011000001111010010100011101110010101110;
#1 $display("%b", po);
# 1  pi=207'b010101110010111100000011100000010100101010110110000101111111111111001101001111101010010100001011111111000010111100001101100001100000101111001011010111011000000100010001011111001000011101100010110101101011001;
#1 $display("%b", po);
# 1  pi=207'b100101000000011110001111010110111010010011010101001111100100101111011110100110110100111110110010101111011010101000110001100110010111101110010111011100011100010001001101101000100111110011011110101111100000101;
#1 $display("%b", po);
# 1  pi=207'b111111001001001001111011001000010110010001100100011100011010001001110001101110110100011101111010011000111010101111010010010110110111111101100100001100000111000101101000000001110010011000110111011010100101110;
#1 $display("%b", po);
# 1  pi=207'b000111010011110101111110000000011000110001000110110100011010101001110110010101110110010011100100010011110101101101100111011110110101101110000000101111010000110110110011110110100100100011110011001101101011011;
#1 $display("%b", po);
# 1  pi=207'b011111111101110001001000110100111001100011001010101101001010000110111000101110011101010000110000011010110011110101100111111010111011011100111011110111110011001111011100011111000110110011010001100010100100001;
#1 $display("%b", po);
# 1  pi=207'b110011001010100000011101111110001110000011001101110000111001101100011110111010011001011000101111000001010101101011101111110011011010111110110010001010001010010101011110001000100100111101010010100011000010101;
#1 $display("%b", po);
# 1  pi=207'b110011101110001101001011101010010010101010110000001111010100011100000111100101110100100101000111101100011101000101101100111011111100110101001110001110001010000010001001111001000100111101001010011101000010010;
#1 $display("%b", po);
# 1  pi=207'b011001011100011111000011001100111101100001011100000100001101101000011011111101101001010100011011100010010010101101101111000000001000110000111010100010110101010011011100101001100011011000011110111001010100110;
#1 $display("%b", po);
# 1  pi=207'b011101011100010000110110010101001000000001110010100100111100001011111001000111111111010110100100111100110110101010111101101011000111010000001110010011001000100010011111111110010100111000111011111010110001111;
#1 $display("%b", po);
# 1  pi=207'b010110100000011001111010101001101100101111000001011110001001100010001110101011001111010010111100110010010101110011010100010000101011111000100010101101111100011000001100101011000111111001101001111101100011010;
#1 $display("%b", po);
# 1  pi=207'b001001011000000100001001100100001010100011011101000100100010100111110110000001110111010101111000000000011111010000001000001000101001110100111110000000111011100110000110101001010011010001000101101010000111110;
#1 $display("%b", po);
# 1  pi=207'b110001010010010110010001110010100000110101101101000011111111011010110111101110101000101001100111011101101101111111111011101110000001011010001010001101100110111000011011011011010100100001110111011011011101110;
#1 $display("%b", po);
# 1  pi=207'b110011011111110101011001010001100111111011100101100111001001010001001111110100110001110010111100101111011001001000111100101110011011110001111010100111110001110110000101100111101110110001101110001100100110110;
#1 $display("%b", po);
# 1  pi=207'b000101100000001111011110001011111100010010001110010101011000001010100100010011000100001000000000100010100000001011000010101100001100100001101011110000111101010011001010110100100001100011101000101110100001100;
#1 $display("%b", po);
# 1  pi=207'b110101001000110000110010010111111011111000110101010001101001011001001101111001011101101101000100100111100010010000111100010000010010010111011011000000011111000110011110111110110001100101110000111101001111010;
#1 $display("%b", po);
# 1  pi=207'b000000111010000010011010000110001001011100111110001101110111011011001011110011001101111000001011001111100110101111010100100100110110110011101111101110001001011110101101110101111101100010110010010111101101100;
#1 $display("%b", po);
# 1  pi=207'b010000101110110001110011010110111011111100110010100100100010100001010111000110001110010001101111111000010001011110010011001000100011010000111111111110111010111000111110001111101111100110111111100101001110010;
#1 $display("%b", po);
# 1  pi=207'b100001100111110101101011000110011001001101101101000100010010010111000000110001001000011111010010011100001110000001010101101100111010110110111000111011101101101101110110111001010010110110000110110010111101010;
#1 $display("%b", po);
# 1  pi=207'b100000100110111101100000010111001101010100110111110001110010111011010110011111000010110011000101011100001000101110011000110101000111010110111010000001100011101110111001100100000110111010100011110110110100100;
#1 $display("%b", po);
# 1  pi=207'b100100110101110010001010110000110011111011010011100100101101011000001010000011111101100010001101001111011110111101000111010110101011011000001011000000001101001010000001110101000001101100100110101000010010111;
#1 $display("%b", po);
# 1  pi=207'b011001101101011010111000001011001000110000000011101100101010111100011110011111101100111000000110010011010110010101011110101100010001010010101101100010000000001010000100000010001110111000010010001110100100011;
#1 $display("%b", po);
# 1  pi=207'b101101000000110000001011111111011101010000010011100100010110010111111101110111001001111011010011011100111001001000001000001000011000011101001011010001100100100111111100100100110111111101101110111001001100001;
#1 $display("%b", po);
# 1  pi=207'b110111111101110000001100101011101101110010110010101110111100101001000011101101011110000111101011010100101010000001111000110110001010101111100000001111000000101110011101111111000011010000001110000011001001100;
#1 $display("%b", po);
# 1  pi=207'b110111101010010100100111111111101100111000110100110011010000001101001011011010100101000001111110011010011111110100000111111110001101010101101011111000010011101011101111111100011100000110110011110001111011000;
#1 $display("%b", po);
# 1  pi=207'b010100111101110000111011011100001100100111001110110101100001101110000000011011000111101000111100101111110000011100100101011001010110010000011010001110110000011011001100001111000011111011000101000111011101010;
#1 $display("%b", po);
# 1  pi=207'b100000001001100100110011100101100011001111101011000011010111001010010011100011000101101000111100010100111000101110111101010001111000110100100100111100011000110110111011111111010101010110100101101000001010010;
#1 $display("%b", po);
# 1  pi=207'b110101011100111000111101010010011010011011000101110001001011110111001101010110000100000101111010001001111001000010001011010111111111000000000100110001011000110000001000000100001100110110101100001000000101101;
#1 $display("%b", po);
# 1  pi=207'b010010101001111110010011111011000101110011001000011111011101110111101110111000101111101010001100100000100110000111110001001101111000111100000110101100111101001100000000000101011111000110110000111101000000000;
#1 $display("%b", po);
# 1  pi=207'b010100110001011100101000000110111100111010001010110010111100101001001100011011010100011111101011011110110101000111110011011011001100101101111110011010011001101000110010100011011110110110101010101000101100000;
#1 $display("%b", po);
# 1  pi=207'b011011011101110010110100000000010010010001011110110011101111000000000100010111000100101011010000111101101001100011000101101001001110101101101111101000111111100000011110101100011011000111000010001010001011111;
#1 $display("%b", po);
# 1  pi=207'b101000001001101001001110011100001100000000110010010111111111101100100001101000111110110111110010110100001001011000011001110001111111100110001000010110010111101110001001010110000110010110011011011000000110011;
#1 $display("%b", po);
# 1  pi=207'b011100110110100011100101010111011011000111000010010000110001000011010011010000111000010011100010000110000100110001010010001001110001110001101011000000100001011100001100010000010101111111100000001000010100011;
#1 $display("%b", po);
# 1  pi=207'b010001011101110100101111111000001100011000011010000000001100011110001011101100101001000000010001011111011101000111110110100101110011110111100001000000110000010000111001101100110110010000011110011010101110111;
#1 $display("%b", po);
# 1  pi=207'b000111001011000010110100000111000111011100001010001100001101011111111011010110001010110111010100101111010111010101010011111000011111100111100111000100100011001000000011001000100010001111000100110010010100001;
#1 $display("%b", po);
# 1  pi=207'b100110101101100011110110000000001100011001111011111000101101000010001111010011110000101001001011000001101001011101110101100100100111000100010011010010011011111101010001111101011101110010010001111001010001010;
#1 $display("%b", po);
# 1  pi=207'b101010101111110111100111010100111111000101000101010110000001111001101100000100101011110111110001011101100100110011100110111001011000011111101011000010011101010011110100000111100011000111010010011011000111110;
#1 $display("%b", po);
# 1  pi=207'b100101011101010101000110000111000001101111011100010001010010001000011110100101011110100100010111010101000111101000110101011110100010100010100000011110001000100100110111101110110111110010111100101001001110010;
#1 $display("%b", po);
# 1  pi=207'b001110110000000010110011001101000011001100101100000101010111010001100100011010011110110110100111000111100011001110000111100001100011110101110100100010100011101010011100001111110001111110101101000000110011011;
#1 $display("%b", po);
# 1  pi=207'b101001010001101011011110111011110011100110010010100000100111101000010101010011110010010010001010010000100011000111111011011010001100100000000011000000011011010111001110110000100000110001010110110111110110001;
#1 $display("%b", po);
# 1  pi=207'b100111000010110010000010001101111001101000000111100001100001001100010111010111010000111011110001101000010011100001010110000010110100101111011010100000110100011001111110110010100010011111110110011000010111101;
#1 $display("%b", po);
# 1  pi=207'b110011001001011001010111101011100010000010010001011111111110001001111111111101001001000001000111001111001011111001010110000000111010011100101100011011001011000010100111101110110011111010100110000000011111100;
#1 $display("%b", po);
# 1  pi=207'b000001110110011101101110110110101001101100001100100000010011110010101001000111010100001000010111011110101001100101101100101001111011110001011010111011110100011001110000011000001101111000011110011101000001111;
#1 $display("%b", po);
# 1  pi=207'b110111110111101001001101110000100100001100010101101000010100000101100111001010101100111010110101010110111001110100110100110101111010110101011101000000110111000100110110101100111101000110000111111101001000100;
#1 $display("%b", po);
# 1  pi=207'b101010011011110010101001010101011011010101011000111011011000001010000000000011100100101010010011100101100101110010100010100100011010111101101011010010001101000011001001000101110111000100110101111000000111010;
#1 $display("%b", po);
# 1  pi=207'b000010011100001010011100110110111101000010010101011001011010100000010011111101110100010010111110010100111110010011111010110101110010111011001010111100010010000011101001111110110101000100001111110100101011000;
#1 $display("%b", po);
# 1  pi=207'b001111000101110001001010101000011001010111010000110110101111011101000100011110000001011010001011111101100110100111000101000001000100100110110001010001101100100110001100110100011001100110110010011101101110100;
#1 $display("%b", po);
# 1  pi=207'b001001001010001010110110010111111111011000110000001101000101101001000100001111110000001111100011101110110000000010011101111000001101000001000011110100111110100110111110100111001010110001101000101100101110000;
#1 $display("%b", po);
# 1  pi=207'b110101000101111010110011010011111101100110111011110011000111000010111111010011010111011010010101111001001001110000011101011001001110010001111010111001001111100011001010011110000101101111101111110100010110000;
#1 $display("%b", po);
# 1  pi=207'b110011000110101111111111011110110110010001010001110001110001101101101100101100001000100010001110000101010111100001001010110100100111001000000110111000111000111100110011101101011111110101010011010000100011000;
#1 $display("%b", po);
# 1  pi=207'b100101010100010011001100010000100101000010010111110001001001011110001001100100100100110000000101001110110101001101000011101010001011001101100100011001010000110100110100101100001001100111001110011010110111111;
#1 $display("%b", po);
# 1  pi=207'b110100111000101001010110011010001100000110010111011111010000010011000100110010010111101110001101010000101110111001100001111010110101110011000100000000011011010110000011100100100100000011011110100001000010100;
#1 $display("%b", po);
# 1  pi=207'b100010110111011101010010001000111001011111001101000000000101011100010010101001010101000000101001010101100011010010111111000100011011111011111101010000000010111100000110111001001010001110110111100101100111010;
#1 $display("%b", po);
# 1  pi=207'b110101110111001111111110110010101011000010000011111101101101100011100011011101000101100111101011100111000010101000111110111001100010011000000101001100011001110110001111010111010001011010111011010110111010111;
#1 $display("%b", po);
# 1  pi=207'b011110110110011000100010011010010111111101000100110010001011011000100110100101101110110101111111010000110010100100101001101010010110000101101100101100000111101110001010111101010111110010101111101001001111111;
#1 $display("%b", po);
# 1  pi=207'b110100001011010100010100001110101101011111100110111011001110111001010100010001111000110010001110000011110010000110001011011101010110111110111000001011111000010100100111110101001111110101100011111001000100011;
#1 $display("%b", po);
# 1  pi=207'b001011001100000000111110110100111010110100011010110010001001011100100010100111000000111001110010001110001000011010110000101110000101111001001000101010010100100000111001001001010111011001000000010010111010001;
#1 $display("%b", po);
# 1  pi=207'b101001110011001111100101011000111111011111010011101100001101100110011010101110000110101110101010111000001010110000100101000000011111010010010011100000011101111000100101011000000110001010110111011010110111001;
#1 $display("%b", po);
# 1  pi=207'b111011010110111011010100101111100100000011011111011011001011111110010000111110010001011001100101011011110001111010110111011001110101000101001100111010000000011101000101010101111110011000000110000101010011101;
#1 $display("%b", po);
# 1  pi=207'b101001010001110111000001110101110101101010111101001010101010001001101011110000110001001101000000111001111101101110001111010000011100111101111101101111111011001010010111011000111101101110100000000011011011011;
#1 $display("%b", po);
# 1  pi=207'b110111010001101111101110110101011110001010111001011110000101010001101010001010110011000101000001100001000100101001000100111111110111110010101001111100011111001000110011010001111000100110110111111111100101001;
#1 $display("%b", po);
# 1  pi=207'b101100110110010001100000010010101000000101010111000110101010100110101010100100100100001011100011110001110000110110100110101001111101010000110101110011000001000111110100001000100111000000111101010000000110001;
#1 $display("%b", po);
# 1  pi=207'b010100000100110010001001100000111101001000011000101000010010011011101010100011010010011110010111100010100001101110110010010001111111100001000101001111110111101111001000101011100110100001110000110101010111101;
#1 $display("%b", po);
# 1  pi=207'b001101010100101001111100010010001111000100010001101101101001011000111100110000001100000010000011100100111011100010111001011010101101101000001001111111001001011000101000001101010101101011111011011101010110000;
#1 $display("%b", po);
# 1  pi=207'b000100001000011111110101000101101010111011010101110110010001100111110110011101010011001011110000001011100101100010001111100011001100011111101011000110001011100111111010111101001100111000111110100100111011000;
#1 $display("%b", po);
# 1  pi=207'b010111111011010101110110010110010101000100001010101011011010101011101110111001101000110101010110110001111000001010101100010100010100110010100011101011110010011011101010101111110000101010010101010000111011001;
#1 $display("%b", po);
# 1  pi=207'b010101000010011111011010101111101111010101010011111111010100101111101010111011011110111111101000101100000011101011001001011011000001111100000100010110001001011100110001001010101011110101111100101100111010000;
#1 $display("%b", po);
# 1  pi=207'b001000000111010100010100000110100100100001010011000100101101110000000000100110011110000110111010110001101001000011101000101101001110001101010110111101011100001110100010000010010111000000110011001000111001001;
#1 $display("%b", po);
# 1  pi=207'b000000100010010011100001101010001111111101101001111100000010100010100000111011101101100111101100110011100011001111101110100101000010011110000000100101100100110011000101101011010111110010010010000001001100011;
#1 $display("%b", po);
# 1  pi=207'b100111110000000011010000101001100111010010110101010101100010110011000001001101010101100011000111011110010101111110111110000010001110001111010001010101100000111011111111101101111111000101001010100001000111111;
#1 $display("%b", po);
# 1  pi=207'b100010000011001101000000111101110001001100101111011110011100110011011011000100110011001010010101111110111101111001111101100111110000110110111101100000011001111010111000010100001011101010111010001011100101001;
#1 $display("%b", po);
# 1  pi=207'b111100100111001110001000010011010011101111100111011000100001011101100111101111011000101011001011001101010011001010110001111000110100110101111100010011001110000100100000011001100000101101100001111101010100110;
#1 $display("%b", po);
# 1  pi=207'b001001011001000100110000000111110110100100101011011101000011100101000110110101011011110101000010100110000001000101001001011110111100111110010001101100011101101001001110111000000011111111111011011010110100110;
#1 $display("%b", po);
# 1  pi=207'b110010111011100000010101010010001001011000000100101110001111010000001001100000001100010100111010010110011110010011101111110010111110110000110011011101111101010100011001010011001000011010000001110010100010111;
#1 $display("%b", po);
# 1  pi=207'b100001101001010001100011010001011011001101000001111110000111101001100010111111111101110110101010100010100011110100011001011000001100100010000000100001010101111110001111100000000101110011001000111011000010011;
#1 $display("%b", po);
# 1  pi=207'b001101100100011100001011000010101011011100100011111101001000010001111100010000101101010110101101000111101101110100100111101110101010010100000110001010010101100110101110110110101001111110000001001001100100001;
#1 $display("%b", po);
# 1  pi=207'b001011110100110111100101100100000100010000101100101110111000010101111101010111101011011101111100101000000011001110001110101010111010111111010010100001001001011011000110100011100111100000110001110001111111111;
#1 $display("%b", po);
# 1  pi=207'b000000000010001010001110011100101010001011110101100111100100010110100100111000011011001000011001001110010111100001010001000010010010000001110001101011010000000101001001110010010000010011100111110000010110001;
#1 $display("%b", po);
# 1  pi=207'b000111101100011111101010001111111010101111010000000111101100000011000111011011110001001111100100001000100100000000010101000110000011110111100101001100101010000001010001101101010010110110111000111010011110101;
#1 $display("%b", po);
# 1  pi=207'b010000000010100011001101001010001000111111010111011100010100111100101011000001100100001101101011001110000001010011110110001000110011110111100100000000100010001001101111100111010000100000000011111100001010111;
#1 $display("%b", po);
# 1  pi=207'b001010101110000101100011000101010001100000111000100110110000011011010000100101010110010111000100111111101110000001010101110111110100110110011101000010101000010101101101011010010100001101110100110000010100110;
#1 $display("%b", po);
# 1  pi=207'b101100110101100001100101110010110001000000001110010000100000011111110111011111000000010011100011100010011101111100110000010000100100010110111100000000010101110010100100000111010010110110001011111000100101000;
#1 $display("%b", po);
# 1  pi=207'b001010100000101000101000111100011101101000001001110110101101010011011101101010100110000010011111100010011100000100010010011011001110100011000000010011001110010000000010111100001011101000011111110000001101010;
#1 $display("%b", po);
# 1  pi=207'b101011100010001100101000001000111001100000010101100110111111111101000000001000100000000001110001001000010110101100001000001011110101101111001011000001001000111010010111000111101101010001010010111100110100100;
#1 $display("%b", po);
# 1  pi=207'b110100010101100101100010001110001000010100011110111000111010000110011011011000011010001000100000101100111101111000011100001000001100111101011010011010010011100011000100000110001110100100100000010110101011100;
#1 $display("%b", po);
# 1  pi=207'b011100000100001000010010111110010110100000101111110011001010110010100101101001010011111110101010000010101101110000101101111110001000101010111111001000100101010111101100101010010000111101011000110000000010010;
#1 $display("%b", po);
# 1  pi=207'b110100001011000111010010010000000110101111000111100110010001100010110011001011000100101010011010101000110100111010101000101100110111010110111100000101100110011111110000010101000111110110101100001010011001100;
#1 $display("%b", po);
# 1  pi=207'b111111110110100010101000000001000001100001101111110100000101100000100111001011000100111011100110010101011010010011001110010111111111011001001010101000010010101100000010101101110100101010001110111010111000011;
#1 $display("%b", po);
# 1  pi=207'b010110001011101100010000101111111000101111000101111010111001010011101000110010011100101001111101101101101011011110101011011011010100100010101101101000000001111100110111000001000110111100100011010101001001101;
#1 $display("%b", po);
# 1  pi=207'b011010110010111100010111010111110101101011010011101110011011101110001100011001011100011011101011111110011110010000010000010010100111111100101100000010011000101101110010100000010010000001100111101110011110011;
#1 $display("%b", po);
# 1  pi=207'b101101010000010111000011001011111000100001010110101110100111001000101011000000000100100010001000011011110100110100001001000000010111000100011001100000101111100001111110011111100000000110101110000000011011010;
#1 $display("%b", po);
# 1  pi=207'b100001010110110111001111110110111111010001001000000100101110100001011110111010000011111011100101111100001101000101101010111101101111010100001111000110110010100100001010000011101010100011011100110001000011010;
#1 $display("%b", po);
# 1  pi=207'b011000001001001101110101010000110111100000000011001111101011010110110100001001000100110111011111001101101110011110001010111111010100100101100111010111001110010111101000000110010001010010010100000111110010001;
#1 $display("%b", po);
# 1  pi=207'b000010010010001000111100001100000101001110101100000011011111101101011100000011011100011111001001110110000110010111100111001011001100010001011100100100001010010110110001010110111110000000100000010001011011001;
#1 $display("%b", po);
# 1  pi=207'b011100100110001011001111001010001101100011000100111101010000001110111001110111001110011101111011010000101111111001001010101111010001011010010101111001010101111010100111100011011100001011101111101010100010001;
#1 $display("%b", po);
# 1  pi=207'b011011001110010101000010001010110011111110001100100111000001010011100100011010010000111101111010100111011011001010100110101101001100000010000011000100101100010010101000101010111010110001111001001100110100111;
#1 $display("%b", po);
# 1  pi=207'b111010100100001011101110111001110110100001010101100000001111110000100100100101100001011001110011011100101001111111010000111110010110111010111111110100100010000110110110111101011011001111110001111101100000100;
#1 $display("%b", po);
# 1  pi=207'b101111001010101111101000101011010101101010111111101011001000001100111001010000110101001100010011011111011000000001110000001011000010001101110110101011111101001110100110010010010100001110110000000111000101011;
#1 $display("%b", po);
# 1  pi=207'b100101101110001000001011010110011100110111101110100101001000101101011110101011101101010110010000111101001101010011101000101111100101000001101010001001001100110110011101000010111000101000100100011110010001111;
#1 $display("%b", po);
# 1  pi=207'b111100010000110001000000000100001010010011000110010011110010011001111001011000011100000111101101011000011110010000110011111100000100110001011010001011110111101011000111110100111100101101011101111100100010101;
#1 $display("%b", po);
# 1  pi=207'b000111001100100110011011011101100011101101101010011110000000000010101001111100100100010110000011010100010110111101110001110101001001000011001100101111000011010001011100011001010001001110001001010001010101100;
#1 $display("%b", po);
# 1  pi=207'b101101100101111110111000110001001000101101101101110001000110000111111001010001000101000001100101100110111010101101101101100011110100001110011000001100000101100110001001001101010110101110110101000010101011000;
#1 $display("%b", po);
# 1  pi=207'b111000101111011101101111011011001110111110000101111111110100101101000101000011010100011011111000101010101101010011001001011100000001111101011000011100101011001111010011101111010000011010111011011100000101001;
#1 $display("%b", po);
# 1  pi=207'b100001101001100010101100001000001000110100000000000000111010101111001111011111000010000001000111110011001101100001101010001010010110110010100111110101100110100100001000000000011011000000011110100000000001000;
#1 $display("%b", po);
# 1  pi=207'b000100000101101010011011100000100101001100010001011000001011001011110101100010000000000011100111100110000010100011000011111110111010000011001011011101101110110101100001101110101000001000001011000001100000111;
#1 $display("%b", po);
# 1  pi=207'b000011101011101000000110100110010110110110000110101001101001010010000000110110011010001111110011110011101110000011010011010000101100011100110100010001000000110000010101111100000000101100101110100111101010000;
#1 $display("%b", po);
# 1  pi=207'b000000110111101000101011001111001111100100111001100100000101111111011100010010011001001011101101101101111001101110110110010001110011011100100111011000011101000011111000101100010001011111010110110100010111100;
#1 $display("%b", po);
# 1  pi=207'b111100110001100001100110111101000010100101001000100000000000001101010000000001110011100100001001011011010100010011000011111111110010000000100010010100011011110111101111110011001101001000010011101001100011101;
#1 $display("%b", po);
# 1  pi=207'b001000100101011000010000101000011101001111111101001100001000101100101010010001001010111111110000101101011010111100111110111111011010001010110001010010000000111010100101001011001101111011000001111110000100100;
#1 $display("%b", po);
# 1  pi=207'b101001101010110001000100000001110100011011111110000101010010110101011100011110011011100111111110111111010111000110000010010000110011010100001110110001000011100010011101000111101101010000110100010010011101110;
#1 $display("%b", po);
# 1  pi=207'b001110011010000110001000001110001011011101110011111100111011000110011010110100011001000001101110010101010100111110101111011111001101000111111101011111000011100010110100100100001100010001111000111011100001110;
#1 $display("%b", po);
# 1  pi=207'b011010111101011111010001001000000000110100001101111010011010110001000110011110010101110110010001111011111011101010000101100000111101001001111100101101010001011011101101101001011111010110110001100000000010010;
#1 $display("%b", po);
# 1  pi=207'b000110001001011000110101000110011100000001011001010111011001110001100110010101100101001111101100101000110000110010011010011110010100111001101101000001011000011011111000111101011111111100111100101101010100111;
#1 $display("%b", po);
# 1  pi=207'b100000101000000010100010000110100110111010011110010010101110101110000110011000100010111110111101010100010110111010001101000001101001001101110110001010111010100010001011011000110001010110011000101010100000101;
#1 $display("%b", po);
# 1  pi=207'b011110011000100000101101111010001001010111101111010100011000101000110101111101110101000110001011010111011111100001111010000100111000010101011001110000010011101110111111111110010110011001001001101010000001101;
#1 $display("%b", po);
# 1  pi=207'b001001111011110000010010111000111111101010101101001001001001000101100001101001111111101100101001001011001001001111011011010101001110110011110111110110000000010010100101010110110100101100010011111010001011011;
#1 $display("%b", po);
# 1  pi=207'b110001000010010010000100010101100110010100111010000000111000010011111010010110001111111101001110000111101001100100100011001100110011100100011100001010110110110100000010110011001011101000110101110101011000110;
#1 $display("%b", po);
# 1  pi=207'b100010101011100010110000011110001000111000110110101110001110100001111011001101100000010110100100110000111100010010111110110001001000010110101000110110010101110100110000000010010000110000110001001011010010110;
#1 $display("%b", po);
# 1  pi=207'b010010100101111001010011000010100011010110100111100101010000101000011101011001001100110111101111010100000110111101101001010001010010100010111010100000000001000011100110110011001111001001100110001011111001111;
#1 $display("%b", po);
# 1  pi=207'b100100111000001000000011111011001101101110110111011011001101101100110101101010001001001001100010011001011011000101110100110111001100100110111101111100110011000010110010111011111000111101111110100001100001110;
#1 $display("%b", po);
# 1  pi=207'b000101001000100110110001110111110000101111110011000010010001100010010111000111001110111111001110101111000001000101101011110101101111011000010100101110101010101000010010001010001001001010110001000000101010011;
#1 $display("%b", po);
# 1  pi=207'b110011011011010110101001011000011011010100001101011000110001111010101101100110101101111101010011011110111110110000001111101101101111011011110001011010111011111011110100111010111110010101000011011100111001100;
#1 $display("%b", po);
# 1  pi=207'b000010111100100110111100100100100010100001000100110100110110111110001101100111011011101100100011011101010001101110110011010101011011111001010100110010001000110011010010111010011100110010101001100011011011101;
#1 $display("%b", po);
# 1  pi=207'b110011011111011000101001110001011000011000000010000001111110101011000110110101110001001100110101011101001011010110011101001101000000110101001000000100000100000100011000110010011000101110010011010001000100000;
#1 $display("%b", po);
# 1  pi=207'b111010100111111010101000100001000100001011000011001111111100100001101010000101111110111010100111001110111100000010010000110000101111001000001111001011010011011010111101001110101011110110001110110111110111000;
#1 $display("%b", po);
# 1  pi=207'b101111000000101110010111101110101110010011111111011001000110101001010100111101001111101011001000100010011000101111011011111001100010111000111110010110011000100110010010011001011001101011011101110010111110100;
#1 $display("%b", po);
# 1  pi=207'b010011110000101001000010100111111111000110010101010110111001110110111111011111011010011111011111100000001110010000000011000011011101001010010010010110011111010100000100111000011101111100110000011110001001111;
#1 $display("%b", po);
# 1  pi=207'b111011110111001100000101101000111111110110000111101001111011110001000010010011111110011111101110011000001110000001001100000111101100010010100101000001000001100010011001110011110101100001001100010001000100011;
#1 $display("%b", po);
# 1  pi=207'b111001010110111011110000000110010001000111101011101111101100111111111100010010011001101100000001110011110100001001001011000000100111011101110100110110001001000010110110001101000101100001110000110100111111100;
#1 $display("%b", po);
# 1  pi=207'b111110001010000010110111111111011000100101000111011011110000101101010100001110100111100011100110000000011110111101110001101010100000010100100010011011000010100001000101010001111101101111001011111101010001000;
#1 $display("%b", po);
# 1  pi=207'b000001110111011011100000000000111100010010010011010000011101000110010100110101001001101001001000011010111001100110101010100100000110101111110110001100110111110100001100011001111100000101100001111110010111000;
#1 $display("%b", po);
# 1  pi=207'b101101011001001100100100000011011101100001000000110101101100001011101111010010001111010100010101010100011010101110010101001010000011010110110110000100011011110011000001010000101010000000110101010011010101100;
#1 $display("%b", po);
# 1  pi=207'b011101100100110111101100100100000011011110101100111011011110011110000000100001011000101111000001100101001101111011110100100010110100000100000001010010000111101111011110101011010000111100000100111010100101011;
#1 $display("%b", po);
# 1  pi=207'b010111010000010010111100001100000110011110101001110111100111010000111010101001010110011011100000001010111111100011101100110010001110011111100101011011011111010011011000110000110110110110110111101011010101011;
#1 $display("%b", po);
# 1  pi=207'b111000001011110010100101011100001111110110111110101010101011110110100000000000111101101111101000101100010001111010111100101001011001111010111111101111010011001101000101010001001011011100100100011100100101110;
#1 $display("%b", po);
# 1  pi=207'b001001111100100101110010000110001001100111110111010101101010100101000011100100100100011001110100000111101101000100010101010011010110011001111011010110011010010111001000011011011110001010000111111001110010001;
#1 $display("%b", po);
# 1  pi=207'b100001111100010001110011111011010110101110001110010101101101011100100101111000101111110111111011010000101010010001110011011100000100100011001010011001110001100000010010100111101101100001110110010001010100001;
#1 $display("%b", po);
# 1  pi=207'b100001110111110001101010001011000101000110000001111110011110100111011111101100101101001110011100010011111101001111010001101111110010111010000110011110001001101010101101000001101011001110000011101101111010110;
#1 $display("%b", po);
# 1  pi=207'b000110101100011100001010010001110001111000100001100001110001111101001001001110111011111100101111101100110000111000000001000000110100010100001111100000001110000100111101011001001110101000011011101010111111000;
#1 $display("%b", po);
# 1  pi=207'b100110010110100100010011010011111001010101000100000111000000110111101111001110000101100001001000011111001011000101111011010100100101011000100111101001100100000000010011010110010000100000111100100000100100111;
#1 $display("%b", po);
# 1  pi=207'b010111101001010001100011001011101100001000100010010101010000111000001101000111110011001000111000011010110101101000101101101101011011001111000101111101011100001110000011010010010011001011100011011100001110110;
#1 $display("%b", po);
# 1  pi=207'b010010010001000110100111100101000011011111001010000111011000100101010110110111010010011110100010011010100000111001100000010101001100001101011111111110110000010010010111001100011011111101101001001110100000011;
#1 $display("%b", po);
# 1  pi=207'b100011010110101110000110001101000011011010011011101100101010001001000111100100100100001010110010101011000111011000001011101110110000101111010001000010001001011000011011111100011000110001001100001001100111000;
#1 $display("%b", po);
# 1  pi=207'b100111010101111011111001100000101100111010100010110000111110011101001110100111111110001110000011000100111111000001110111110100110101110100101000010100011100010100011100000001001110011000001101001101010001001;
#1 $display("%b", po);
# 1  pi=207'b101100100011110110110011000100110011100010111000100011110110010000000011000101000110111001010111111111110101010111000001001110011100011101111011110001101001000010110111010110110101011010000111010011000101001;
#1 $display("%b", po);
# 1  pi=207'b110011101110111000111100100101011111001101010001111011010000111000110110111001101111011001111100101001001000111111101111010111111110000111111001001110100011100011100000111101001111001010011100000110000111001;
#1 $display("%b", po);
# 1  pi=207'b101110010001000011100111110001111001101001100101001001000011111000101111011010100001111111110111100011111010110001100110111011111001100101010111110111110111111001011110011001101010101101010101111100000111011;
#1 $display("%b", po);
# 1  pi=207'b111000111100111101010001011101111101000010011101110010101000111110110000000001011001011000100100110100001010101010001001000101011110011101110101011101111100111011010011100111010100010011011101011011001111001;
#1 $display("%b", po);
# 1  pi=207'b000110111011101101111000100000011001000111100011001001101111111010010011001111110111001111111101100110110011110010101110110110100100101111010010101100101101110001111011110110010110101110111111100111100000101;
#1 $display("%b", po);
# 1  pi=207'b111001100000000001001001000001001111111000011010010100111100101111010111010001111101100001001101111111101000000001100101110101010100100000001110110001000011001000001111010000100001001010111100011100000001001;
#1 $display("%b", po);
# 1  pi=207'b000111001000101111000011111010010010010000111100010010000101100100110000001101110010010000010010000011111010000001111110101100100010100100011101111100110101110111101011100111000010001111000001110010101010100;
#1 $display("%b", po);
# 1  pi=207'b110100001111010110000010010101111001111011100000110100001110100100000010101100100110101110000110011110111111011000101111100011111111111000100000001100100000001111010110001011011100101101011011010001111100101;
#1 $display("%b", po);
# 1  pi=207'b001001010011000010010010110101011101110010000000010100001100101000010000101101000111101111111101101010110011110001110111001100100010011101011010100101100100101111011000010000101110110001110101110011110010111;
#1 $display("%b", po);
# 1  pi=207'b111111110010101111011100001110110110000100001000010100100000100100001100011011110110000000100001010010111101001110011001001110111100001100110010000100001111000110100110111010001000000000000101100000100111100;
#1 $display("%b", po);
# 1  pi=207'b011011011010100110001011100100111110011000101001011011010010011110110111010111000110011001100111101010110010000101111101011110000111111110110000011100001100010000001110000100010010011101110010101011111100000;
#1 $display("%b", po);
# 1  pi=207'b011000111010001101100000110010101100100001111000001101010111011110011110111000100110111011111101000011010101010011111011110010111110111000011100010100011100100000111100101011000100110001001110010100110000100;
#1 $display("%b", po);
# 1  pi=207'b111001011101001110110101011010111011100111001111000010001101110111000110110110101111010110011111010111100100110110100001110011001011000110010000101000000011000110001110101011101001111111101100101000000011010;
#1 $display("%b", po);
# 1  pi=207'b011000011100011100110111101001110011111110101001100000110000111011010011111110001101100001101011011110001010011111000110111011000111001001000101101101000000110000100101110010000101110010111000101001111011110;
#1 $display("%b", po);
# 1  pi=207'b100110101000110111001001011010000100110010001011100111011110011101001001000011010110001101011111011101100010101011001010100100110111000000100010111101110000110011011100001011001010010010110111110000100000011;
#1 $display("%b", po);
# 1  pi=207'b011000001010000111101010011010011010110111110011100010101110010011000000011001000001010011100111000001001010110111101101001101000111010111111010000111010000101001011111101111011001110101000100001100010000110;
#1 $display("%b", po);
# 1  pi=207'b011101110011001111001010111000110001000010110010010110011111010110101000111100001110011010110011101010000101011011111100101000100010101111101010111001010101101001001101000101011100111010011111000110010110111;
#1 $display("%b", po);
# 1  pi=207'b000110011111110011001000100101110001101110010011001100011111110110011101000101101100010110010010100000100000011111000010001011011000101000100010000000011001111011110010000011001011110011011110101001011101111;
#1 $display("%b", po);
# 1  pi=207'b001100010001011001110000011010101011000111111101100101110011100000000110100000000001010101011000101010111011010010001101000000000011100001111010010010011010111000001000010111110011001000101110001110100111001;
#1 $display("%b", po);
# 1  pi=207'b010001011011011011100101011101000111111111010111010011110100100001000011111001000000111111101001111000010001011001100011011001010011001001010010100101010100010100001010111100011101111011011000011111100111010;
#1 $display("%b", po);
# 1  pi=207'b101011100011000111001101101011101110111111010101011011010100000010011001010011011100000110111000101111000110010100001110010111001101100111011111101001101011100000000011000010010110110001110010010011111011101;
#1 $display("%b", po);
# 1  pi=207'b011011001000101000110011100110011111011000011100100110011111100010011101111000101100011111011010101010011010100111111111111001101011100110111001111110111010010101010001000100100110111001111100010101001111010;
#1 $display("%b", po);
# 1  pi=207'b110100100010101111010101100110011000101111111001001100011111110101100101111110100011100000110101010110110100101000011001000100010000001110010100110010110111000000110001110010000101011010101000001100001110110;
#1 $display("%b", po);
# 1  pi=207'b111101111101110010101101010011000011111010110100100110111001101001111010000111011110101000100101100011101001001100011100011110100000111001000100001100001111010001000001001000000110110000100010010100011111001;
#1 $display("%b", po);
# 1  pi=207'b000111000110000010100100000101110000100010000011010100001000100011000000111011111100010101101111000100111101010101100011001101000001010100011000110101101101000111111010110000100100010100111101001110000110110;
#1 $display("%b", po);
# 1  pi=207'b111111110110111111100010111101001010100011001011101011110111111111111100000000000000010001101111010011001110101101000100011100100001010100101100100101011011011011010011010101010001111001000100110000011111001;
#1 $display("%b", po);
# 1  pi=207'b100100100110000110001011010100101011001101011101000010110011000110111111101110101000011011101010011101000110110011001001111100001111110001000011110010101011111001000111100111001001111101000101010100110011100;
#1 $display("%b", po);
# 1  pi=207'b001111100010101111100111011111011000110000011111110100011101011110000011010010010011010001011011010001101001101110010101100100110010100010101001100110010010101000111100110000110000010101001110001011010011000;
#1 $display("%b", po);
# 1  pi=207'b011011100111101010000110101110000110000001000010011001100011111110001111111111100000001011001100001011011101001011111110100111010111001111001000000111010000101100101101101011001101100011000100101101111111100;
#1 $display("%b", po);
# 1  pi=207'b001001100011001100100010111110110100110010001100010110011011000000111101100000110010001100010001010111001111110010100010111001011000110101111001111001101011110101101000110100110100010110011001000010000111111;
#1 $display("%b", po);
# 1  pi=207'b100000100011011000000000101000001011001001110101100010010111011101101110010000001001111110000100100000100001000100100001011010010011000010010111010001001010011101111100101010101101011011100100000111100010011;
#1 $display("%b", po);
# 1  pi=207'b011010011001110011000010000101100000000011110101001000101100111000100101010011001110000101111101010101101110010110000010000000101010101100110100111111110100011011010111011100110001101101110111110100111010010;
#1 $display("%b", po);
# 1  pi=207'b111011011001100010001010011101101101100011001011111000100100001100010100110111001100110101001001001000110100110001101001010110100001000011111101011100010000010010110100010110111110110101101001110111100101111;
#1 $display("%b", po);
# 1  pi=207'b110111001011110101110011000010111000111000111010110011111110010000000100001111100100000000110101010001101101111000100100101011110000101001001101001101110010101100011110111000001100010000111110110010111110101;
#1 $display("%b", po);
# 1  pi=207'b010111110000000010100110101011110110110100010010110101110111100010100101001111011011100001100001001100111101111011100000110001000100011010111100010011000001101010100110111011110000000001111111100110000000010;
#1 $display("%b", po);
# 1  pi=207'b000101110001101100101001011100011011001010110110010111111011110000111001110010011111111111010100101100111011100001110010011010001000010110000001001000000011101001011000100011111010101110101010010000000100011;
#1 $display("%b", po);
# 1  pi=207'b001110011011001101010010100110111110100010011110111101111001100011001001000111001010110111101110110000100011111100010001101111110001011010100001100011111000010100110011000011100000011111100100110000010001000;
#1 $display("%b", po);
# 1  pi=207'b111110110001100100110110010111000010100000011010110100000011100000100100001100001111111110010111010000100010000000100111100011111101000010001001111001010101000010110100100011100101110101100001001111001001110;
#1 $display("%b", po);
# 1  pi=207'b010100100110100011101010110101101100011111101001100011000111011111001111110000100101011101001100010111010001100110010100110000011000111101111011000110001011111001101101001011110010101110011011010000010000101;
#1 $display("%b", po);
# 1  pi=207'b001011000000000111100000111010000000000000110100011110111011011111000111011100110011100001011111001000110001000000010100100010000010010100111001100101001111010011100011110011011010011011001001100101100010101;
#1 $display("%b", po);
# 1  pi=207'b101001001110000001111010001011011111110111011101100010111110011000001000000100100111010101010101110111011000010010000000111010001101000111111001101000001001011110010101001100110100101001001010100100011111100;
#1 $display("%b", po);
# 1  pi=207'b100100000010100100110100100100111101001111011001001001010011111001011100111100101100100001110101110110011101111110111011100111100110101100101111110011101100011100100100011101101011111011011101010111011100110;
#1 $display("%b", po);
# 1  pi=207'b110000001100101011110010111110000111010011101111111001110111010011101110100100010110100011000101110000010001101000110111010101111111110000110101010101001100100000001011001111001011011101101000101011111111001;
#1 $display("%b", po);
# 1  pi=207'b001010000100110110110111011010010011011000001010001100110000111100011010011011010101011000100100110101010000011100001101000001001100100000110110110001111101010110011010000101001111100000001101000001100110100;
#1 $display("%b", po);
# 1  pi=207'b001001010001110100010000011101110100001110000010011100000001011001110100001111100001001110100011110101111111110110101110100011001111001100101011000101110000010000000110011000000000110111100010100101000011101;
#1 $display("%b", po);
# 1  pi=207'b000000100010001001111100101111011110000010111011101010001010001101011110101010000001110011101000000000110010100110111001001101010011000011101100001000011011111000110100001110001010100011111000110111010011100;
#1 $display("%b", po);
# 1  pi=207'b011110101111011110111101000010011010100001101000110011010001110101000011010100100011011101010001101010111110000111010111011110010011110010011100000110000000100100101010111111111101010010000001100001110110001;
#1 $display("%b", po);
# 1  pi=207'b001011000101101111011111001100100100001110011100101011100101001111010011000001001111001011101010110100010001111000101111101000000001001000000010111011100001010010110011000111111011000001011000000011010111110;
#1 $display("%b", po);
# 1  pi=207'b000111110101001110100010010000000001000001001101000001111011101101111001010010011001001011111110111010001010011010101000010011010101101000011100101100111001110111001110000001011111011011000010011011000100010;
#1 $display("%b", po);
# 1  pi=207'b001101011011001111111011011001111110000100011001000111111111011011110100010101101011010000110111011001010101101110100011001101101010000000011100010011010111101101011110010011100010011111011100110010011000011;
#1 $display("%b", po);
# 1  pi=207'b100010110011110110010110100000110100000011100011001110001001011101111000100000000001011110101010011101001000100101000000110111101001100110110000111111110000111100110111111101100010101010010000001101101001011;
#1 $display("%b", po);
# 1  pi=207'b100100001111011110101011010101001010001110110000110011000111111111100100110110101111111101101010011000111101111011000000010001010110101100001001001110100011010100001111011010011101000000011111101111100000001;
#1 $display("%b", po);
# 1  pi=207'b011010101111111101010111100001101001101110001110111100101101001100101101010100111001100101110100101001101100010111010101100001111001011101000100000011110001111000001101011110010100000000100101000001101010110;
#1 $display("%b", po);
# 1  pi=207'b100001010010101000101011110110010101010001011111001011011100011111110110100011111000011001000001001101001010110001100111011110100111101110010000101100101001001010100000011010111111000011001111000111000111010;
#1 $display("%b", po);
# 1  pi=207'b111111101010101110000110011001010110011001111101110111100000011001111100011000010011101101100010110010101010000110111010111001000100100001000000110001011010110110001011011000001010100110110101011101010101001;
#1 $display("%b", po);
# 1  pi=207'b100001000111001001111100011010111101100011001101110001000111110110010000111001111101101000110110000111100110011101100011000000011010010010011101010110011110111110000000111101101101111001100011010110010001101;
#1 $display("%b", po);
# 1  pi=207'b001000101101010001010000010010101011111011101011011001111111111010111001110110001011010101101011011110000100101100011011110101010111000011101110101001011011111010100101111110110001000110110101101110010010110;
#1 $display("%b", po);
# 1  pi=207'b000110100010100101011101011001011001101101100001110000010100000111100101000011111001010110101001100011010011010110011110101001110010110111001111001001110111001000011111101100111110100011101001111100000000001;
#1 $display("%b", po);
# 1  pi=207'b010011100100100011000000100111110010010011001000010110000011101100000100110110000101101100011001010101111110001111000111111011100111010011110100000011111000000011001011110010111100011101100010001001001001100;
#1 $display("%b", po);
# 1  pi=207'b101110000000010000100101110100101100010100101111010000101101000010111100000000101011110101101101001110100000110111000111000000111010111000111100111101100011000111011000000001010101000111101111111001001100011;
#1 $display("%b", po);
# 1  pi=207'b110101000001110111100100110000100010001001001101110011110110011100010010101110011010111001010110110110111110000001001101010101101100011101110000111010101011011001010011001001001000010011101001001000000110010;
#1 $display("%b", po);
# 1  pi=207'b011101100001000001100001110111100100011111011100110001010001000101110110111010110001010011111000101101111010000101110001000111010110000010110000011110000001000101011110101110000010100110110001011101110111000;
#1 $display("%b", po);
# 1  pi=207'b110101110100111101010111000101001101111011001111000110001000011110000111000010011101011111001100000001010100010100000101110011000110011000101100101111010111000001010110001010000011000101100100110110100000001;
#1 $display("%b", po);
# 1  pi=207'b010011001000111010100011010001011011001110100111101010011101101110011011001010011010000010011001000111010010110000111001100101100011101110111010100001100010111000011011011011100000011001011010000101110110001;
#1 $display("%b", po);
# 1  pi=207'b011010010111100011101011010110100111101100011001010000110101101011000000011100001100011111111000100110100111001001011111000100100010011100100011001011011100000010000010110010111111010011100010110011101000010;
#1 $display("%b", po);
# 1  pi=207'b010100111000010001111010100100010010001011110101011011011111000001001001110000100110011000101101111010000011010100110101001011001111100010110010100011111001110000110100001010111011000111001000101000101100101;
#1 $display("%b", po);
# 1  pi=207'b011101010010111111111000001000001100100011110110111111100111100100000101111100001001111111001011101101011111000010111111100001101011001110010010100011010011110011100011001100111110011111110000101011111101101;
#1 $display("%b", po);
# 1  pi=207'b000010011100001011010100110100010110100000101101101000010110101010101001111000101000001101101010111111001101001000101010111111110001101100100101110111011000001111111110101011101000110000100000100000101010111;
#1 $display("%b", po);
# 1  pi=207'b000100110001100011001111010101010000100000110111000111010010010111010111011110000001100111110100001001001011110110110110100111111111101101100010010010100110100001101111101000101110110111101101001100000101001;
#1 $display("%b", po);
# 1  pi=207'b000000010000111010011100110001110110110010100010001001111111011111100100000111111100001001101100000111101100110101101001100011100100100111010011110101101001110011001111100101101100100110000111100010000011011;
#1 $display("%b", po);
# 1  pi=207'b111000100011110011110100111001111110100001001101100001101001101001010011101011100110101010001111101010100101001100101010101001011101011100100001010011111010011010111111011001000001011001100010110010110011100;
#1 $display("%b", po);
# 1  pi=207'b010111000101101111010110010000100100000101010010011011101011001111110010100100100110000000000101111011111010101101100001111001001101100010110000110111010010011000110000111011110000000011101111100111000001001;
#1 $display("%b", po);
# 1  pi=207'b011000110111110011100111100001100101101001011100011100111000011010100101011100001110110101100000111101111101010011101011011010011101010011010010000001100101101110011101000000101110101011010010010101010100110;
#1 $display("%b", po);
# 1  pi=207'b011111110001011011011000010110011100100010101111001010001000111010010010001111010101000000111100110111000110000101100010000011010001010000000110100011101101101011110010000010100101110101111110101000000010010;
#1 $display("%b", po);
# 1  pi=207'b000011100001101110110001001000100001110010010110101111100011010110100100011011001100010100100010001100111010111111001011101100000001101011011101011100010110010111011101010010111000010111001001010011100101111;
#1 $display("%b", po);
# 1  pi=207'b000000001100100011101101010000000100101100010101011000100010011101100010110010110000001010011001101110100001000011010000101010000001010101110000110010101000110110001001000010100001001001000001110001111111111;
#1 $display("%b", po);
# 1  pi=207'b000000011011110000101000111011010110011010010111110010011010011010111000110111001000010001011011111010011100100011111111001110111001111001011000100101100000010110010001111001001010011010011111000011001111110;
#1 $display("%b", po);
# 1  pi=207'b100111011110010111011101011110001000010110011101010001101111111011011110100000000110010111111111011100110011010111010011111011101111101011100001011010000100110110111000101000111101000111100111001110100111011;
#1 $display("%b", po);
# 1  pi=207'b101101110010011110010010111101101101000000000001011001010000111110100011100101101100000000111011001100010100010000101000000100100000100001110011011010011110010101010110101010100010110011101101001010000111010;
#1 $display("%b", po);
# 1  pi=207'b110001100011101110001110100001101110011010110111001100110110101110011011101101100011110110011110001010010011010000101101110101111011011101011010101100101100111001111101110001000000001010100111100110110000100;
#1 $display("%b", po);
# 1  pi=207'b001100111011101011001010011110100010110111000101010000011110001010100010111010010000101001111011001010101110100100011000110111110000011111000110110011010101111001100001111101110110010110110111010010001110111;
#1 $display("%b", po);
# 1  pi=207'b111000011110111011100100100000010010001010101111100100111101010001111010011110101101100001011101001100110111001100101010001101001100011001101110101001100110111001111110001101101111010111110001101010001100101;
#1 $display("%b", po);
# 1  pi=207'b101010001100111100111111111101101100000000101011101000000111000011000110001010101111010011000000100101001111010101110000010001011000010111100111101100000001000110010101001001110001101110110101011010000000001;
#1 $display("%b", po);
# 1  pi=207'b101010110100100001111100111010111101000001101001111000100110110000010110010010110000000000101011000101011011011010000000100010001110010110101000001111000011111000011101010110000101010101011110100011101000011;
#1 $display("%b", po);
# 1  pi=207'b110010001111100001011111100111011001101100110111000011100100000111010100001101001010101011110001100110000001001011001000010000100011111011110111001110010011110111101001011111010101100100110110111010001100010;
#1 $display("%b", po);
# 1  pi=207'b001111100110110100110000010111000110001010010010010111101111111010111111111001011001101101100111011100000010001001011001001101100001000010011100100110001011010101100110010110010000101010110111100101001111010;
#1 $display("%b", po);
# 1  pi=207'b000111101011001101110010111011111110000110100111111111011010111010100000100010100010101111101011111010100001101110001010000000111000101010011101101011111110100010100100001110100111010001000101000111000011010;
#1 $display("%b", po);
# 1  pi=207'b110110111001111011111101111110100001111010001010101001010011110011111010010000011010001001011110110111100110111101010111100110000010011110001110010110111011010011111110001010100010001101110001000010110111000;
#1 $display("%b", po);
# 1  pi=207'b011101110011101111000001111110000110001000010111000000011100000101110110100111100010011100010000000001101111110100010100011100111000111000000011110100011010001000000010010000100100100001110010100111000111000;
#1 $display("%b", po);
# 1  pi=207'b100111011111111000110110100000100111110110101111100010001101000001010101111011001110010100111101101101001110111101110100010011001001001111111011000110110000100011111111110110100001010011101000111010101101110;
#1 $display("%b", po);
# 1  pi=207'b111001111111111001111000010010000000101111011110101011010000001001011001001100000110110010111100110000010011001011100011111111111011010000110010101011110011111111011101010101111110000010010000001000110101000;
#1 $display("%b", po);
# 1  pi=207'b110111111011011110001010110000010100101011110101010110101110111011010000011011000011011100101000011111100100010111110110000110101010000011100001000000101101001111101011000101010111001011011011110001000110001;
#1 $display("%b", po);
# 1  pi=207'b101010010101001001011000101001110101000011011001010011101111100110111010001000001110011001110110001101011100010111010000000001110111011010101110000101001100011100000111100010011000110110110000110010101111010;
#1 $display("%b", po);
# 1  pi=207'b001001001111000010100000101010011011110011111111010011000100100110001100101101010001110000100110011000010000101101111010111000011010100001101000000101001000111111110111000110000001110000000101011000101010110;
#1 $display("%b", po);
# 1  pi=207'b100111100001111111111011001100100100010001111100001010101011010101110001000110110010000111010000000110110011000110101010011101011011010010100110010000100001001101101001011000111101110001110101101001110100000;
#1 $display("%b", po);
# 1  pi=207'b100010001111000101100001111011010101101110100111111010011001000101001111010111011111111010001010011000111010000111110000000110000001110100011111010111111011010100100000010000100001101100011001001111100011001;
#1 $display("%b", po);
# 1  pi=207'b001101101101101010111111101001110101100011111111010001001010001110101000111001010011010011100100011111111100110111110101101101110001110110010010100001100001000101010010010101110001001100110100010011001110001;
#1 $display("%b", po);
# 1  pi=207'b110001111011000010101100010100010100000001110000010000010110010011010111011011100010101110101001101111100001110010101000010010001110100001110001100110000110001100111000000001011010100001100011101111000011011;
#1 $display("%b", po);
# 1  pi=207'b110001110010100001001110011000000110000100000111100111101101101111101101100011100010111000011111011001111101111101111001101010101100101001110111010010101101100110000010100100100101111101000110100000100011001;
#1 $display("%b", po);
# 1  pi=207'b111111101100011010100110000011010010000111101101101100101111110001111011110100001100011011111010011010010001111011001010001100000101110000110001000000111000101101110110100011110000011100000001001111000011100;
#1 $display("%b", po);
# 1  pi=207'b100000110000111110010100111110101101011110100000000111100100101000000011101110110111111100011111101001000000000100101000111011111010100110010011001010000101000111110101111100111101010011000011111001011010111;
#1 $display("%b", po);
# 1  pi=207'b001100101110000100001111011000101010111100010110001001101101000000110101000001001101011100101010000000100111000010101010101001101000001011111001100100010100011010011001100111100011011001100101101000011101000;
#1 $display("%b", po);
# 1  pi=207'b110111000001100110110011011001011111011010100001000101011110111101111010000101100100000100000111100010110001110011001100011001110000011001010011111100101101011110011100111010110010101101011101000001100000110;
#1 $display("%b", po);
# 1  pi=207'b110110001000010011110000110100011101000001011001101001100111101000001001011000011001011011101101100010011100001100011011101110110110011000000001100001010000111100001011000000000011111111111101101011011010110;
#1 $display("%b", po);
# 1  pi=207'b011010010100000010000010111011100101100110000111010101101000011101110111010011010101001100111000111101100101001001100100010100111100001110001110100111000101010110010111011010111001110011011100010010110110101;
#1 $display("%b", po);
# 1  pi=207'b100111001110011001111000000111001001111101000111101010011111110110110011111010011100010001100110010011011111011110000111110000101001111110000101001001111000100101100010010011110010100100000111000001110010001;
#1 $display("%b", po);
# 1  pi=207'b110010001001101000010101000001110110000111011100111111010100111111001100010011000100011100011010001011100010011001010011000111101001100000010011010110011011001110101110100010111010000010101110011101101011111;
#1 $display("%b", po);
# 1  pi=207'b101100100000010011011011100111101111110111011010111110101011000111011111001111010011001001001110110100111010001100111101010111100011010011111010110011111101101010111001001100101011010010011101001011111011101;
#1 $display("%b", po);
# 1  pi=207'b101111001000111010111111110010010011101011011110111010100000101000001011100100101111101001110011001010001101001011011000100100010001101011010000001100110111011000000100011100100010011010011000100011111010011;
#1 $display("%b", po);
# 1  pi=207'b101011111000110011001011001111100011101001111010001000111001011110110101110011110100010111100000110100111101001000011101110100100101110011001001111001111111101000011011110011110011010101000011011000000000001;
#1 $display("%b", po);
# 1  pi=207'b000011100101101010110110101001100000001011100100101001100110001101110010010010010001010001100100111100001010001111010001110010001100001000000011001101110110110000101101001101111010000001000100100010001010010;
#1 $display("%b", po);
# 1  pi=207'b100011111101111110111101010001001111011111101001000010001111001100010001001111001100100101000001001010110110110110100101100110101010001000010000101110101110000110000001101001110100100111011101010011111111000;
#1 $display("%b", po);
# 1  pi=207'b101000111110100000101100000010100011100000000000001101100110001100011100001011000010011101100110110100011111000010101110110110010101011111010101101010110100001000000010010101111100001111000100011101101110101;
#1 $display("%b", po);
# 1  pi=207'b110001101110011010001110110011101000001110100100000001110100011011000011111110011000101001011100111111001011101110110110111011110000010111111101110100110000010110101001011111010110101110011101111110101010011;
#1 $display("%b", po);
# 1  pi=207'b111000011101110000111000011101101011011111101001110101111100010000110011111101001101101110001001011001000010100001010110010000011101111010101111110110010011010000001101000111111010001111101011001111011010010;
#1 $display("%b", po);
# 1  pi=207'b001010101001100101011100000110110000101111101101111111001101000101011001110000110000101001100100110000011100100111111101111010011111111010011101100110100100010111001101000010111101011101010101001111011011111;
#1 $display("%b", po);
# 1  pi=207'b100101110100000010101101011110101010000100100011101100100001110011100001110001100000110000100101100100111010011101010111010100111000110001111101100001010000101111011110000100111000001010000011111010000100011;
#1 $display("%b", po);
# 1  pi=207'b110011001001010110001001010110111100010100001011100001000000110001001110001001011001001010101110111110011101001010111001001101100010100110011111000101011110001101111001100111011011001001101111010011001110100;
#1 $display("%b", po);
# 1  pi=207'b111011000100100101100001001001011011001010100100110000010000100001001101001100110110010010000000100000110010101010100101101101001111111110101000110111110011101000010101011001010011101011001111101101111101101;
#1 $display("%b", po);
# 1  pi=207'b100011011011110000111001110001001111110001100100000011000100110100010010011110010100100010010011001000110111001101011001100100011010100010010010111001011101111100001011010110000101000111000000001110110101111;
#1 $display("%b", po);
# 1  pi=207'b011100110000100001011111011001011000001100011010110111001001000100110111010001111000101000001001001011100001000101000101101111100110000011100101110110010100101000100000000110101110110100011100010101000000001;
#1 $display("%b", po);
# 1  pi=207'b100100100001001111101010000110101001000001111000011011011011011010010111101111101010001101010011101111001000110111111011111001011100101011111011101101010101101100100101111000101011101101000011010101110001100;
#1 $display("%b", po);
# 1  pi=207'b011110001010010100011001010010000001110001011100010000110010110001100011001010011101011110110011111101101010110101001010110111100000010101101000100100001000101100111010010000111111110101010010101101011101111;
#1 $display("%b", po);
# 1  pi=207'b111111000010100011101000011100010000100100010110000100110110100100001001001110001010001011111001000010000001010000000000111111101000110000111101000100110100100111010110110001110111100110110110100100100001111;
#1 $display("%b", po);
# 1  pi=207'b110010100110110011111010000111100110001110101001011001011011101100000001000001110100000000010010110111000101010001110110100100110001001001011110101010001101101101100111001100111011000111001111101000001101000;
#1 $display("%b", po);
# 1  pi=207'b101000011011001000111110000010001011010101001100001011100000011111101110100100101000100111011000110011001110101000001001101101110111010101001111011101001010110111100101000100011100100010011110010000111101010;
#1 $display("%b", po);
# 1  pi=207'b111000000101001101010110010000001000011101000010100110110011111101101000100011100101000001011011111000010010010110100110000101000110101100101011000100111110001110111110011000100111111100100100001110111001011;
#1 $display("%b", po);
# 1  pi=207'b100000001101111011001100000111101101010010011011010111101000111010000100011001111111011101110110111111100000001111110010111010100011100100000110110101011100100000110000010111000010100000000000101010111000010;
#1 $display("%b", po);
# 1  pi=207'b000011110110010011001010111101011001000011010111100010110111100000000100101111111110010100110000101101011000101101110111110101011000101101110100000111011000010100011100101100110000010001111011010110100101110;
#1 $display("%b", po);
# 1  pi=207'b111011010010111111111000001001000100110100000010110100011101000100010111110000101111110101011001101110110101100011010000001110100011011001000111000000001110001111011111000111100100010011010001000010111000000;
#1 $display("%b", po);
# 1  pi=207'b000100001111011110110010100101100010011001110000101000000100101001011111111110101001101011100011011001100100001000010001101000011100011100010000110001011100000100101110101010100010001101100101011010111110011;
#1 $display("%b", po);
# 1  pi=207'b111111000111000010100111010001101100010000101000111111100101111100000010011111000110001000011001010101000000111111011101011111101111111100000100100101101100110001100011001000000011010010100100001001101011101;
#1 $display("%b", po);
# 1  pi=207'b101001110000111011011001010110001000100011000100100010100001011001110100111011000100110100101110111000100011111100000010001101111100100010100101100110011110100011101011010110010000110010000110100111000100110;
#1 $display("%b", po);
# 1  pi=207'b000010000010111000100010101010110100011010001011100111101100100001101111100100110100100111011010001100001001010100110011000100011101001001001010101001111011001000111101011001000110111100011001111101010100001;
#1 $display("%b", po);
# 1  pi=207'b000000101110011111010011100111101011111010111101000111111110001101101001010001100001001111001100001010110100110101000101010110011101101110001010011001111100110011001100000010011001101010100001010111110101011;
#1 $display("%b", po);
# 1  pi=207'b011001111110001010111110001010011101111011100110011101001100100111011011011100111000000001000101010100011110100110110101111110111000100111011101111100010100011111001110010010111101110101101010101011000100100;
#1 $display("%b", po);
# 1  pi=207'b001110010110111100010010100000001010011010111000101100101011000110101011011100010101000100111000111111101110100010001101000011001100000110101000011111010100110111101001001010101100010001010011011010000000100;
#1 $display("%b", po);
# 1  pi=207'b001110000100000111011101000111111010111010001100101010111001101011001011000110111111111001000000100111010010010000000011011101110101011010100111011011001111010110111011011000001000111000110101011101001101110;
#1 $display("%b", po);
# 1  pi=207'b010111110011000111001111010011100011110111000100011110101100000101001011110101011001101010000010011100111011101101110100100001111110110001111101110100100001001101001000011111011000101101101100111011111100111;
#1 $display("%b", po);
# 1  pi=207'b111000101111011001010110110110000011010100101100001100011011001111011110101111011000001001101000010011100010000000100011111010110111011000111001011000000000010100100111000100010000100000010011001011010000001;
#1 $display("%b", po);
# 1  pi=207'b110110011000000110010011101010000111001011000011011010011001010100011111001110100111110111010111001010101010100001101110111100000010010011110100001110101010111001011100110100110111100001111001010100100100101;
#1 $display("%b", po);
# 1  pi=207'b011010101010101001111101111000101001101101011110110100111000001000000001010000000000100010100101100001001011011111001101100100100011010011110110110110101111110100010011110111111011111011111011110101110000110;
#1 $display("%b", po);
# 1  pi=207'b101100101010010100010011011011111111011101001001100110000111011001110111111111010111110010011100001110000011011010101101011001000010010110001100100000000111011100100010000011101111111100001001001100011111011;
#1 $display("%b", po);
# 1  pi=207'b010100000010100100010110101001101001001010101100000110000000000111110100110010111001101100010011100111000001001001001110111110011110100011001101010011000111100010010000111010101111011101101010110101000110111;
#1 $display("%b", po);
# 1  pi=207'b000100100001011001110100100110011011100010011100000101011100101100110000111101110101000000010011010110010111000000001111011001101111001011111000001010100011110010000100110100110000000010011111110111111001101;
#1 $display("%b", po);
# 1  pi=207'b110111110001001111111101100111010010111010001100110001000011000110100111100000010011000110011000000111101111101111100010111111100001100011101111111010110101000111001100111011000010010011001011010001111000011;
#1 $display("%b", po);
# 1  pi=207'b011111001001001100111010101000000100101101100100101100001110001100101100110111111010000001101101111100101100010101001110010110101010111000010011111100000011000000000000111111101110001000011001011011100101100;
#1 $display("%b", po);
# 1  pi=207'b000011111101110111101100100000101100110011001101010111111001111101111110011011000010100010010110000111001101100101011101000100111101111010110000110111011010000011010101000001111111100000100110101110110011100;
#1 $display("%b", po);
# 1  pi=207'b001011000000111001110111100100001010100100001111010010011011110100101111011100000011100101011011111000110010001001111101001011001010010001111100001010101110111111010001010000000111010010010010101010010010111;
#1 $display("%b", po);
# 1  pi=207'b100000100000110010001111000111001011100001110000001100011011101100010000010001001110011110111100000011000110110110110111011111101001111011111101101011100111111010001101100001100001101010101100110101000000100;
#1 $display("%b", po);
# 1  pi=207'b010001101010100011110110101001110101001011011000111101101000010000110000010100100000000111101000011100001111011011100011101010111111010010010101001111101010010110101010101001111100110100110011011101001011111;
#1 $display("%b", po);
# 1  pi=207'b011100110011010011111101111110101101111001100001100110010010110010000111001010111101011110101111111110100011101111101000101110100100000101011110101010010000100101110010100001111010001100111101111101010110000;
#1 $display("%b", po);
# 1  pi=207'b101010001111111100001010100111011010101111010011010111101011011100100111001110010111110010101101000001001101000001011111000110001001011101010111000100110100000011001001100100011110111001110011100101010111111;
#1 $display("%b", po);
# 1  pi=207'b101110000011010010101001111000010111000101010000011100100001100010010000001010010100000010101101001111000000010101001101111100000011100001101110100001010110100011000110110001110001011011111011001001110010010;
#1 $display("%b", po);
# 1  pi=207'b100111000011001001111000010000100100001100010011000000001110100011011011000011001000100001001000100101101101001110000010100001100011011000100011110100011010101111011001111000011001101111111010001110011000111;
#1 $display("%b", po);
# 1  pi=207'b111111111000010011010101101111111110011110101111000001111011010001000011101011110001110011110100001001111001100110101011101011110000010000111010011101111101011011110001110001110001110111110010100101110000001;
#1 $display("%b", po);
# 1  pi=207'b101110000111111011000011011000110100100001000000000101100001101000111000100010110100110100011101011100101101111010010111000010001011000001110111010001100010101100010000111010101001011111000111000010101010011;
#1 $display("%b", po);
# 1  pi=207'b101101111101000000000000001000011001111001011100001110000100000011000010111010001001101101110101101110010100011011110000111010100110100101010001100111101111001011011010000100111010000100010010010001010000011;
#1 $display("%b", po);
# 1  pi=207'b001111010100101101101111010111111001100101100110110111110101000011110111011001101111000001110110000001011010111111011101100000000111011010111111100100101010010111111100100100100111110001101010011011000000100;
#1 $display("%b", po);
# 1  pi=207'b011001011100010101010110101100111011100011000100010001010100000111000111000111010101100011111001000101100110110101011111000101000000011000111011111010110111110001101110101101000110010011001000010110011110100;
#1 $display("%b", po);
# 1  pi=207'b011011111000010000101101010101111110111101011111010110110100110011001001110001000111010101101110111010101100100001111001000101011110001000110100101011001001100000110010010111111001101001101100110101110001010;
#1 $display("%b", po);
# 1  pi=207'b000011101110100001111011001011011010011010101001111010111100100000110010111011100100110011010010010101000110111100110100000001100110011110110110111001111111100000011100010111110001000111011010100100000100111;
#1 $display("%b", po);
# 1  pi=207'b011111111100000111011110000110110110111110111010110111100101111011011011100000100111010100001000011001111001011100001111000010110100101110010101010011101000010010100100000101010100110100110111000011100111101;
#1 $display("%b", po);
# 1  pi=207'b111001001011001111111111010101101100010100011101010001011111000001000110000011101111011011010100000000011011110100101000010011011101101101001000111000101010011010100100001111000001111110011101001101100010000;
#1 $display("%b", po);
# 1  pi=207'b111110111111000101110001000100111010100110101000001001110100111111010111000101111011111110101000100111110111011001011011010011001101000110001010111110010101001011011100010101101000000110101011011110010011000;
#1 $display("%b", po);
# 1  pi=207'b100000011000010111111111001011101010011010100000000010001011000100101000110111111111011000101100001000011101000111111110110011010010000000100100100110011100010000100010101000000111010011111110001010011111101;
#1 $display("%b", po);
# 1  pi=207'b001001101001010011100000101000111000111010110111001011001010010011101011000000010100011111010000010110110001101111100011100100110001010010110011010101010110000101011111010000110001001011111000101111000100000;
#1 $display("%b", po);
# 1  pi=207'b111000101010111000000110011010111100110111111001111101011010001101101010111000011101101100010001100001011001100110110101101100101000100011110011001011010110000110000011000010001110110100010011010101110110010;
#1 $display("%b", po);
# 1  pi=207'b001100101101110000110111100000011010111110100110011010010100110100110010100111111011001100111010111100101110111000100010101101101011011010101101111110101101100101101101010101101111011011110010011100000110010;
#1 $display("%b", po);
# 1  pi=207'b101011010001101010001011001010001101001111111011001000111100000110100100111001010011100000010110101110000001001101000110010000010010111111101110110101000000101110111101010011010100001010100010011100001111000;
#1 $display("%b", po);
# 1  pi=207'b011110110111010010001000111110001101101001010010111100001011010100011011100010001101010101010100101001000001110111101100101101000000011110100100000100101010001111110011110101000000110111110100101110010100000;
#1 $display("%b", po);
# 1  pi=207'b111001010111010000101001111000101010101111010011100101010100110100111100111111100100111000000101101001010101110100000111100110000010001010110011100000011000100011010000100001111000010010100011011111111011101;
#1 $display("%b", po);
# 1  pi=207'b111000011000111100000011011111100010100101111101000010010010111101011100010101111001000001101111001001110011111110111010010010011000101000001101010000000001010011100011000101011011110101001010011001110110000;
#1 $display("%b", po);
# 1  pi=207'b000010010010101110110111000011000000010111000110000100001000001000110100011111110111101001011100011111111101010100110110010110110110001010111001011110100100001110101101010000111010100000000010001001011010000;
#1 $display("%b", po);
# 1  pi=207'b100010101100010100010001110000110000010110000001011110001111110010110100111000001101101100100010011110010010010110110010101000100101110010010111011000001101011100001000000100000010011001001111111101101111110;
#1 $display("%b", po);
# 1  pi=207'b001100100001010010000001101010010100000101111001010111100100111111000010111001101000111101011001000011000000000100100111100000000110010101011010011100001101111010010010001110100001001110111100000000110001101;
#1 $display("%b", po);
# 1  pi=207'b101011101011110110000000010110100110100011001000000111101111101100100111100010010001000101101001100110000101010010010000001111001111001010010010000101101000101100111111011010001100011110001100000000001111011;
#1 $display("%b", po);
# 1  pi=207'b010101010100101010010110000110000010111101001101110011101011101111110100000110011110110100001111011011000000010001010010101001110100010100011010100001011110001001110100110011101111011100010111010000010001001;
#1 $display("%b", po);
# 1  pi=207'b000000110001001100011110010100010000000011101000110010000101101100011111101010001100001100001101011111011101100010111101011011000011011101010010010100110101100111010010001111100101110100101000010101110110001;
#1 $display("%b", po);
# 1  pi=207'b011001100111101111110011111001111010000000111001100011011100001111001101000101100111000010100011100111010111001000010100010100110110110000001110110001011010101111111011010100000010101000001000000000001011101;
#1 $display("%b", po);
# 1  pi=207'b100101100010001001001111100111101110100111001001100010111010110000011100110110101111010011000000000111101100100001001110000011101010100101110000000110100111011100000011101101000101111010101111111111001001111;
#1 $display("%b", po);
# 1  pi=207'b011001011000101111101110010110001101011100111001100010111011110001000101111100100100100101110010011000101110100010100100100010001110100001010010011100101000101000001010101001100100001110000010110100100010110;
#1 $display("%b", po);
# 1  pi=207'b100001110000010000000010011111111100011011010101000100101101010100001100111011110000001001110011001101001111110111100101000001111000100100001110011111011100101000111110100101100001001100100010010110100100001;
#1 $display("%b", po);
# 1  pi=207'b000111010010100111000111110000001110001011010001111000011000100011011110010001010101000010110011011010000011111110100100000001010000101011111110110101110000110101100110110110000110000101010110010011010100010;
#1 $display("%b", po);
# 1  pi=207'b011110001100100000001100010010111101001000000000001010111010010110010110000100000011111110011100011001000010000101100000000011000001101101000110101001100100001110100110011100100100000011001101101011101001010;
#1 $display("%b", po);
# 1  pi=207'b110000100110011000100010100011111010100111010010101010010101010111100000000100001110000110001100011011010111011100000000100111111010001111110000110100111000111101101010100110011010011101000011000011110100001;
#1 $display("%b", po);
# 1  pi=207'b110000010011111011001001010011000100101100001011001000010111010100001001111110001010110110110110100000100010010011101000010010110010010110111100000100110111110010000100101011100001010011001110111100100001010;
#1 $display("%b", po);
# 1  pi=207'b101110100110001000110101000100001101000001110110011011001010101000111010000100001000101111000000110111000001001101000010111001000010111000111011111010000001100100010010100100010100011100011011001011111101100;
#1 $display("%b", po);
# 1  pi=207'b000111001001100001001010110000100000010110110010111101111100100000100110000001000110100011001111010010111011110001111010001010100010001110010100011010001101110101010011110010000000101001100100010111000101110;
#1 $display("%b", po);
# 1  pi=207'b010111100110001000100001110100010110010000100110110111000110100001100110010010000011101010010000001100111100100111000001001011101000110000111101000001000011101000101011110110101110001111100110001010011010100;
#1 $display("%b", po);
# 1  pi=207'b010011010110010000110000010001100001100010010100000101101111110010100001000001101011001100110000111001100111101100001100000010100110010011011001011101001110010010101100111101101000110010101111101111010000000;
#1 $display("%b", po);
# 1  pi=207'b000000100010110111110110000001101010000100101100011000111110000100101111100010010001100000000100001001011110000110110010110100000010110010011110100101100100110011100001011101100110111001000011011101001001101;
#1 $display("%b", po);
# 1  pi=207'b110011110000100100111000101110011001011100110110110000101100001011010101101101111011111110110000100101000000110000101101110011100001000111100010011111011011001000101101101001101010100000000110011111101000001;
#1 $display("%b", po);
# 1  pi=207'b101111100100010011110110011101001111101011001101110101000011011011101010100010000111001110110011011010110001101000100101001010110111111100101000110111100111110110010100000011010111000100011110000000100100001;
#1 $display("%b", po);
# 1  pi=207'b111100001000010111101001111100010010110110000000111001111100100101000011111010111001010101101100000101010011011101101101110010111001010111001111000000101001010100110011001111111100010100101001100100000101010;
#1 $display("%b", po);
# 1  pi=207'b011110110111010111011001101100011100111011011100100010001100010001000011010000001101001111110010011100100001101011111100101001111110000001001101010101100110001111110111000011000001110100111001000110011110010;
#1 $display("%b", po);
# 1  pi=207'b101010001000011100000100011001101000111011001111011100001110010111000001111111100010010001001111110101110011100110110110000100001110110100111110001000100100100100110000001111011110001111011111110111100000010;
#1 $display("%b", po);
# 1  pi=207'b011101110100001110001001101011100111110111110110101110101101011000001111010101110010101110111101100001010001110000111100100110010100101100110101111000001100100010011111100011010010111000001110000111001011101;
#1 $display("%b", po);
# 1  pi=207'b000111000011110011100101111011001101111000000001001110111001000011111101010010010111101001110110010101001100110111000100010100101000111100100001111000011001000011011010100001000110100111011111101111000001001;
#1 $display("%b", po);
# 1  pi=207'b011110001001100100000111000110101010110010100110110111110011000101001000000111110011100110101101010010101101010100101110000011000000110000000110000000101010001101110010111011111010100000111010110100110100000;
#1 $display("%b", po);
# 1  pi=207'b101100010001001011111000110000100101101001111010011010111001010001011001101010100111100000111110001000111111101100010110101100110101101101111110110101100000001000101111100100001011111101000000011101111110100;
#1 $display("%b", po);
# 1  pi=207'b100010010101111001110010000010111110001001111100011111101100111101110011010010111011101110111001111101100110000001110100011111110011001001101001000101010000100011111111111111011110111111101001111010010111110;
#1 $display("%b", po);
# 1  pi=207'b010110101111000111110100010110001111100001101001000111110110000000000110101100011010001100110001001011011110110000111000100010110100010001100111100101000000011110001111101010111111010110110001010100000111001;
#1 $display("%b", po);
# 1  pi=207'b111111100111101001110110111110110101111101111101111111000111101101000011111111000101101011110011000010111001101111011001000101101001100101100111101110011111110100000011001111011001111110100010110010000111101;
#1 $display("%b", po);
# 1  pi=207'b010000000010110011110110111001010100010111100001001001001100000100110000100111000001100101110110101010001111101011000101011010011100101100001100111100011000110011101101000011001110001100000011111000000000001;
#1 $display("%b", po);
# 1  pi=207'b101101000001100100110000110010011111000110010010111100111011010111100111110101111110011001100111000100010001001101001111010010011000110110110111101001010010100011010100100001010101100101101111101000111101111;
#1 $display("%b", po);
# 1  pi=207'b111110100111101111000100100100111000111111100011100111101111010100100000011111011011100001110010111001100111001010001011011010101010100000001101110001010001100001010001001000010101001101000000100110101000000;
#1 $display("%b", po);
# 1  pi=207'b000100001111110101110111011001010101001000011100110110111111110101111111010001010000011011000000001100110001001100100001111000111000101011101100001101011001111110011110110101111000010110000100100011100100111;
#1 $display("%b", po);
# 1  pi=207'b101000100110101000000000110101001100111110000010001000000001111000011101111000011010010000000000010001101110011111010101101001011001101010001001001001011011011111001011001101010010001110100001011110100001101;
#1 $display("%b", po);
# 1  pi=207'b010100011011011101000100011011111110010011000110100110011001101111001111101011111001110010101100001000110100011001101001111000111001110011111111010010100111000010111010100101111101000100010111010011101001011;
#1 $display("%b", po);
# 1  pi=207'b110111111111100110000110100111000100001010111100010111000100011111010111000101010010111101110101101110100011000010110101011011000001011001100101001101100101001110101100010010000000111100001001010111011110100;
#1 $display("%b", po);
# 1  pi=207'b100001011001001111010010110000000110101001110001001001010000111011010111001101010100111001111111000110110001000100100011111011110000111011011110000001001111101111111101101100110001001111000100111011101100000;
#1 $display("%b", po);
# 1  pi=207'b001101011111111100010001001010011101101100011100001110011011010011110000010011010100011001011011001110101100100100100101011100000001100000011101101000100101000000110000110111000000100001011111010010010011100;
#1 $display("%b", po);
# 1  pi=207'b100111100000111000000001111100101000101100011100000010110110001111001011000110001001000111100000100000100110010110101110110000011000111011000100000101100111010100100110111011010111110010110110111000101001001;
#1 $display("%b", po);
# 1  pi=207'b000001110101100000110101110011100011011001001110010010000110001000011000010110111110101011100101101001001100110010101001010011100100111111011100110111011101001100010011010001011110011010111110101001101110111;
#1 $display("%b", po);
# 1  pi=207'b011001001001110000111011001001101100001001001100001010001110110001011000100000110001110011011101101110111101010011111101001101100001100001001001101100100010111010101000101011001111000000101110111101011111011;
#1 $display("%b", po);
# 1  pi=207'b000111100110111010100110011010101100011111100111101010100111101110010011110111011110101101100101111010100101010010000100011000110110111101101010000010101011101111100000000110111010110001100000101000011000111;
#1 $display("%b", po);
# 1  pi=207'b010001110110011001001001000101100100010001100101000110101110100000001011100101110100011111011001110100000001101001010101110101101001111100010111001010100011111010111011010000011011010001010110100100110010101;
#1 $display("%b", po);
# 1  pi=207'b001001101111011011010110100010110001010001011111010001011011001001000001011001000101110101011011110010100110010101111101110110110011010011011100000101011111110101111001101100011000011100100011010110001000100;
#1 $display("%b", po);
# 1  pi=207'b001000011101011110101111110011010101101000100010001101111011100001000100000000011101011110101111011110100110001010111100100000010000001110100010101101011110011100011001110011000110011010100010011100011000001;
#1 $display("%b", po);
# 1  pi=207'b110010011010011000000111100010100111110110101100001010010011111110001000101000100000010111001110001100110101000110111010101010000100010100101011100001100010000111001001101110100111100100000101001011110110111;
#1 $display("%b", po);
# 1  pi=207'b011011110001000101001101100100101011100000010001000101101001100000111101100010011010011001001101100001110110100000011111111000010000000100000011101000011010100011000100111011010111001111101000011001001000100;
#1 $display("%b", po);
# 1  pi=207'b000001110001010100110001011110100110000011101101101011011111011111011010010000101000001100011100010101111011010100010101011110010011100111010000011110101110100100110111001111100010110101100101100001110011110;
#1 $display("%b", po);
# 1  pi=207'b000001010011101100111101110111011101000100101010100101100101101010001110110001000110011010110100010101101100011010100100001011111000111010101000010111001000110101110110001000111001011011011111001010010010100;
#1 $display("%b", po);
# 1  pi=207'b100000111001011001011100010111000101111101001100110111001010010110110000011000010110100110000000011010110110100010110011100000110010001001100000001001000100110100000101001000011011110000101011010100001101111;
#1 $display("%b", po);
# 1  pi=207'b001001010001011101101101111111110110100010110111110100101111101011101001101101001000111001101100010001110100100101001001110101100110110001001100110100100110001100011111110110011000010111011100111101001111100;
#1 $display("%b", po);
# 1  pi=207'b101011111100101010110100011110011110010111000101010000011010101001010011111010100010100110001010000101001000111011011111000110000111111001010100010001111010010011111000001000010001010011010001111100111001001;
#1 $display("%b", po);
# 1  pi=207'b010110111011101000001110011101001111011101101100100011101101100110110101110100010111010101001011101101000111110110010101010111101100110000111110000100100011010000001101000100011100100111000111100001000000010;
#1 $display("%b", po);
# 1  pi=207'b111011100011111010000001101011110100101110010000100111010000111010010100111111000101001100111110010011100001111111000010010011000000011100101000101010000001000011111111100111100010011101111011111010110011000;
#1 $display("%b", po);
# 1  pi=207'b010011110001000000011000100000010000011001101010110110110100010110101001010000100110010101111010001010101001000000101111110010100001111100100010110101100100011100010011110011001010000101001110111111110101001;
#1 $display("%b", po);
# 1  pi=207'b011010000111111001110011001001000010000010001011110011101111001001011101110111110000000101101001001011000110001011010101100011011010010101011101011110100011000101001110101100010010010000010100100100101001000;
#1 $display("%b", po);
# 1  pi=207'b101100001101101001101111100111001111100110101000011000010100001001011110001100011011100011110110010001001001111100010100101111110010001001001001101011011000001111111011010110101110110101000100001101011111100;
#1 $display("%b", po);
# 1  pi=207'b101001010110110001000010000011011110110000101100111011011100011010101010110011001110000001010101001101110111100011100101100100000111011001011111001010101110100101110010100110000011000000101010101001011111110;
#1 $display("%b", po);
# 1  pi=207'b110100001011101010000110000100101110000011001100110000101000101011010011001010000101100110111001001110111011111001101000101110010000000010111011111000011101001100111001101101101010111010111111011011100110101;
#1 $display("%b", po);
# 1  pi=207'b110110010011001100010100001101011001010011101101000010000010010110000001010110010111110111000110101101101111100110000001010101101000110100111001000100100000001011011101101111110110010001101111000100101101010;
#1 $display("%b", po);
# 1  pi=207'b000110001110010000101001100000000110101010000111010010000111100011110111001100010101000110100110010010110100110101010001000110101111011100000101000100110001110001100010001011011111100111111001111000110000101;
#1 $display("%b", po);
# 1  pi=207'b000101100010100101111100111011110001011010100110101100001001010111101101001010100111100011111010101001110010001110100101111010110110110001001011100011100101010100111000110110011000100110100001000010111110101;
#1 $display("%b", po);
# 1  pi=207'b110001110101111100010001001011110110111011100101011111001100101110110110000111101110011010001110000100101101001101100011010111110111111010111001011100111001001010010100110101011000100111010110010111110000101;
#1 $display("%b", po);
# 1  pi=207'b100111100000111101100111000110010100010101000101001110111010000010100010100010001011101001110001001101110101000010001111000010001011100001011111110100001000001000100100010100100010101110011110110011001100011;
#1 $display("%b", po);
# 1  pi=207'b101111100111010101100000111110001110010000110111001011111001111001010110100011111111001000011111011110101101000100110001111101100001100110101110000110001100110000101000001011111010111101011001100010000001010;
#1 $display("%b", po);
# 1  pi=207'b011001100110010101000111100011000010111000101100011101010111100011110111110000100011110110011001010100100010110011010001000000101100100010011001110110000110011011101110011110011110101100101011101100001101101;
#1 $display("%b", po);
# 1  pi=207'b101100010001010000101111010001011011111101000110110011100110100001101000000101001011111110010010111011110101110000001110001000001101110001101010011111000010100000001011100011111111010010000011100001111110110;
#1 $display("%b", po);
# 1  pi=207'b111111101001111010101000100011100100101010100011100000010100011111100111100001100001101001001010110001001000111001001011100111101111010100000111001111000000001001000110011110101111000010001111100011110110010;
#1 $display("%b", po);
# 1  pi=207'b100101100111111010011001100001100101011100000011010110000110101010001100010001101110110100111000100111011011111111111010000001011000100000000010011111111000101011001000101100011111001110100010000101101111011;
#1 $display("%b", po);
# 1  pi=207'b010100000010110111111001111101001101000001110010000011000100101001110001111010011000110011010000110010001011110000010100001111111001111110110111111000011100101011000010010101000001010111101000001010000111101;
#1 $display("%b", po);
# 1  pi=207'b110110111001100001101110110011100101101010011111001001010101010100100000001101111101001101010010110101010011111110110110010000111001110010001101011001110011010011111110111111011101101010110100001101010000110;
#1 $display("%b", po);
# 1  pi=207'b000100001010010111000011000000110010011010100010010010110011000010100001101110011101100000010000100011111010010001010000100111100010000011111101100010010100010101111111100010101100010111011110110111100111110;
#1 $display("%b", po);
# 1  pi=207'b001111011011001110100111000001101000011100011000010000001101101101110000110010001100110110101000110010010001000010100100011001110110010000010100111101101010101111000110110110100101011011010000100010101000010;
#1 $display("%b", po);
# 1  pi=207'b001011110000000101011101100010001011001110010110100000111001010110111001101000110010111011000011010010100001000000010000110111011111010110111010100000100100111101111011100111001000100111111001110000101111000;
#1 $display("%b", po);
# 1  pi=207'b001101111101100100101011000101111011001001111011100110000110111001011010011110101100001000010011101111101000000101110111000000010101111010110111110101100111010011000110101110101010100011010111011001111101001;
#1 $display("%b", po);
# 1  pi=207'b101100001000101111001011001011101011001011001001101111110110101000010100011010001000000111100100001100010110001001101110010111010101110001011101010001110010001110001101011010010101010011000101111000000000101;
#1 $display("%b", po);
# 1  pi=207'b111100100001110011010111101101010111111111101000110111110111011000001010011110000010010010110100000011101010000111110100010000001100000011111111101010100101100101110110110000101111010000010010010101011101101;
#1 $display("%b", po);
# 1  pi=207'b110000100110001010100001111111111101100011010111111101110101111110011110110011001011101001001100001111110001000001110011110001001111110111100000001111100000000001001111001111010110001100111111101010100011001;
#1 $display("%b", po);
# 1  pi=207'b000000001000111000001010111110101000010010011101100001000101011000100010010100011010010101000111010000010110100101111000110100100110110101110001110011100011000011110011100110111111011011000110000101100001001;
#1 $display("%b", po);
# 1  pi=207'b111101000100011011110100111011000100100111111111001110100001000000011001111000001001000000010101011110111001111110111111000100110001110000100000101011000001010000000101100100011100010110000001000000011100111;
#1 $display("%b", po);
# 1  pi=207'b101110000011000111011000011100000111011001111111011110101101110110101011111111110000010101010011001001001100101111101000010000001001111100100001010011001001101001000011000011000011001010011111011011110011000;
#1 $display("%b", po);
# 1  pi=207'b111101110011100100101011111001000000100001011101101100110011011010011110101000110101100101110110110111110110110111100011010110001100001010101001111101110010000100000010011111100101101100010001110011101111000;
#1 $display("%b", po);
# 1  pi=207'b110110110111010001010011110010100100000010000011001110111101101001000100100011110011101001111110100010011001100000011000101101110010111011001101011011101001011001100110000011011001111100010001111000110111110;
#1 $display("%b", po);
# 1  pi=207'b011010111011010000011100011110011100010101111000011101010010111111101010110001011101001111000011111110010101000101110001110000101001100000010111111111001010010111110111001101111001011110100110011101100100011;
#1 $display("%b", po);
# 1  pi=207'b001000100001111100011000011111001100111110110101010001100011000010101100001000000100000000111101001000011100100001010110111111010001001101011011001010110110110101111100000010001011001000001100110101111000101;
#1 $display("%b", po);
# 1  pi=207'b000111011011100011111100101100110101011010010011110111110111100101110101001011100101101010100110100101011001011100110111101100101110111111101000111110010101010000111110100100010001010111100011110110010001000;
#1 $display("%b", po);
# 1  pi=207'b111001100110101001010101001110010110010000010111110011100101110001111100001000000110101101000101100010001100000000011110110011111001111111000110111001100111000110110001100010000001101000000111010010011010110;
#1 $display("%b", po);
# 1  pi=207'b111000110011010011001111111000101111101100101111001011101001110101111000100111100010000101101010000100011110100011111110101010110101110101000101010011000011000110001010001011111111100101000011110100001000101;
#1 $display("%b", po);
# 1  pi=207'b110110001101000101010011110011001100000100101000010000010001111110000010110100010110011000001010010100011011101110111000110111111001111001010000001011111011010101100010001001000101100010100011010101010110000;
#1 $display("%b", po);
# 1  pi=207'b110001100011111010001100111010101000000001100111010101101011101001001110100101100000101001010110101000110110000101110110011001000010111001011100110010110011001101001110100111001110100010000111000001110001110;
#1 $display("%b", po);
# 1  pi=207'b110000101000100111011000111011011111011111111111010101000101001111000011110100011001011000011000100011010001010000101100101010111100110101111111000001010001001001010101110011010000011110000001011111011100011;
#1 $display("%b", po);
# 1  pi=207'b000000100101100101100110001111010001100100011001011010000110110010100110001110001011110001001010110110101101111110000000010010001001011001011100000000011110100010011101101011110100111011001011000011110000100;
#1 $display("%b", po);
# 1  pi=207'b111111011110110101011101100001111010111011100000001001001111100101001010110110011100000001010100101001000110111000011110001101000101101010101101111011000000101011001101111010110100000010100100001001000001000;
#1 $display("%b", po);
# 1  pi=207'b010011101010111000101010111100001111111101100100110000011001101101010110011101100001111001010001000001001000010011010000011100011010110101001110011001011101100111111000010010001000101011010100110000000100011;
#1 $display("%b", po);
# 1  pi=207'b011010011011101000001100011010001000001100100011110100101110001001101011011001011111101001110010110010110100101011010101011110011001010001010010110000101011000101011100101110101010010101100011011011111011101;
#1 $display("%b", po);
# 1  pi=207'b001111111100110100101011001110111010101001111101011000111100010110011011110100011000001110001110000110101001011000110111111011111101010010000011110011001001111001000001101110110010101000111100100101000010110;
#1 $display("%b", po);
# 1  pi=207'b011110000010010101001111100101000110010101101110000000010101110011001100111110010000010001110000001101011100110110101101001101001001111111100001101110001100101110000000100011000001110100000010000101100111100;
#1 $display("%b", po);
# 1  pi=207'b101011111010110111011110001011011110010011101111010000111101000110101100001010111100100000001010111101100011001001100110110010100100010101110010110000111100101001110001111001001100111110110100100001101010000;
#1 $display("%b", po);
# 1  pi=207'b001000000011010001110111010000100010100000101001111010100001100011101111011010011001000110011100000001000110010001111111000010110101010011110111001110100001000011101111111011011101100101100100101101110011111;
#1 $display("%b", po);
# 1  pi=207'b100001001010010010111011001101111000010101011111100010110010100010111100111011110100000111000101100100101100111011100101110101001100110011010011001101010011001101111100000100110011110001000000010101001110000;
#1 $display("%b", po);
# 1  pi=207'b100010101110101010111010000000011000110011011110101000111000000001111111000100101001100010100101110001110111010101001010111101101101001110000011010001101000011001110001101110010111100100000101111001100110001;
#1 $display("%b", po);
# 1  pi=207'b101000010000001011001011011100011111111111110101000110000000110111001110101101101010001111101111011111010110010101101011011100101111001101101001101011111000110010110111111001110000111100011101110110100011010;
#1 $display("%b", po);
# 1  pi=207'b111110001101110010010100001011110110111101000000000101111001000001010111110011110011010110010001100100100111110000011000010100100110111110010000111011111100000010010101111010111100010110000011101000101001111;
#1 $display("%b", po);
# 1  pi=207'b111110100100100001111101000110010000110111001101111111111101010011100000001011101010001000001001001110101101000100100001101010001111011100001110101001000100001111110010010011000000000110101101110111000111110;
#1 $display("%b", po);
# 1  pi=207'b001110100111111001100011011101000000101001011110010101100001000011110011000101010001011011110010110100011101101101000001011111101111101101011101111111110001101001010101101011001110000011001010001000011111001;
#1 $display("%b", po);
# 1  pi=207'b011111100101111010100111000100011011101111000000111010001111000000100001000101011110100100110000010100101101000110000111110000101010000011000100001101011011100111011110100110001101000100011101110101111100110;
#1 $display("%b", po);
# 1  pi=207'b010010000101111100000111000111100000110101111111111000011110101011100001000000001111010011010010100111110101100101000111000100101111101111111001001010011001000001101100110111010001100111000000101001100100101;
#1 $display("%b", po);
# 1  pi=207'b000101001011000000010101100110010011101100001011110011110111001110001111001001011100100001100011111011101111100001100011001010100011111111111101000001100000110010000101001111111001111101100110000100000100000;
#1 $display("%b", po);
# 1  pi=207'b100001000110010010101010001000111100101100110110001111101000101101010111011111100001001110101001101111011110010001111001011001011100001111101110010111010111100000000010000100000011010011111100110000111001001;
#1 $display("%b", po);
# 1  pi=207'b101011111111010100101011001111000111011111110001011101010101100010100111001000001010110111100111001100000101100010111010001000100100011100011111111001101101110011111010101100101100010001010011011111110101111;
#1 $display("%b", po);
# 1  pi=207'b000110100010100101011001010001111111111100011110100111001011000001101111000011110111110011011011000011011001010010111001000110000111100000000010110100001010110101001010111001100101001101001101110100111100011;
#1 $display("%b", po);
# 1  pi=207'b100000101111101100101000101110111001010110011100101010100110011000001110011000011111110110001011010110010001010111100101111111111110101000100010000000000011100010010000001111101001111110111100011001001111110;
#1 $display("%b", po);
# 1  pi=207'b010100011101010100010011000111011100101001000101111001011101001110111110011000101100111001111001100000111010111110000100001011010001011110010111011001110110001000111011000000011101001011010000010011000011100;
#1 $display("%b", po);
# 1  pi=207'b101110111001100011001010011100101110000110100110011111101110100010110110000110101101101111110110101111111000100110100011001001000000101100010001101111001110001010010001001010010011110100100111011001100111001;
#1 $display("%b", po);
# 1  pi=207'b111100101110010000101001111010011100110101001111101000001110011110010110010111111110011110011111101100101000000000100100001011111000001110000100000111110011111011111110101110111100010100010001010000000011101;
#1 $display("%b", po);
# 1  pi=207'b110011011011010010101010100111011000100110101110001111110011000001000001110110111100000001001001110011011001010000111110101010000110000011011001100100110111100101000100000100001011001001010111001101111000011;
#1 $display("%b", po);
# 1  pi=207'b000010101000110011000101110010000010000010101010111100111001010111111011000011001110110110011011101000111001001100111111100001000011111100001000100000101001001100001110000011000101011100111001010000000111000;
#1 $display("%b", po);
# 1  pi=207'b000100110111010111111110101001011100010101100010001011001100010110101010001011110000010100111001110001100101101001011001011011010010101110100101111111100011101010110011100011000011101100101111100011011100011;
#1 $display("%b", po);
# 1  pi=207'b111000011011010110001100011110101110000001010011001010001101000110100011101101001111010100000111100000101011000101010011110000011111000010110100011111011100110101000010101101010011111011101111111010100101001;
#1 $display("%b", po);
# 1  pi=207'b100110011011100000000101100101110100101110010111101011100000011000110111111100111001001010100111111101011101100001101000100001100000100101010100110100001100011011101110100111010111001000110111010010110010101;
#1 $display("%b", po);
# 1  pi=207'b000010010000101111100010001110000101010110010000101101010001110001110100100001011010101101011000010100001001011101101000000001110010011111111101010111010110100111011101000011110011110111011001110001101100110;
#1 $display("%b", po);
# 1  pi=207'b110010010110101100010000101011001100001011110101001010000101011010000101101010000001010011010010100001000101100100011100000111101111101101111110011000011111010010100111000011000110000111000001110101101001000;
#1 $display("%b", po);
# 1  pi=207'b011111110000101110110000110100110010001010010011001111110110010111011111111101100010110111110110001110000011000111110101101010011111000011011011100110101110101110010011100001001111000001010011001111011110111;
#1 $display("%b", po);
# 1  pi=207'b001110000010111011000010100001000011101000001011111010101100000110010100001101100101111011011100101001010001101001110100011101011100111011101000111101011100100100011000101011111101100010100111100100100100001;
#1 $display("%b", po);
# 1  pi=207'b001101000000000011000010111111001010111001010110111110001000010111110101101101000010010101111011001111000101011001010001010001001011000100001001000101001100111011001001111110000100011000100010101101101011111;
#1 $display("%b", po);
# 1  pi=207'b101000000001101111100101000000111100101100010011111001001011010011011111010011110000100100011101111111000000110001011000110000000001000111000000011001101001010011101100010100001010011001010000101011101010111;
#1 $display("%b", po);
# 1  pi=207'b111101111000101010101110010111000110011101010010100110100100100111000100111011010011000111111000110011101011111100101000011110110001111010001100010100010011011100011101000000101001001110101100010100010001101;
#1 $display("%b", po);
# 1  pi=207'b101000010001100000011010010100100101100001000111101100011110011100100110000100010001111111111111011101100000101101111001101111111001000001111110001010110010101111000011100010100110000101110000011001111000011;
#1 $display("%b", po);
# 1  pi=207'b000111000000110101011000001011011010011010000111111110001100100110000101000001100100010110001101111011110111000100010010001101000101100110000101010100001101000101010101010100100111000000000001001001100011111;
#1 $display("%b", po);
# 1  pi=207'b110001110000101001100010011001111001010011101011010100111111101111110000000001110100100110110101101100010101101001001100101111101101110100110010010001000000000011101100100000011011010000001111100110011010100;
#1 $display("%b", po);
# 1  pi=207'b011000100000000001110110000110001111001100011110100001000110111111001011001110110001110000010101001101100010000001000100110111101001100100001111011111101001000001110101011000101011100001111010000111010011000;
#1 $display("%b", po);
# 1  pi=207'b110010001110100010111100111110011110110100111010001101011001100100101000000110110000000100001011010011011110000110110011101010001011110010011001110111000010010101000110110110111001110010010110010101011101100;
#1 $display("%b", po);
# 1  pi=207'b111000101000001110101000001111100010101101100000111000110010010110001110110110000111101100111100110001101100101000011001010000110011100111000100110111000001111011111110111100011111011100010110010001101010001;
#1 $display("%b", po);
# 1  pi=207'b100000100110000110000000110101011010011010100111100110100100110010011001001100110000011010000001000110010010001011100101001110001001101110100110010010010110010110111111011010110001011101111111111101010000010;
#1 $display("%b", po);
# 1  pi=207'b111101100101010000001100010101010001101000001110100001001001100001110001111101010110001100111001011100111001110011011110000000001111101111010110110011010111111001100010110100001101101100011110011000110011110;
#1 $display("%b", po);
# 1  pi=207'b111101011100011110101110001011111011110000111000000001110001000101011011100011010100000100100110100111011100011110101111011001011100000011111010101111010000100010100110110101000111101111100001010110000001110;
#1 $display("%b", po);
# 1  pi=207'b001101111000111011101010011110001011001001000101111101010110100100111001101000100101101000110010000011100100001011011110010111001100110100111111110101110110111111110000001001110001000101010111110110111000000;
#1 $display("%b", po);
# 1  pi=207'b110000100101110001100101100001111000010010110101001101110100010011111010010111101110010110000100001001111011011001010101100111110001110011100111111010100101101011001000010101100100001101101000001001000100010;
#1 $display("%b", po);
# 1  pi=207'b110100001011100110011001001000111110110011010101001010110000101111110100010100101001000101010101100110000110011010111011110000111101000011011111100000001000101101010000010000111010001010001011100101000101001;
#1 $display("%b", po);
# 1  pi=207'b110101000000010111111110001100100011111011111110001010110100001110110100000110111100010001110111111001100010011011100111010110001011001000001110111101100001000010000011110111100001101101100001001010000111000;
#1 $display("%b", po);
# 1  pi=207'b111100101101011110001001011111010000011111010111000001000000110101011110101000010110001001000101000001001110000110011011010111011000000101111000100111001111101110111001011011001010111101100111111101011101001;
#1 $display("%b", po);
# 1  pi=207'b001100111000011100001010000100010001011010111101101011100111001010101011010110000001001001111001001101011101101110011100101001011101000000110001001101010110111111010101001011101001100010110100111100011111000;
#1 $display("%b", po);
# 1  pi=207'b100011100100100001011101000100001000101010000101100110010100010010000010001011101111111010010111011001111010011011110101010011010000101100000001100111101011010100100000111010111110001001110100000011110111000;
#1 $display("%b", po);
# 1  pi=207'b000100110000011101011101010000011100110110101001100111010011101011111111100111101111110101000111001101100101111010111111100011000110111000000011111111101001111101100010010101011110011010000101010100110110010;
#1 $display("%b", po);
# 1  pi=207'b000000111011011110011001100011010000000000101001101010000001111010100011000110001101011111100111000101100010100000011011011011001011110001001010000111111100011101010010011101110101001001000011101000111110101;
#1 $display("%b", po);
# 1  pi=207'b000011100010100011001100010110111011010010011111001010111011100001100101100110101000110010100110101110010101011011101110110011101011001000101001101010001101100100101110011111100001001110100000010001111000000;
#1 $display("%b", po);
# 1  pi=207'b000000001111011111111110110101001110000011100011001011011011001111111000001010100101111111010010000100100100100000001111110000101001110001110001110000001011101100001100000011111010010010011100011011001011000;
#1 $display("%b", po);
# 1  pi=207'b101100011000010101010010001111011100000101011010111001110000010110101110000011111111011011101101110110100011001011011111110000001000010110000011110111111001110100111101101111000100110110010100001110111010001;
#1 $display("%b", po);
# 1  pi=207'b010011110010100110001000110011001001001111010111110100011110001010000101101100000001110011100000101011111001101010110100001000110001001001010001010111000010110011111000110101010000011001011111010001101001000;
#1 $display("%b", po);
# 1  pi=207'b010011100111100101101101000001110000111111100000000010010110001001110100110111100110101111111101111001101000100100000110000011111001111010110000010110010001001011100000000011000011011011001101011110001101110;
#1 $display("%b", po);
# 1  pi=207'b110011110110101010111010101011001100000011100110000100111011110001011000011111101110000011111101010011011110010001111011110011111111101011101010010101110001111010010101011100110110100011011100111001110000111;
#1 $display("%b", po);
# 1  pi=207'b101001100101001011111001101011101010010110001100000100010101111011111111011010110011000010100101110010110001110100001110000110010110101101000011010001101110110101000111110110100111000110110101111010101011011;
#1 $display("%b", po);
# 1  pi=207'b001100101011010010010011100111111101110111101001000001110001011011101111000100000011010101010001101110001010111001111001101001001011111101010001011111110001110001010110101110110110011101011111111000001100000;
#1 $display("%b", po);
# 1  pi=207'b101110111011000100100110010100001011011100011011111001010110110011111000110111111100111100000111011000111110100110110101111011101010111100010011100110111110000100011001000111101000100110011000001010101000011;
#1 $display("%b", po);
# 1  pi=207'b001101100110010000101010111111000111000000111001110000101100010010000110000011111101100101001000100101001111110010110101101011100001110111100111111100110010011000111000011100110001101000010111000101001111100;
#1 $display("%b", po);
# 1  pi=207'b110110000011101110111011000001101110000111110000100011111001010010101011101101010010100101101011000011100111001100110110100110000011011111000110010100010001001011101111110101110101101000111001010000010011111;
#1 $display("%b", po);
# 1  pi=207'b001110011000010001110110100000001000100001111111101000001001010111001101110000001111000111101011011110100100101100010001100011000001000010011000011111110001110010101001001010100011111011101011101001000000110;
#1 $display("%b", po);
# 1  pi=207'b101011111010110110000001001100111111010000110110100101111001101000011010101010111111011001101011011011000101000010001011010001000111111111000100100011000100110110100010010111000011111110011010001010011111100;
#1 $display("%b", po);
# 1  pi=207'b111001000110101100100011000001000111000000111010011000000100011110011110011100010010110000011000011010111110101010100010001101100110001001100001010110010101111110000101100100101010110001011001000110001100010;
#1 $display("%b", po);
# 1  pi=207'b011010001000111000110101100001100100111111001000110111100011000011110100011100011101010011000110100000010100101011111001110110110101000111100011000110001011010110001001110100100111001000000111100000101011111;
#1 $display("%b", po);
# 1  pi=207'b101100011110110010010110001000110010011111111001011011101011001010001011001101101011101110110111010001100101011010100010111011011111111010011001000111010100110010001000000001111000111001001001011101000111100;
#1 $display("%b", po);
# 1  pi=207'b010000110100001001110100000110101010001100111010101000000101011001110111001110101001010101111000010010001101011000010010101001111101010110100111111101011010110100011110000001000111110010100011110000001100111;
#1 $display("%b", po);
# 1  pi=207'b010100110101110001000011010011110011111011101010110101110000101000110101111010111110011011100001011100100101111001111001101101101010010101011010000111001110110011011001000110010000101011110010101011001011001;
#1 $display("%b", po);
# 1  pi=207'b011100111111100000101010000111001011101011101000111011101111010100101011000100111110111110011110000000101101010100100100010101011111011000111101100011111000110100100110010011111010101111010001000010111101101;
#1 $display("%b", po);
# 1  pi=207'b100110100001101000100100110011101000000110101111101101010111010011100010100111101100011000110100111010000010101111110110110011001100111011010101010100001011010100100010111010100101101110101101001001001011100;
#1 $display("%b", po);
# 1  pi=207'b101111010110001100111000101111110000000100001100110001100110010000001111101110111010000110000100110011110010000010111111111000111100011101101000100001011010001101111100100001111010010010110111011100010011011;
#1 $display("%b", po);
# 1  pi=207'b010000111011110110111001001010001001000110010000011010100101000100110001000001100010100100111011010011101000001000000011011001001101010101001000010001101110100101100001101101011000101100101000100111110010001;
#1 $display("%b", po);
# 1  pi=207'b011100011000010111110000011100011010011101111110100011010001110001101001000000000011101010011100100110100000000100000000010001001010001110110011110000011110011100100110000101110001000000001011111111000110100;
#1 $display("%b", po);
# 1  pi=207'b101000010001000100111010010100001001000101101111101101100000110111011110001011101110000101101111110110001110001111001011001011010000001111010111111111101011100010111011010101111000011111110101101011110101010;
#1 $display("%b", po);
# 1  pi=207'b111000101011000101111110100010110011000101100110001110010110000110101101101001110101101001000000010101101011110101110100000001101111100110100111010100001001101011001011101100111101111111010010111011011000110;
#1 $display("%b", po);
# 1  pi=207'b100101110110101001010111000011101001010001101111010110011100000111111000100111010011110110010101100010110000111010000011111011010001111011101010010101000111010111001001010111011100001100011111100000110110000;
#1 $display("%b", po);
# 1  pi=207'b111000000001100100111001101010011111100100010001011101110010101001101101001001011111010101101011111110111111100011011100001111010011100101101101111111010011001110001110101100101010001010101000100100010011111;
#1 $display("%b", po);
# 1  pi=207'b101010110010110100101101100011011001100001010111001000101111101110111101010100010001110011010010110110110111000000100101100110110000111011001000101010100111000100111110010000111011101100101000111011011000000;
#1 $display("%b", po);
# 1  pi=207'b110100000010111101011111000011011011111110111100110001111110110101100101000101100010010111010011110011010000101110111001111111110000101000000100110010111100001001010001110101111111110100000101001011111110001;
#1 $display("%b", po);
# 1  pi=207'b111001101010011001000111011111110010010001010111011100010010000111001001100010010101110110010011001010000111010110110011111110101110010100011101101111101010001111001000010111000001111000010101001100111110001;
#1 $display("%b", po);
# 1  pi=207'b111100111000001000010010000110001100110010101000000000110000101101001110010110100010111001010000101011100110011011010111101010010111111000001011000011001110111111011101010011001110001101000100101011000010010;
#1 $display("%b", po);
# 1  pi=207'b100010000001111001111111010100000100000001000111110000010100110010100111110010000001111110010011001101101101101000010000001010111011100000110100101101011000001100101111001110010001010101101101010010011000001;
#1 $display("%b", po);
# 1  pi=207'b010111101111000111110000001100110010011101001011100110000001111101011100000000011010011111011000010011010111010011010111110000100110000111110001010011100111011000111001011100010000010011111110100110011100100;
#1 $display("%b", po);
# 1  pi=207'b110011100101011111110010111011001101011110101110001101101111100111110100111001001110001010100111101000101111111110100111111101110000011101000101110100111011011000001010100101101100011011111001011100100010000;
#1 $display("%b", po);
# 1  pi=207'b111011111001100010010010100100011001111010111111001000011101101000001011111000000101111110101010001100001001100110110000011101001000101000110110111000100011001110010010010011011001010011000101110011010010111;
#1 $display("%b", po);
# 1  pi=207'b010010010100011101010010111100011100100110110110000000010110011000011101110100101101010000000111000010110000101001001100101001110010111011000011111010010110110110110111110100001100010010001000001010001000110;
#1 $display("%b", po);
# 1  pi=207'b001110010011001101000010001001000111011001111110100111101110011100011110110101011011100101001010110001110010111011001111011010001010111001110100000001110011010100011000110100011100101011101101111110000100011;
#1 $display("%b", po);
# 1  pi=207'b111101011001100111110001111100001000110010001011011100011100000111001000000001110011010101111111001111011010000010101111111010111111001101010110101100011110011111101011110110011111110000110001001101000101001;
#1 $display("%b", po);
# 1  pi=207'b001110100010011000010100111110000111100111010101101111001111011111000111100100100101100100000100101010111001111110000111110100000111101111101010001010100010100110010100001101101100100010100101111111000010000;
#1 $display("%b", po);
# 1  pi=207'b111000110011010101101000001101011101000011001111010011100100100111011100100011100000000010101100000110100010111100100000001001111101000110010110001111100000100101011100111100101010000001100011000100101011111;
#1 $display("%b", po);
# 1  pi=207'b010010000001001011000110000010010100101001110011110111010100111001010011001010111111010000001111010111111111000010100111010101000010100100001111110010100101011110110111010011010110001011010001010110011001011;
#1 $display("%b", po);
# 1  pi=207'b110001101011111011011010111101101110101011101010001111101010111010011011111000110111011101000100101000011101001000110111111111000001001111110010111010010000100000101001011011101110001000100101001100111101110;
#1 $display("%b", po);
# 1  pi=207'b010101100111011111101111111111001000011111001010100111111101110001010000110000111011110101101110010111001100101011101101001100111110100101001000010001000001110111010011111110100011010010101101100011100110100;
#1 $display("%b", po);
# 1  pi=207'b001100101111011101010000011010010010111010100101011101110110000010100110000000111110010011110101101011101010011001011011100000000101011110010010111100011111101000110110010111111110011111110000000100111100010;
#1 $display("%b", po);
# 1  pi=207'b101001111110111010101000011110100011101101101000110110111101110010000100110001011010011010010011011000111011110101001011100001101101011001011110100001100000100011001000110010111100101101111110001001000110111;
#1 $display("%b", po);
# 1  pi=207'b001101100100010000111001011101011101010100001100000010110001000100110001011100100011000110100000111000001001101001011011110011111001101100011100000010101101000000101111101111100101010011110010000011101011111;
#1 $display("%b", po);
# 1  pi=207'b010100111001110000000110101010011010100100111100000000010110010101001001111100000101011110110101101010101011110011000110110101001001011110101110011011010101100001110101001001111111111010001110000010101011100;
#1 $display("%b", po);
# 1  pi=207'b101010010010111000001100101100001111111101000110111000000111011000011011000011010101000011010101111100110010000111011110000011110001110011001011110011110111000110000111010000100011100101101001000001000000000;
#1 $display("%b", po);
# 1  pi=207'b100011110101110100100101011111100011110111110001000000101001001001100000100011010011101111110110101110011100000000010110001101001110011001101100111110001111111010010110100011110101011001110100110101010101101;
#1 $display("%b", po);
# 1  pi=207'b010100110110001101110110110011011100111101110000111000001101010101110111101101111111010010011010001110111110001110001010001110011110010101001001010010001000001110011010001001001000110101010101000000000010111;
#1 $display("%b", po);
# 1  pi=207'b010110101010010001100000001011101110010010010011110000110110011000001011010101110101001111011110100001001100001111101100110000111111000011111100001010101011000111001011100000111011001000001110111100100101100;
#1 $display("%b", po);
# 1  pi=207'b110011100110001110111101011100101010100000000110000011100101010010011001001000011100000111110000010001110100100011000000100011001100000000100111110111010001000111110100011111001001101010111101101101111011010;
#1 $display("%b", po);
# 1  pi=207'b110100011000011110000110100101010110101001001111101111111111101110111000011100001001000110011101100110010000010110110001101111010000011000011111101110001011001100111001101010111010100001010110111111111111110;
#1 $display("%b", po);
# 1  pi=207'b100000111100001100110111001000011000001101010001010110101111110110000001100101001111100010101111110111101010011000010111010101010111110011011010001111000010111011001010000101001010010001101101100101110010011;
#1 $display("%b", po);
# 1  pi=207'b011100010111010110101110010101101010111101001001000111011001110010100010110101100000001110000111100111101110111110111110100101101100010111011010100001111100000000101010011011110001011001001000101111101010000;
#1 $display("%b", po);
# 1  pi=207'b101011101001111100010000110010010111100101111011111000000101110110001001011010101110001001011010000111100011100110100110000001000011000001010001100110101001010001110111111111000010100010101011000111111000010;
#1 $display("%b", po);
# 1  pi=207'b111110111000101000111011111111101100110100101101101000101111100110111001100000011110010010010001111000011111001111100111101010011110011100111001101001101001000101001010101011000011001100000001010010010110111;
#1 $display("%b", po);
# 1  pi=207'b111101010111100001110100010111111111000010011101110011111001001011001010001000000100111110010101001011100000010010110001111110100111010011100011101010000000001000111011100100011000111001010000101111100111011;
#1 $display("%b", po);
# 1  pi=207'b001111000010110001100111010000101000001000111010110001001110001101001000110100100101011101010001100000011111111010100010010111000110000101110111010100011110100011000111100000100110100110100110001010001010110;
#1 $display("%b", po);
# 1  pi=207'b100011010110100010110111000110000100010101001101100010010100111111100110110111110011011011011011010111011001010101010111011101010010111001011010110110110001101010100101101010110000001011111110011000010001110;
#1 $display("%b", po);
# 1  pi=207'b011101110101010110011101101011010110001111110100010100100110000100111000110111001000000101011001100100000000110100111111011010000101111000100000010100001110010101100111010100001100011110000010010101001011100;
#1 $display("%b", po);
# 1  pi=207'b110010101000010011100000010010011111110011011111011000001001001100001001011000000001100110000111110011001110101001011101111010111100101111000010010001011110101011000001111010110111111000010111011001001101001;
#1 $display("%b", po);
# 1  pi=207'b110100001010000001000011000100111111101111000101000111101010000001100101101000010000000011111001100100010011001111110011011001011000000100000001110001111001001111011001101101100000110011111011000000011111011;
#1 $display("%b", po);
# 1  pi=207'b010100110101111011111001100110001001110010001001001011100011100111101111000101110000100001001001101000101100110100101110101011010000001010100100101010001101100011100000110011101011111100001100111111011111010;
#1 $display("%b", po);
# 1  pi=207'b011011101000101001011111111010110001110010011001111101111111001010111100111001101101110001000001011010101011001001011001001100111001111001001010100001001000100101100100000000011111000101100010011011010000010;
#1 $display("%b", po);
# 1  pi=207'b100101011101100101000110111011110111110111110110100101010000011010100010000110100000011001000011000010011100000001110001000011001110111111011111111001100011011111010001011001010010000001011111010000110101101;
#1 $display("%b", po);
# 1  pi=207'b111010000100011111110101110100010000010111110001101110110010001011111001011110000010101011001000110011010000101111111101011100000110111101111100011001100011110111001110101011011000111100100000111111000001111;
#1 $display("%b", po);
# 1  pi=207'b100000101011110001010010101110111010101000011100011010001000000011010110011110110010101011110000001001111001001110101111000010100000110111111011100001111101110101000111110100111011110011000111001101011000000;
#1 $display("%b", po);
# 1  pi=207'b011010111110011000010011110101011100000101001001110110100010100001110101000011111110001110110100100010010110011100100001111100001111001101100101111110110100111000100001000011010001001100011000101100000101111;
#1 $display("%b", po);
# 1  pi=207'b000000010101110010000110000101101011000101000010111001000110001100010100110101010111001011000011011011100001101000010111111100001111101101000010110101000011110001111010010000101110001010110001110001010101011;
#1 $display("%b", po);
# 1  pi=207'b000111110011010011111111011110101001000101000011101000101111111010100101111111111011011011111110101001011011101011100101000100000101011110010110101010111111100100111100111111011110001100001000011101000000110;
#1 $display("%b", po);
# 1  pi=207'b001101101011010100001101100100100011111000110000101011111111000101000100111010111011000001110110000011101110010000000010100010110100100100001110011000101100011000000111111011011010111010110000001100001010011;
#1 $display("%b", po);
# 1  pi=207'b110000000110010000000010011010010010100010100001011101001010011001110011000001010100101010001001001010001011100110001110100111010111101100111110111101100001000100000100011000100110110100100111000111001001100;
#1 $display("%b", po);
# 1  pi=207'b010101000011100101011100110010010100001011000100111101111001011000001000110010111010101100001101100000111001100111110001101110101000100110100101101110010111001001110100001100111110101010111111001010001010100;
#1 $display("%b", po);
# 1  pi=207'b100011011100110001000100010000110101000010111101001011001110111011010010001110101101000100011100110100011000010010010100100100110110101110101100010100101011101100001000111100001000011011100000001000100100100;
#1 $display("%b", po);
# 1  pi=207'b100010110001001000111100100010100111000010000110011010000010001111011100011000100100001000010001001001001100111001101011111110100000100001101100111100111100101011110100011111011110101011110011100110101110110;
#1 $display("%b", po);
# 1  pi=207'b010110111010011010011010111111110100110100101011000101111111110000111010001000001111010111001101011000100101000101011100010100101010010100111100011011001000000011101101011010110101011000011101001100001111001;
#1 $display("%b", po);
# 1  pi=207'b000111111010110100010011111100101111101000100000001100000101011000111100110010010110000011011011011001100100111100101011010001101011110110101001100000010111101100101011011011001100010010011100011101111000101;
#1 $display("%b", po);
# 1  pi=207'b101101100000100101001100001110011011101110011110000001100011100101110000110001100010111110000011111000001010100000000010011011100101011000001110000011000000000110110100000100101110100111110000011100101001111;
#1 $display("%b", po);
# 1  pi=207'b100001101000110000101100101101110100100000111110001111010111011000110010000101101110111001011111000000101001110101100110000000111111011111111101001001100001000000001111000110111101011000011010011101100011111;
#1 $display("%b", po);
# 1  pi=207'b110100000100010101001111001101101111010100100101000011101010011110101110111111000011111110001110101000011110010010011000001001001100101001110111101010111111111110011110000111010010001000110010100110000011000;
#1 $display("%b", po);
# 1  pi=207'b100001111001011011110111011101010010011110111000100100011001001111101110001111000001111110111100101101111100011011100000111100111000000010000001111100110111001101100001001011110010101101111100001010000110111;
#1 $display("%b", po);
# 1  pi=207'b110000011000100011111101111010110110000111010111011011000010110001010100001111011100010110101000110000100001000011000101100001001011001010000010011110111101101001111010010110001101110011000100010000111100100;
#1 $display("%b", po);
# 1  pi=207'b000001110001000111110001100101011010001000010100111011010011100110111001010100100110001010011011011100001010010001110000000000100011110000101111000000001010010101001011101111010100101000110001100000000111101;
#1 $display("%b", po);
# 1  pi=207'b110001110101110101010011100110001010100101100011000111101100001011011010011001000110011111100111111000111001010111100011101100001110101111000110010101101101100001100010101101111011111111001101011100100000110;
#1 $display("%b", po);
# 1  pi=207'b111111010010101100100110101111001100000011000000100101101010001001011111010010011011100001010010100001000010101110100010011011000001111110101100101110001101011001101000101111000000100011011100000000000000100;
#1 $display("%b", po);
# 1  pi=207'b000111111000100111110001000001010011100110001111010110011011100110110011111110101111111101010101100011010010111001010101010110011011110101001101001001011001000011111100101000110011100101010100010010111111010;
#1 $display("%b", po);
# 1  pi=207'b110110100101110111100011010010111011110110100011001111011011100011010010111011000101110001100110111011010111011011101110000001110101100000101100010100010111011100010010100011110001000010100101101111101111001;
#1 $display("%b", po);
# 1  pi=207'b010101011010001011011110011001011101100101011101001111110000101101011000100001010110011101111110100110110111101000110011010101001001100101010000011011101101101011010001010010100111110100000010100001010110011;
#1 $display("%b", po);
# 1  pi=207'b001100101011001011110011111111110101011001000000111101110001000101100000101101100110000001111000001110110010111011111111101010111000001101000101111111101011111011111011110000100100010010010011011100101011100;
#1 $display("%b", po);
# 1  pi=207'b101011110001111111101000100000001100100010010100011100101111110010010101110010110110101101000110000110100111011111110100111111001100001110100000010111100010101010000000110100001100001100110001010110111101001;
#1 $display("%b", po);
# 1  pi=207'b011011010110110000001110001010111101111101110001000010011111110000100110101001101010100100110000110001000110010100110000111011010011011101101000101111000010011001000100111010111110001111110100000011111101101;
#1 $display("%b", po);
# 1  pi=207'b110011011101011011001110000111000010101010100111100111111100010000101101100000111011111000001100011100110000100111101011011101110111110010111000010001101110100011110111110111011010110010000110000110100111010;
#1 $display("%b", po);
# 1  pi=207'b000001001101000000000101000001100100011110010111111110100100010010001000000011011001101011011010001110110111011011110111000110100101010101111000110111011000011111110011001001001000010110101001011011001111010;
#1 $display("%b", po);
# 1  pi=207'b010000010110001101011010101001101100111101011101101000001011010110101100110111010111011011100010101010110011100101001010000111101001011111101001001101001101010011010001111011010010010110001100110010000001011;
#1 $display("%b", po);
# 1  pi=207'b011110000110010101100110011101110111010011001000100101011011001111100011111001010001011111010010101111011101111001110010111111001011010010111010011110110110100111110011011111011011011101110101100010000010111;
#1 $display("%b", po);
# 1  pi=207'b011110111000000111001011000100010110101110011100011111100101011111111100011010011011010001101010011101011111000010110011001111010110111001000110110110111111100111100010001100000010011000110101100100001110101;
#1 $display("%b", po);
# 1  pi=207'b110110110111101111001010110111010011101111101001111101000101110010100101010011001101010110011100001001000000001101111110001110011000100000011000010011101001101000111101011101000010101011101000001010011001010;
#1 $display("%b", po);
# 1  pi=207'b000010100010111001011100110011010100000011111010110100010010100001110100111001000100000001010111101101110101001010110100111000011011111000100000010000001111011100010110011110110101100010111101101110101111110;
#1 $display("%b", po);
# 1  pi=207'b001110101110100000011011010010011110111111000100100011110001011001010001100101011000000010111100000111111111001000110100111010101011000010010110011011101000111011011101001111110111000000111010110101001000000;
#1 $display("%b", po);
# 1  pi=207'b011111101000000001001100001100101100101010001101000100011100110110111010101100011001000101010010010100111011111011100011001001001110000110001111110100000001111010001101111010100011111011110100011011010101000;
#1 $display("%b", po);
# 1  pi=207'b000011111000101001000000000001110001110011010000110101101101010100111100001100100100110100010000101001001010001100111011111100101100110011101010000011010101010101111001000110100010111100100100100100111101001;
#1 $display("%b", po);
# 1  pi=207'b101010000010100100011111010011011111000011110101100010000011101111001100101100101110100010101010010000010000101001000101110110001010011011000111110001110000001100001110001101010011011011011010000011000010010;
#1 $display("%b", po);
# 1  pi=207'b101001101110110100000001010001000001110001100000010001010111100101111011101011011101101011011011011000111010110111110100000011000010101000101111101111011001000111101001100000110000000000100110000001100010100;
#1 $display("%b", po);
# 1  pi=207'b000001011110000010101001011111010001110111101111100110010101101100110100101111010000001110011010001001110100001101001001000101110011110101100111010100100110111010101100100111100100100010111001101011111110001;
#1 $display("%b", po);
# 1  pi=207'b101011010110010001000001110111011001101010111110100111100110000001001100011110010100010100110110001000100010001000010111101011011001001101100001111010010010000001111110111001001011000111000111110110001001110;
#1 $display("%b", po);
# 1  pi=207'b101000011110001101110001100000011001001010111100100100010100101000010111101111000010111101001111100011110000011100010011101010101100101111100011111011110000111110110000011001111010101100111011110010110000100;
#1 $display("%b", po);
# 1  pi=207'b000111111001100001010101110101000011100000001110101010111010111111111000101111111111101010010111101101001010000001111011110111101111110110011110100011000001010101000110100010001001010010001000101001111111100;
#1 $display("%b", po);
# 1  pi=207'b010000011111111000011110011110010011100111011000111110010001010101001100100100110011101110101011110001110110101010100111011001001101000000010001001100010110111100111101110011011110010010111101000111111011001;
#1 $display("%b", po);
# 1  pi=207'b000101000100111100111001011101000000010101100100100110111100111101111011100010100011100110100000001000011000100011100110100010100100100101000100100001001000101100000110111111010010011111111111100101111101110;
#1 $display("%b", po);
# 1  pi=207'b111001111110001110001001111101110001110101100010110100000001100110111010010100010010001111111010011000001101001101100001111100001000110000011111100100010101100101111100000101011001101110101100110100000101010;
#1 $display("%b", po);
# 1  pi=207'b000001001001110100110100000100011010100010111111000111111010010110100111111001110100010100011101011110101000000010000110100100100011000111000011110110010010111010000011111110000001000101110000100011111110111;
#1 $display("%b", po);
# 1  pi=207'b100011001000100010001001110001111001101010010001100001100100011111011100111011111100100010000100110000011111101101000101101100100110101010101100001010111001100110111000100010110101000011000110011101101010000;
#1 $display("%b", po);
# 1  pi=207'b111011000100110101001010101100011001011011011011010001000000100010001011101000111000010000101001010010111000100011100011110110101100111111011010101101001101010110011100000110010000101110001111010010110110011;
#1 $display("%b", po);
# 1  pi=207'b000111010010000110111100000101001001001000110000100111010010111101011000110001001001000000101010110010110101011111111101110110001011110101000011100010000010000110110100111011011000000110010100010001110110111;
#1 $display("%b", po);
# 1  pi=207'b011101111110101011101011100111001001000000100101000101101001111011011010110001010001011111110101010111000100011100111011011100010001111111100100100110110011101111111110110100100111010100110011001010001100100;
#1 $display("%b", po);
# 1  pi=207'b111001100110001101001011010100011011101101010100110011100111001110010011000101010000001110111100110110111010111001001110100010011011111110110011111110100001100101000111000001100000111010111000110111010111110;
#1 $display("%b", po);
# 1  pi=207'b001010111011001010101001000101000001011010100001111000001000101011011010101110100110110000010010111111100110110010010110001110101111111011000100101000101010110110011101101000101011001101011110101011110110110;
#1 $display("%b", po);
# 1  pi=207'b000110011011111100111011010011000001110001000110111011111110010100111011111110101010001110101010011101000011001010000111111000010101110101100000101111110111111000111000110001111110101110101011010111000001001;
#1 $display("%b", po);
# 1  pi=207'b000101101001010001011000101100110111001011001100111010010001011011101010101110100011000011111110010001010111110010110101000100010001110010001100101001111011000110000010101000011000110101010101011111010010110;
#1 $display("%b", po);
# 1  pi=207'b001001010011101011100010101111111010101110010010011110111001010001010001001000111111110100110101100011110011001100100000100001001100011000001011010110101000111011011010010101111001101000110101101110011111110;
#1 $display("%b", po);
# 1  pi=207'b001111000010101001111111100110101001000110010100001110000100010011100010111111100101110010001001110010110011011011101110010001010100000001101100011011000111110011011100001010001011111100001000110001001111000;
#1 $display("%b", po);
# 1  pi=207'b111011111001011000001001000111010100111110001010100101001100000101001000111001001000011110110000111011100000100010011111110101101000011011111000110100111101100101111111001100011010011100010100100110110100110;
#1 $display("%b", po);
# 1  pi=207'b110110001101000110100111111110101111010000100110110100010101111101000011101100111010001101110011111111100101001010100110000001100001110010101011100001101110100011100100011101000111110111001110010001100010001;
#1 $display("%b", po);
# 1  pi=207'b111010011000011000011110010111010110010011101010111111001111001000001111000001100100001100011011011101111011001101011101010110111101101000100001001000000110101101000110001100101101001000110010101011111111011;
#1 $display("%b", po);
# 1  pi=207'b111010100110110101111100000010011110100101101011101111010111010001111110100011110010000011001111010110011010110111111010011111001110100110111000111010001000011001010110010010101110011111010001010100010111011;
#1 $display("%b", po);
# 1  pi=207'b101111010101000000110110111110111001110110101111110111111001111010011011001001000000011000100000000011011110010101001110111010010101000010010011101100011010100101001111110101011111110001010010000001110010010;
#1 $display("%b", po);
# 1  pi=207'b101111010001011000101110001011101001100110000101110001111010011011001101100010010010100001011111111000101111010110000100111000101001110001101110110000101000011000110110000111000000110110111000111000011101010;
#1 $display("%b", po);
# 1  pi=207'b110100111100010001000101010010100011000010000011000011111111101010011011111100111111111110100101101010110011010110000010011010110101010001110011111001100011000010011111110001010001101110010011000111010000111;
#1 $display("%b", po);
# 1  pi=207'b001110000010011110101001000000011001111010110001001110011000001011000100100011101111001110010101010101011000111111110011110111100000110010101101100010110110000010010000110101100111110100001110011001100110101;
#1 $display("%b", po);
# 1  pi=207'b111100010101011101010000010000010111111101001011010010100000111010101000110100000110100001000001111101011000001010000000111001000111101100100101110001011111001110011100001100001011010110110101110111100110110;
#1 $display("%b", po);
# 1  pi=207'b000111010001010111010001100100010001100110010110111110101001011111001100111110100001000010000100011100011110010110111010100100010110110011000001011101101011101101111011001110101111010100111110110010110111001;
#1 $display("%b", po);
# 1  pi=207'b001111101001111010110110110100101110010111110110110101111001000101110000111000010101111000111111110001010010101000000110001000101000110000001000000110011100110000010101010000001011010011111010011011110010000;
#1 $display("%b", po);
# 1  pi=207'b110101111001011000101101100011010101001110010100001000100101110011100011011000011010101000000101010000111111011110111110101000101101000110010001101111001010101010110101011001010111110100110000100111000111010;
#1 $display("%b", po);
# 1  pi=207'b010001010111000110011111110010100100101101001110111100011111110010110011001101001100111000001110010000000101101110001110110101100001011110011100110011010111111111011101101001011111100000100111101011101001101;
#1 $display("%b", po);
# 1  pi=207'b010110111000011110100100100011100110011001001110110010101101001011101000101110100011111101100101001111001111110100000000000011100010100100001110101101100010101011001000111011010001011101010100110010000110110;
#1 $display("%b", po);
# 1  pi=207'b001011010100111011010100000111111001100001010110101000111001010100010000011010001000101000001101100010111110100100101001110100010100011101001011011100101010101101110011001111010000011001101010011010010010101;
#1 $display("%b", po);
# 1  pi=207'b110011010011011111011100110110011101001110010011100101100001100100000111100100101101101010001111110001100010011000010011000111010010100000111110010010110001100011011010001101000011010000011000001000010101011;
#1 $display("%b", po);
# 1  pi=207'b100111011110100110111101111111110101101000101100000000100100101010101111011111011001100100001000101010000100000110011000101011111010110110111010000010111101011000110000011110111010100000001110010000111101110;
#1 $display("%b", po);
# 1  pi=207'b010010110010100001101100110000110110111110101000111110101001101101000011111110000110101000111111011010101010010001110111011100010100111110110011001010101000000010001011010000001011110101111101010000110111100;
#1 $display("%b", po);
# 1  pi=207'b000111001011010100101100011011010011110011101010111011011110101010100001101010000111001000110101010101010110101100110110011111011100110001110000011010000000101011101010000010101000101100101010111000111011010;
#1 $display("%b", po);
# 1  pi=207'b001100101001011001010011011011010000011101010010011100000001000100011011011000000110110011000010110111100111000111111111100101000011010010011001001000001001100110011000010111110100111011001111010110110101110;
#1 $display("%b", po);
# 1  pi=207'b010110000110101100101010000000111101111110010010001111101111101111111010011101111110011100000110100000001111110100111001110101001000000000011101101011011110101001000000001001100010100001110011011101100001101;
#1 $display("%b", po);
# 1  pi=207'b001100111110100101001101010100000111100001110100101000000011011101001111100101000111110110010011011010000011101001110110110011100111000101100011001101110011011111101100001100110000100000010110010111010111111;
#1 $display("%b", po);
# 1  pi=207'b011000101011001111010010101101000011110001101110001001010111001111010001000010101001101000101000011010100110101110101011001111100101111110100000010111111100101011111000111000011100000011110010101110110011111;
#1 $display("%b", po);
# 1  pi=207'b101101010001000111011000000101111010011011001110101011111100010010100100001011110011010111011000110101100011010100000101000011101100110000101110000001111010111100110001011100111011011011011101000001001110010;
#1 $display("%b", po);
# 1  pi=207'b100001001001100111000010111100100011000000011101111110101101100101111000110011001011011100110010110111111101001111000101011100011011111101111101101011010100101001110101101110010001111100110100011101010010011;
#1 $display("%b", po);
# 1  pi=207'b010000010001110000110000101011111110101010010011110010000110000101111111000000011010011111000101000110101000001101101110101101100100010110010100011100000100001011101011010011000100110001110001000010010011101;
#1 $display("%b", po);
# 1  pi=207'b111101011000000100101110011000100100001101100110011111111100011110001011000001111011011110010010000011011100010010011111101111101110000101111001000001111000001011010001110110100011011110110001011110100101011;
#1 $display("%b", po);
# 1  pi=207'b100000101010111100111000110100110010011100000100000001000111000110100110111111000101000111101111010111101111110110111000111011110100110001111111010110000011011101110111100000011101111110000011110011111100110;
#1 $display("%b", po);
# 1  pi=207'b101111010101110111110111110000110001110001001111000101110100000000100001101010110010011110001011010010000100110011111100110010110100000100111010111110010001011001101010010110001000010000100111110110110011101;
#1 $display("%b", po);
# 1  pi=207'b110110111110000001010100000001001011000001010110011000010101001010011001110000000100000011101010011101100001010100101111100111111000000001010000000000111110100011100000100101000101100110101011011001110110011;
#1 $display("%b", po);
# 1  pi=207'b010000110001010001011101101001010001011011001101111001110011111010111000000010011110100011111100001000000111010000101000011000010010010111000001001111000000111010010010101100111111111011010000100011110010111;
#1 $display("%b", po);
# 1  pi=207'b100001011010001001100010111111111010101001010001100011011100001111111110110001110101010000000010110100111000100000010000010101001100010000001100100001010001110001101100111101011010010001110100000011111100011;
#1 $display("%b", po);
# 1  pi=207'b000001000111001100111111101011000001001110110110110111100110110011110001110010101100011101001101000110000010000111110100010110000010111100100001000011101111101111111001101100010010101100100011001011110001011;
#1 $display("%b", po);
# 1  pi=207'b001000101011011010101000101111100000000100011011110000111100010110101001111111000100010000100110001111100110010110010101100011010010010011000001010111000000000001110000111101001001100111110000001101000000101;
#1 $display("%b", po);
# 1  pi=207'b110110011110111100010011011011100110101110100011010000110000111110111010101001100110011100011011110001111010000101111111001011010010011111100100111101000011111001101010101100010001100110101110011010110100100;
#1 $display("%b", po);
# 1  pi=207'b000111100000000110111101110101110100100001001011001011111011101010110010110000001110000110001101101011001110100011100111000110111001111000111111011101011100111101110111001100101010101010011100001001100110111;
#1 $display("%b", po);
# 1  pi=207'b100001101100100100100011011001010111111111100100110010011101000000100011101011100011001011101110111011110010100111110000100111011100010011000010111100010000101111011000101001110101011000110101011101011010011;
#1 $display("%b", po);
# 1  pi=207'b110101111101010010010100111111010010011101100001111111101101100011110100110001000000111100111101110000001100000010101101011101101001111100110011000111100110000110111000101001111100100101110100011100100100101;
#1 $display("%b", po);
# 1  pi=207'b000110000000000001011101100011100100100001101111000010001001010010110000010100110100000101010110110001001011111101100110100011111101100101100110100010001001100110001101001011101001001100111011001100010001001;
#1 $display("%b", po);
# 1  pi=207'b110110011100101101100011010000011110000000101110100011101111000111111100010111110111101101000110011101110000100010111001100011101110000100010000001100011000100011000111111011101100010101100000001011010111010;
#1 $display("%b", po);
# 1  pi=207'b111100110100010110011011110010011001110101010010010111110111101001000101100110011011101100100110001110011111101001100001100101010100101111110110101110000101100001001011011001111010010101111101000110101110011;
#1 $display("%b", po);
# 1  pi=207'b100000101000010010101101000101111110100011011111100010011100000111010011100001111111101111111010001010001111111010011111001101100110110100110110001000000010001010110110111010000110111011110010101010110000000;
#1 $display("%b", po);
# 1  pi=207'b001011111000000101111101100111011010000100100100100001100100011110000010001011111110001100100100010001001111110010101100100110000001111000001100001011010100110011101011011110000001110010010101100010010001001;
#1 $display("%b", po);
# 1  pi=207'b100101000111111111001101111101011110111010101111011011101100001110100101101011111111011000000000101100100000010010000111011111001100011001001010101111000000111100100000000100010011001001110000110011010101000;
#1 $display("%b", po);
# 1  pi=207'b000101111000101101000001100011001111101000010101101000011100101110101011011101111101110101111101000011111010101000101000100111101011100011100110010000110110000001100011011100111011001001001111111111001011000;
#1 $display("%b", po);
# 1  pi=207'b110011101111111100111111001010101111111111001101010110101101011000010101110010010000110011111011111101101101101101000000010001010011101001001100110101001101100101000101010100001010100000101101011100100110101;
#1 $display("%b", po);
# 1  pi=207'b010111100101011010010010010111100110101110111111000000110100010101110110111101001000101000000000101111011110110001011011001100000110110000101100101110010101011011010011001111111100110011001111100001000000011;
#1 $display("%b", po);
# 1  pi=207'b000100001011011000110110111011101111110001011010010001010010010010100010110110010110001110011110101011111110010010000111011100111110000001011101110101111101011011001110011011100001110101100011111010011101000;
#1 $display("%b", po);
# 1  pi=207'b110000100111100110011000000000001100111100111000101110110100010101000110010111000100111000011001100101000001000000010010011111010100110101000010100110000101000000111110100001100010000101001000100111100001000;
#1 $display("%b", po);
# 1  pi=207'b110111111001110111000100001001011011111011110000001011011000000110010110010011011100010001110111110101000000010101110010100000000110101101011011000010010101011111110110100011001000000100011110111000101100111;
#1 $display("%b", po);
# 1  pi=207'b010001011111100111110001011100100111011000011110100101110110000110000011000110111010000110111110001011101011101001011100110101101001110011001011011110110110001011001101001000010001000111001000011110001001100;
#1 $display("%b", po);
# 1  pi=207'b111000010100010100000100010011001001100101000011111010111111000101001110011110011101000000110001100101100110111111011010100110101101111110000101111010010010010010011101000101001100101000000001101100010110110;
#1 $display("%b", po);
# 1  pi=207'b111011000101101111100000011100100100110011100000001001001111010000000011001110100001000111111000010111001011101011001100101111101010000000001111111111010011010001011111011001010101111111100000111001100010100;
#1 $display("%b", po);
# 1  pi=207'b011111111110110010001100010110100000001000010101110001011010110101100101111010010001110001111000101011001110010100010110001010100000000100000000011101100100000000000111001100011011000111101101100010100001010;
#1 $display("%b", po);
# 1  pi=207'b100111011101010111001000010000100111010110101110000110100011100000001011010010000011000000011000100111000011011011010110010000000110110111000100110111010101111010001100110101011100110011000110001001010001111;
#1 $display("%b", po);
# 1  pi=207'b110111111010011011110011010110010001011100111001011101011100001110100000110000100011011101011101001111110001110101110100101001110110101111001101011001100001110110011010110001010000000011001111011010011101110;
#1 $display("%b", po);
# 1  pi=207'b001100110000111010001110011010101000010111011010100000101111110011001010100101011100000011001011010000111011011010000010001000100011111001000000011011100000001010010100101010110111000110010010101110100100010;
#1 $display("%b", po);
# 1  pi=207'b010101110100010110101111011100110011111000100111111111010001101000000100110101000000011011000110000100111110010011001100001011010110000110111010110000110111101100001110101000101001000000101010000111000110001;
#1 $display("%b", po);
# 1  pi=207'b000001011100001101110000001101110010000010110101001010000000010110111000100100111000101001111110111110111100010101001111110010000110000101010001100010011111101001010110111010000011001101111111110111100000000;
#1 $display("%b", po);
# 1  pi=207'b011110000101101101000101010011010000110010011010000001111100110000111101001101110010010000011111011000000110101100001001110100011011110010110110101100110001101100100001011110000011101111111000101000111001011;
#1 $display("%b", po);
# 1  pi=207'b001110111110110101110001011110011100100001110110111010110111100010110001000100100000000111110001110110010000000100110110010100110111010111011000010110011011110000001011001110100000011010000101011110011001101;
#1 $display("%b", po);
# 1  pi=207'b010101001101010100000011010111011100100000001010100111110010110010110010100000011111000100000000010110010101010101101000110011110101110110000001001000001001011110010100110101101000010100110100101010000011101;
#1 $display("%b", po);
# 1  pi=207'b111101111011010100000101101110010011101111011101110000111101011111110011100100110101010010100110100110011011111100011001010111010000011111101111001110010010100100000010101001010100111110001101000111110100110;
#1 $display("%b", po);
# 1  pi=207'b000111110001111101011110011010000001011101000100010111010001010110011101110010100101011110010010010111110101111100100110000000100111000010011111110111110100100010111011011010000011111100101001010010001111100;
#1 $display("%b", po);
# 1  pi=207'b100111110010110001111010000101110110100101010110110111100000111000111111000010000101100000100100110110111011101111011010100000110001000101110001110100100101010000011100111000100000110111100101111101100111011;
#1 $display("%b", po);
# 1  pi=207'b001111001000010011111101111010100011000010011001010101010111011110000101100011111011001000101110101001010001000001010001111100100000011110110001001101001000001101101001101001001000101001110101011101110011111;
#1 $display("%b", po);
# 1  pi=207'b011010000001001111010011001001010100011100011000010110100101010010000101001111100110100111111101100011010110000001101010100110011111001100111001100010001101101011001000000100111001001010000101001100101000000;
#1 $display("%b", po);
# 1  pi=207'b001011101111001111000110110101100000111010101000101110101110110101011111001001110101110110100001011010100100111110100011000111100110000111110100011101101111110100110111110001000011100011000010011011110110011;
#1 $display("%b", po);
# 1  pi=207'b000010101011101110111111101101011101001110001101111110001000000010001001010100111111010101111111100110101100111101101100100110000111000000111100001101011111001101011001101001100100001110101101111010010111010;
#1 $display("%b", po);
# 1  pi=207'b011100111001110110100111001100110110111000110011111111111010001110100111101101000111101111000111001100110111100010100111010000001011011100111101001010011011101110111101101101011000000110011101001010101010101;
#1 $display("%b", po);
# 1  pi=207'b110010001001000000111111110001000100110000000011111100011000110110011101111111100001001111011100100010001101011110010010000001011111100011101010100110011010101110010100101111000110110001110110001101101100110;
#1 $display("%b", po);
# 1  pi=207'b001111000001110011011011001101001000010100101000100100110110011111110011011000001010001001100001110011111110101110111100000000011010100100000110000100011010000101001011000001010110110111001110110000011010011;
#1 $display("%b", po);
# 1  pi=207'b001000111100110101111011010000001011101111101011101011110101101001011100111111110100110001010111000110010011110110101001111000001101100011011001100010010101111100001101000000010101111001011000101000101100000;
#1 $display("%b", po);
# 1  pi=207'b011101000010101011011100000100011000100100001111101011101110011101100111101010110100110010000011100101100000000010100110101000001010010000110000110101011101100011010111011111101001001010010001101100100010110;
#1 $display("%b", po);
# 1  pi=207'b100111001101110010000101110100111101000010010110100101100110001000110011110111000001000110011000001100011100101111101010010111101101111100110101000111111100011101111000011111101000100101001001101111111000010;
#1 $display("%b", po);
# 1  pi=207'b010000001101111011001001000000011100010101101000001101001110001110101100010111100011000111000101011000111100011100011000011101001001111011011111001001110101110111100000000111011110110110111011110100000100110;
#1 $display("%b", po);
# 1  pi=207'b010100000100111011000001000101010010001011101111100011001010110010001001110110111110011100100000111010110100000010000010111100011111100101000011100000000111111001000001111000000001100101011010101111110111011;
#1 $display("%b", po);
# 1  pi=207'b000101101010101111010001110010010111111001010100111011011010100000101100010010111111011011001010000010000101101010001001101111100101110100111001001101001011010011001010110100101101010000001100111001110100000;
#1 $display("%b", po);
# 1  pi=207'b101010101000010011101011001010111110010100101101111100010111011010001001100001111010100111011001101001001011101001000101011110101110111010010110001101101001001010100110000101001011011001110111010111101001000;
#1 $display("%b", po);
# 1  pi=207'b100101011111101111111000011110100001011001010101001001010111001001001101100111000000010110100100000111001100010111101111001001111100101111100101100011101010111001111010101110101010100000000000101011111110110;
#1 $display("%b", po);
# 1  pi=207'b101110000011011000100100100011111001010010110111101011101001111100100011001111110111110000110010011111110111010010011001100000101100100111111100100011110000001111010000001000101110111111011001000110000100111;
#1 $display("%b", po);
# 1  pi=207'b110011111100010010011101100000110110001011111110001000010000010010010101000010011110100100101000100010010101110101111101010101110110100011011111100111001110001011111100110101001010011110110011010101001010100;
#1 $display("%b", po);
# 1  pi=207'b111001111011011011110110001011010000011000111100001100100001000001111111001011110101111011111010010111100011011000111110100001010000001111001001111110101111111100100011011010010111111110100100011111110100011;
#1 $display("%b", po);
# 1  pi=207'b010101011010101100101010100110000000110001000111001000010001110011110100110111011010100000110010011001000010111111111100110001000110100001111100011000111010101100001000010001011000101101100110110100100101110;
#1 $display("%b", po);
# 1  pi=207'b011011100110000011011111111101010011000011100001110100110000100001111001000111000010011001001110111101100110001100100111101010101011100010110101101010111010000100111011000001101000111110110000110110110100110;
#1 $display("%b", po);
# 1  pi=207'b011101110011001110011101001011011110000110110000100110011110100001110001101111011010101111111000010111000001001000111010011000100001011111001001100110011010001000110100011111010011110101000100101011111010000;
#1 $display("%b", po);
# 1  pi=207'b110111101010010110000111100111100001011011110111010111000100010010011110010000110110111110110101001100010100001101011111001010101111110010000001110010000101000110011011010000010010101101110000100110100100110;
#1 $display("%b", po);
# 1  pi=207'b000101011110101010000001010111000000000011000100001001111011110100111111110010000111000000010101011100001000101001011010001100100001100010111110011101111011111001111100011100110101111111011101011100011010001;
#1 $display("%b", po);
# 1  pi=207'b111010110111001110010000010100101010100001100010000110000001000110101010001111001011001000000011011100010100010010000100111001010101010110100011101000010011001110100110010000110111110000001100111000100010001;
#1 $display("%b", po);
# 1  pi=207'b010101101011100110000101011001110011010000010000111010100111100011000001001110010101111110101111011010111011001000101001100011000010000110110000010011001001011010001100101000101110101001100000111101110011000;
#1 $display("%b", po);
# 1  pi=207'b000010001111001000010001000101101101110100101000001001101101001001101101001001010101011000110010001110000100011111110011111110100100000100000000010110010110101101010100100000111001100011100000100010110100000;
#1 $display("%b", po);
# 1  pi=207'b101110001100001011100110000001100110110110111011001011001010000110001001001101011011110001000011110001101111000100011010010010011101011101000001011011001110100111011011100110101000000011111001100100000000100;
#1 $display("%b", po);
# 1  pi=207'b110001110000110110101111110011000111100101111001110001100010101110001101010110110110010110100010010001001000001011001001011000101011001101010010011100000001101101111111111110011100110000111010111110011011100;
#1 $display("%b", po);
# 1  pi=207'b001101000001001110100111011100010101110100010100110001001001011010111000010111111110100001010011000011000110011100100011011111001010101110001011011010100011001001101110111100011111000001001011010001100011011;
#1 $display("%b", po);
# 1  pi=207'b000000100100000010010011001101010101000110010000010011001101010100010000010110100000000111010111111101010000000001000011111001001111001111011000100100110011011010111010100011101001110000010011010110110110001;
#1 $display("%b", po);
# 1  pi=207'b100000010001011011110000011101101000110010001101000000000111111000111001001110011010001010010000001010100011110010110011110111000100111111111101011100111000111100110101110101011000000111111000110110000010100;
#1 $display("%b", po);
# 1  pi=207'b100001001001011100111000101000000111100010011100001000011011000111111001001000011100001100000000001110011101101000001100110100011111110010111001011111100101111110111110010100111111100011010011100101001111110;
#1 $display("%b", po);
# 1  pi=207'b110000111000110010110110000111000011010010100101101010000100110001001000111000010010010010100010001001011110000100000110110010101000000001010101100001110011110111000111000000000111101011000101101010010101010;
#1 $display("%b", po);
# 1  pi=207'b000000110011000001011101011101111010110000101001000110111111100100101100000100001011100011101011111110100011001110100011000100110100101101110011110011100000001010010011110001111001101111101111111011110101100;
#1 $display("%b", po);
# 1  pi=207'b111010011111101111101011010001111111101110111001010100001100110111011000101010010010011101001111101010111010010010000111011010000000101010100001101000100110011010111101110010011100101011011001000110100010110;
#1 $display("%b", po);
# 1  pi=207'b010010010001111011110111111010101010011011000000101010000010100100010000110101011111101101100110100011100001111110100111001110110110100111111100001110101101001010110101101100110110101100110110111110110011010;
#1 $display("%b", po);
# 1  pi=207'b111100100110000110001101000101101010000001110100010000110011100110110001010110100100011010100010001110000111011110111101001001010101110101001010111110010100000010011100101110011001110100000100100010011001001;
#1 $display("%b", po);
# 1  pi=207'b100011010001110101010001001101101101001000100100101101111111001101010011111001010001000101010010010110101001001100001100001111001001001010011010100001110011000101011111001000011111101111101100000000100111010;
#1 $display("%b", po);
# 1  pi=207'b101001010000001000011010110000000010010011111101001001110110011000010101011010000011110100100010111011100001011111111111100011000000001110011000100001101110001011010100000001101101110111001101011000010000100;
#1 $display("%b", po);
# 1  pi=207'b100101001111100110100111101101010001111110001101001010011010100110100010000100000101111110011010110000111101111111101000100011100000110011000000110110101000111001011010110111110011110110101111010101011100000;
#1 $display("%b", po);
# 1  pi=207'b110010010000010100010100000101100111011001111101100010001001000011100010010101010011111001111100000001110111100001001011101011100000011010101100011110001101001111010000010100010101100100100001101000100010011;
#1 $display("%b", po);
# 1  pi=207'b101100001010110001001000110010001111001010110101000110101001011000111000001110001100010010110100100100100110011111011100111000100010011100000100001011010100011001101101110010000001001100110100001001001110111;
#1 $display("%b", po);
# 1  pi=207'b101000101001011111010011100010010100100101001101000110101010111111001101011010010010101100001010111000111001100111010101011000111110010000100011110101111100111100010111100100010010111100000101100110110100011;
#1 $display("%b", po);
# 1  pi=207'b111100111100000110011001011010011010000101101000111010111110100100000011110101010111101011111100110001101100110100001001111100111100001001011101110011110111110010001010011101110101111100111101100100111001011;
#1 $display("%b", po);
# 1  pi=207'b010111111010111111001111011101111001110100101111110110001101011111011010010000000110001000100101100101011110000010001000100001000110000011111111100110000100111111100101100000010100001111011000110100000110100;
#1 $display("%b", po);
# 1  pi=207'b011101110010101111111000101010001111001111101011011101011110000001111111011101101011100000011100000011111100101011101110010001100000100111100111000010011001100101001000011101011111011101111111100000011010000;
#1 $display("%b", po);
# 1  pi=207'b000000110001011111101001000101111010010011110000011101011001111110100001100100001000000011000000000100100110100100110100111011101101110001101010010110100111001010110100010111010110100110100001100000110110000;
#1 $display("%b", po);
# 1  pi=207'b001001110100111110001011010110100000010111110111110110000000011011001010011000010100100010100101000110010101100010011010110100110101101001101100001011000111111000101101101011000010011111011000010000011111011;
#1 $display("%b", po);
# 1  pi=207'b011000101110110101110011010111011101011011000110111101011010100001100110101100011001110101100010011010110101000011010110010111111010110011011001101011011000100100111011011100001010110010010011000001010100000;
#1 $display("%b", po);
# 1  pi=207'b000110111101001100010111101011011000100111001110100001100001110010001111100100110010101111101010011011001011100000100100100000111010010000010010110011100100001010010100011011100011000000010101101001101010110;
#1 $display("%b", po);
# 1  pi=207'b001111010111110110001001100110111101100111010011100111101101101110001101111100111000111111000111011010010001011100111101000100100111010111000011111101011101000101010111111000000000111000111111000100111010001;
#1 $display("%b", po);
# 1  pi=207'b000011000000000101001010101011111010100111101001111110000001110000100000110000011101110110000101100010000101000110101001011011010111101000101000100110010101101110001010100010100000010001100111010100010010010;
#1 $display("%b", po);
# 1  pi=207'b100000111110001000100010011010000011100111110100100010011010111000100001010110101100101000110101111010001000110111010101100010011100100010000000011001110000010101101110111110111010101000101111000100111000101;
#1 $display("%b", po);
# 1  pi=207'b000101100001001001110100001001101000100111101000100110001100110110110100111101100100111110000100001111101110011110100101011010010101110101101011100100101000111010011000011001000010010110010001010010101111001;
#1 $display("%b", po);
# 1  pi=207'b101011011011010001010110001100101110101001010110011100000010110100010000101000011101001100011010001011000001111001101101110101100010100011000110010010001100011000011111000000100001110001111100101011000000001;
#1 $display("%b", po);
# 1  pi=207'b011101110000010010001101011010011000011100000111000000110111100101110111000000011100000100111010010010011110100110101110110100100010100101001100100111000010101001010101011000001001101110011011110010011001000;
#1 $display("%b", po);
# 1  pi=207'b100101010110100100000111011010110101111101101010101011100101111111000011110111011111011110110010011011011110011001111001000010111110111000101100100101110010100011111011000001010100110101010111000100110110100;
#1 $display("%b", po);
# 1  pi=207'b100010010011110001000011101111101001111010000101010100111010111001101100101010101111111000111010111101010101001000001010001110101000101100110010110011100101011011110110010010010100110100100101111111010000100;
#1 $display("%b", po);
# 1  pi=207'b010110111101101110100000111101011110010011001110011010011101010011011011000100101101000110001110000010111101111110011000010011110011010100111000111110111000100010110000001100101100101011111010011011000110001;
#1 $display("%b", po);
# 1  pi=207'b000011011011000010111001011010001000101110001011000011000101010000000101011001101010111101110100111010001000100111110001100110011100101010000011111100111011111000110110111001001001010101010011011110110001100;
#1 $display("%b", po);
# 1  pi=207'b010110111100101101000101101110001101101111011000100001001001111111010010001011100100101110101100010001001010000001100100001111111100110110101000101100100000010101011010100001101010000001100001100010111111001;
#1 $display("%b", po);
# 1  pi=207'b001011101100001011011000111111001000111100110111000100001000111111000000010000111111111110101111010110100110101011101011011110001010111010111100010010011001101001110000111010110100110110000101110000011001010;
#1 $display("%b", po);
# 1  pi=207'b111101110011110110100110010101100111101100110011010110010011011001101010010001010111011100011100111101111000110100001001000001100111011010111111010110011001110011010110100100010001111011011101010010100011111;
#1 $display("%b", po);
# 1  pi=207'b100110001000101010111011010100010000110100111111001111100110111100101010111101110100100000010111001111110100101010000100100101110111101011010000000101001110111011101111000101110100110000100111110000011111001;
#1 $display("%b", po);
# 1  pi=207'b000100111111000001001101010001100101000110010001111011000011011011001101110111000100101011110000000111001000011000000010010111010000101110100111111101101110011110000101101011101100110000011111111011101110000;
#1 $display("%b", po);
# 1  pi=207'b101111011101000000100100101100000010100101100011001111110001000000101100110011010010111011101100010110111110100101100011010011110110001111101111010101101010100101111111010000110010010111101110000010001101011;
#1 $display("%b", po);
# 1  pi=207'b000111000100111011010001001011000011110000111100010000111100000111011001010010110000001011110010010000011010000111100001111110101100001001101000111100001110000101110010101110111101101011110111000110001010101;
#1 $display("%b", po);
# 1  pi=207'b000110011010100111100011010010100010111110110100000100110111010110000100100101110111101001111100010100100100001000001110111010001010100011101011010101111011111100001101001110111111111011001001001110001101001;
#1 $display("%b", po);
# 1  pi=207'b101001000111100010000000000010110010101100100100111010000101010111011110010101110110111100101111100000100100100010011110010000100101111001100010011111000000011110111010111101001111111111001101000111100111111;
#1 $display("%b", po);
# 1  pi=207'b000000010110010110100011010110000010110000101111111001001100101100010011001110110100110000001010100100001000101111100000101001000111100101100011111010001001100101000101111101101101101011000010000110110100011;
#1 $display("%b", po);
# 1  pi=207'b000000100111001001111100110001111111110000100100111101111100110011100011110010000010001010001101110100111011100011100111110000110101101101101101110000001111110110011011000111111011110111001001001101000010111;
#1 $display("%b", po);
# 1  pi=207'b000000011100110100110000101011010000110100011010001110110001011101110011110010110101110101011110010100001110111000010101011000010000101110111011101001101111010000100111011100111111010100010001101100011000010;
#1 $display("%b", po);
# 1  pi=207'b011111011000010011110000110101011111001010010010111100110110000001100010110111100001100011010100001111010110100110011100000010001011011110110001010001001101101001111100101011101001101100000001010011111010000;
#1 $display("%b", po);
# 1  pi=207'b011011111110101000000001000010111110110010110111100110010111101010101110001001011011010010101001111110010010010110001110000100001111110101010101111111101100010011110110001100111110101111111101001101011000100;
#1 $display("%b", po);
# 1  pi=207'b010101100011111100111011101010000100101001111000010011111011010100100010110010000111110001000001101000101100011010111101001010111110001110011001110110011000011101100010100101011010101011111101111000001100010;
#1 $display("%b", po);
# 1  pi=207'b001001111010001111000110011001010001101010011101011101010111001111011001111100110100111010100010001101101011110100001001100101001110111100011111110100011100110011110011110101010001010000100000001100001000010;
#1 $display("%b", po);
# 1  pi=207'b001001111000000111100101000111110010011100001001101100100101001011111111010101101010011001111110011000101101011011111101000011100100101011001101110100001100010101011011111100100000110001010011010001100001100;
#1 $display("%b", po);
# 1  pi=207'b111001111111011010110111101110101000101100001001101000110010100111011001101010110111110011010010000101010101001101010111101101011100010001100111111000000011111111011001010010011100110001110100110100101010110;
#1 $display("%b", po);
# 1  pi=207'b000111011110000011000000111100100100010110110100011010101010101100010101010101100110111111101010110110101110111100100101101001011011011100010110100000011101110110001011101110010011100011111001111001000110001;
#1 $display("%b", po);
# 1  pi=207'b011001111010010000110010000110100011000111000011001100011100100001011001001001011110111111100111000110011101111001011011101001011101000011010011011100111001100001011111101001111011001100011101001101101111001;
#1 $display("%b", po);
# 1  pi=207'b111110111001010100011111001010010001000110110010111010011010001101001010010010101011000001111001000100100010110110110100110001100111100010010101011001001101100011011011100110100110011101110010001100110111010;
#1 $display("%b", po);
# 1  pi=207'b111000101111000101100010100100000011010101011111111111101110110010000010100100111011001111000100110001010011000110101000100011111101110001100101110111001101001110111100000100011110101111100001100000101101010;
#1 $display("%b", po);
# 1  pi=207'b111111111000101100000100000000000100011100011011001110111100010001101001111100101100100101010101101011111100101100010100000111010000100101001000000010110000010101010001000111110010000001111100011011101010000;
#1 $display("%b", po);
# 1  pi=207'b010101110111000001011000100000100111011100111010000010101101111110010111110000001110001011101001100000011010101001100100010000010000000001010010001100011011011110001000110110011110000100010011011111111111110;
#1 $display("%b", po);
# 1  pi=207'b010001011110010010100111101100001000100101100100101011010010100011100010110100010000101011000001100010001101110011001001100010010110001100011001100111101001110010010000001100110110001000110010110010111110001;
#1 $display("%b", po);
# 1  pi=207'b000100101101111011000010000101111100100000001100001110100110001001111110100010010101111000011101111111101110001111001111111101110010010100101101111010000111111010101001000010010010101010101111000100001110110;
#1 $display("%b", po);
# 1  pi=207'b100011010110001100100111100010101000101101101010100011001001101110001010111110101110001111010001100000010000111100010101000010101110100011100111111001000110111001101010010101001100110000001110111010100011011;
#1 $display("%b", po);
# 1  pi=207'b101110010101101101001011011011111110111011110110011010111001001001111111110110110001110010000111111010011001011100101110000011101001001101001001001101100101000101001100110100100100000000000011000111100110001;
#1 $display("%b", po);
# 1  pi=207'b111110101100001100111100101100000010000100101010000100011100010101111101110111010011101111101100111010111111111100011100001111000001011110110000000110110100010100011011110010110111010110110101000001110100010;
#1 $display("%b", po);
# 1  pi=207'b011001000110010101101000101110011110010001000000001111010110111001111010111011111110010010011101000110001111110100110110011100100111000010010011011110011110111010001100100010011000101001101001011111010111111;
#1 $display("%b", po);
# 1  pi=207'b111010001011001101011011011100111001000110110001101011100111000110100011110011011000000100100001100000100011001101110010011000111100100000011100011011100100011001110100011001101111101100011010101101111110100;
#1 $display("%b", po);
# 1  pi=207'b001011010000101001010001110001100011000110111111111001000110101101111001011001011101100001000110111000110011000110100001110110010111010111100101111011111010000101100001000111111111010111110011010000110011011;
#1 $display("%b", po);
# 1  pi=207'b001000000011101000011011010111011001100100101011110101000010100101100001101101001001100101000000000001000000000001000001110110101100000101110111001010000001111011010001000100110010101001001011111100110111111;
#1 $display("%b", po);
# 1  pi=207'b001100111101000110011101111110000100011101100111110011100001001111011010011001111111100100000100001111111000001101001000001011011100101110000100000110010101101011001111000111010110000110010011111100111100011;
#1 $display("%b", po);
# 1  pi=207'b011000011001111100111011111110100101111110110100000001110111111010110110100000000111111100111000011010010110110110010001010001000110010111010001011100010110010100111010100010101100001010010110000100101011010;
#1 $display("%b", po);
# 1  pi=207'b000101010010111001100010101011001111100110110111000100000000101101110100101000110010001111110101100101011101100100000100011110101100011100111000000010110100000111111110011001011101001111010111101100001100010;
#1 $display("%b", po);
# 1  pi=207'b100111100101100010110100001000000100001100000011000100000101111011100011110011101010010011010010101101100011011011010111100111001010010110101101111011101111011000101101000110010111110100111100001010011110001;
#1 $display("%b", po);
# 1  pi=207'b011011111100010001100010111011010101010100011001100001010011010001010000100011010110111110111000101000101010101111100011000111011010000101111110101110000010101001010111100001011101001110000000001001000010000;
#1 $display("%b", po);
# 1  pi=207'b100011010110111000110111010101110001101001000010110011100101111010110110101100000000100101011000011100110100000110001001101111010110000110110110000000001101110011011010001101101010110001001011010100000000011;
#1 $display("%b", po);
# 1  pi=207'b001010110100011000110111000001011101101101101001001110101001100010010110001100111101101001101100010110100101000101100011000010000111111000010000000011101001001111110000010110010100110001100100110000010011100;
#1 $display("%b", po);
# 1  pi=207'b001110110110101000101111000110100010000011011100101110011110100001001111001001010101101110011101100001000000000101001011101011100110001101011011010100100110001011111101001100010011000101001101111101000100111;
#1 $display("%b", po);
# 1  pi=207'b001101101100001110110101100011100001011010001010000001101111111110010001110010111010101111101000010110101110011111000011000111010111110101000011110110100001000011101000101110000011100110010000001100000010101;
#1 $display("%b", po);
# 1  pi=207'b100101111011011111011011101011111111111101011110101000000110000110110011110100011100001111010010010110110001010011001101000011101101001111011110101000000000000111111110001000001010100101100001001100110101000;
#1 $display("%b", po);
# 1  pi=207'b100010111110101100010101101111000110000100010000101000011011000111100101100011010000101011110101110111111001000111100100110111110010001101101001101000110001011011001011110111111110100100011001101001001100100;
#1 $display("%b", po);
# 1  pi=207'b001010001100001011000011000001001000100001110001011111000110011100100010110000011111101010011000110111101110010100011000110100101011011100101101000011010101111110000101000001000001010001110111100101100011101;
#1 $display("%b", po);
# 1  pi=207'b100010001100101101001100100010100001110001101011011111001100010000110111110000111010000101010011010000011001010001111000100000001111010101110011001000110011101100001010101011000110111110110111100011010101000;
#1 $display("%b", po);
# 1  pi=207'b010101101000011100100101001010000111000100101100000101111011001111000101001011110100001111101011111111011001111101111011001110000010101111001011110001000011011110100011100110101011001100001111100011011011001;
#1 $display("%b", po);
# 1  pi=207'b110101110001111111000100110000010100011100100011111010111111111101101000000011000100111001101100011000100101100110101001010100101100110000011001100000010110000100100001010001111111010100110111001011101011111;
#1 $display("%b", po);
# 1  pi=207'b011110100011000101110101010101000010010111011101110000001001101000111000110010101001011010100101110110011010000100000011001010001010000101011111011001001010110111000000111001010010010110111001011110101010100;
#1 $display("%b", po);
# 1  pi=207'b101001011101110101001110111001000011000011011111110001010100000111001111011001100101110110111101010100010000110000110010101110001110011100001111101110010101101001101100001111001011100011101000111010101001010;
#1 $display("%b", po);
# 1  pi=207'b000000111110100011001001101000110001011011001001111011000001000010000111011110101111101001101111011100110011011110110001000010101100110101011100000001111000001110110000101101000111100111101101100100110100010;
#1 $display("%b", po);
# 1  pi=207'b011011010111000101010010011111100111000100110000111001011000011101010011110000001101001010010001100010111000011101010001010101001100001011101011101000010110100001100011010010010110011101101001001001010111000;
#1 $display("%b", po);
# 1  pi=207'b101110100101000101111110111010111111101101110010010111010100010001110000101100100111101011000101110100001000010000010000000000010000101111110001011011000000101010001110111100000111101101100010011110001111110;
#1 $display("%b", po);
# 1  pi=207'b101110100000010010001100001000111000011001111110110111110111100011011001010000011100100100111101101000111101000111111010011100011011000110010110101011111100011111001000000011111100111110101000001001100101011;
#1 $display("%b", po);
# 1  pi=207'b000101011101100110001001111111010111010111111111101101011110010101110100111100111100101110000011010000110001111101101101000101101110101101000100101100001011100100100001011001001010100101101000011011000101011;
#1 $display("%b", po);
# 1  pi=207'b011111000010101110100000100111100111010100110101000011101101111011110011100110001011010001101010101110101001001000011010000000000110111011101101110110000111011110010111010110000010111100011110110010011000000;
#1 $display("%b", po);
# 1  pi=207'b001110111010001100001111100010001011110000111011111010000001001100001110100100000011101110010001111000100011011000101100101011011000100000110110000010000000001101111010000011100110100011101001000100010101100;
#1 $display("%b", po);
# 1  pi=207'b111101011000010111100100001011011010110111100111100110010111000010110110010111100011111001101101001110000110100110001111010000011001000011010100110110101101010110010101001010111110101100100101010010011010111;
#1 $display("%b", po);
# 1  pi=207'b110001110111111111100101110100010110100001110010101100100100101010100100011100010101010011110000111100001100110001010000111101111100010100010000011010010011111011001101011101001100010110111101110011000110111;
#1 $display("%b", po);
# 1  pi=207'b010000101001101010010011111011010110110011100010111101110000111001110010100111101101001110101111010011110011101100011100100110110101011101011100001011001111010111101101100101101111010011111001110000110100001;
#1 $display("%b", po);
# 1  pi=207'b010101000001011110000000100011011010010100111101101011011111010001101000000000100001111110010100001011001101011011110011001001110011100010000001111001111010100111101000011010000111111001001001111111101011100;
#1 $display("%b", po);
# 1  pi=207'b011111011011100000101110011000111110011010111101000001001110010011001010011111100000101101110110000000000111011101110001110111000011101010101100111110001101011101110111110001000010101010000011010000100000101;
#1 $display("%b", po);
# 1  pi=207'b011011101100101011000111101100010111110111101110110010110001001101010010011000100000111000110001111010010011010110111001100011101110011001011111100110011100110010100111011010010110110101001010010000010111010;
#1 $display("%b", po);
# 1  pi=207'b101110011110011101110011111001111101000010010100111100101101101010001010010100111100100000010010000110010100000010001100011001101111000101100100111001000000000001111110101011011100000000100001100110000000000;
#1 $display("%b", po);
# 1  pi=207'b111011000101010110100100011011101100000011001100100111110101100011001110111110000101001010001111010011110110101001011100111101101110110101100010010000011111010111111100001101100010001001001100101010000001100;
#1 $display("%b", po);
# 1  pi=207'b101000011001000101101101100011101101110000001110110111011010110000110000000011110000010011011010000111100101101000101000010001010010110110011011011100000101110111011000001001111000010000101111011001001010111;
#1 $display("%b", po);
# 1  pi=207'b011101101101111000010110011100001000100001111111100101111010110101010010110001110011010100010111100110110000010110000110001010100100101000111100110101101100111010111001100110110110010001110010000001001101111;
#1 $display("%b", po);
# 1  pi=207'b011110001011111110000111100011100011101000000011100100100010101000101110001011111000011011110001010001010110000111010101101010000110010111110000100110000000110100110101100111000110011011100010001001110110010;
#1 $display("%b", po);
# 1  pi=207'b110000101000111111010100100011111111011111001011110011011101100001011001011010101001010010010111111010111010011011001100101110011101111101011110100000111111111111011000011111100110100011110110000100001100001;
#1 $display("%b", po);
# 1  pi=207'b010100001011111001001100001001000101001101001011000001110000100000011111101100011010100000101101011101100000100010110100011100110100011001111110001011001111110011101010000110111101101011001110100100111100000;
#1 $display("%b", po);
# 1  pi=207'b010011100100000111000001001001110011011100000010011100100110111000011010111111011011001111110001000010001000110000011001111000000010111101010011110100100001100110010101001001110110011000001111001001111001011;
#1 $display("%b", po);
# 1  pi=207'b110000111101100011100000110000110111010111110001001001100011100001100100001011100010100110101001100000001101000100001000110100111010101111000111110011011010100011010111110110100010000000100110001101100110001;
#1 $display("%b", po);
# 1  pi=207'b001110001111111010111101001101001001101001101100110101011010111011000011000011010000111011101001010111001010001111011000011010001001100111100101001110101001000000010100001100001001010110000011110011101100110;
#1 $display("%b", po);
# 1  pi=207'b101011101100100101110000001100101100110010101100001100101011010010101001000101100001101011000001110101001001000001011001011100100100100110010000001111001100000001111100001001101111110000000111101000011010001;
#1 $display("%b", po);
# 1  pi=207'b000000111011010010100010001100001011101000000101101001011101011110110001001011110111100011010001111011001100100101111000001000001000110110010000110110010010000111001100111111000011000000000110001110011001101;
#1 $display("%b", po);
# 1  pi=207'b111101010010000110101110001001111010111000010101000000010100111111101101100011001001100110011001110110000101011001001110011000000000100101011000011000100101110111011000100111011001110110100101001011110110011;
#1 $display("%b", po);
# 1  pi=207'b101110000010100011111101011101100010111100000100101010101001001110011100011001100001011001111001010010010010101011101000011101010010100100110001111001111110011011110001101100110001001001000001100000001110100;
#1 $display("%b", po);
# 1  pi=207'b101100100100100100101010101101011111001101101111110000011001011011100000111110101110100011111011000001001100111110111011110011110110000101111111110000010011000100011000010111111011000110011011011000011010111;
#1 $display("%b", po);
# 1  pi=207'b111100110101110111001011000001001001011101000111100111011010101111111001011101001010101001101101011110011010101100100100010110101101111011100001111111001100100010110110010011110111000010110110110001001001111;
#1 $display("%b", po);
# 1  pi=207'b010011111001011011011111101101110111111011010011010001000011001011010111000011010111111010000001101110101110010000100100100110111011001101111111001101000101011101001000111001101000000111010100110000110100110;
#1 $display("%b", po);
# 1  pi=207'b110111001111010010011111110011101100001000101001000001111101101110101000001000111001100110011000100100001000000010110011110010101010100010001100111100000111010110110100001111110100100100010100101100100101011;
#1 $display("%b", po);
# 1  pi=207'b110101101001011100100100110011101011001110101001101110001111010010011110111010011010001101111000000010101001001100110101011101001101001001111001111110001101000011110010101111100000100111001000010000101001101;
#1 $display("%b", po);
# 1  pi=207'b110100011111001000111110011110111111100011110000000001111010111010101000010010000111110000001011000011110100011101101100100000101011100101110010011100100010111010101000001000101001001010011010101011001111001;
#1 $display("%b", po);
# 1  pi=207'b011101101011001011101101000011001000010001011001110100100000110010001110011010101001111100010000111111000111110010011010101111010110000101000101111011011100001010000011001101011001000110101111110111110011010;
#1 $display("%b", po);
# 1  pi=207'b010110111101000111011011011101010111011101011101101010010100000110000101111100011111011010110101010000001100110101101100010001000101101011101001110011001001111010001100110011110100111100001101111101101101110;
#1 $display("%b", po);
# 1  pi=207'b011110010000110010011000010000101110010100100010100000010111000111110100000011000110110110000101011100111000011001011010011000010000010101111100100011101000011010110001111100010011001101001111011010011001101;
#1 $display("%b", po);
# 1  pi=207'b110000110100111001010100111110111001100011000110100100111001001100010000011111111010011011000001010100010011111011010100100111100011100010000001101010100111111101110100000100100110010100011110011001110000001;
#1 $display("%b", po);
# 1  pi=207'b100101101111110111100111110000000011000100110110011100100110011101011011110111100101001111111010110011000000010001010100110010011100000111100101101000000101101001100100110100101011001000101111101011000010111;
#1 $display("%b", po);
# 1  pi=207'b000001111101111010001000111000000111110100011100111100000100011111011100000001001010100100001110111100100011110000011011000111011101111100100000001000011110100111000010111101101011100101100101001001011010010;
#1 $display("%b", po);
# 1  pi=207'b110111010101001100110111010011011000000100000101000011110111011011011001110111110011111110100110010011001101110001001100100011110101111010111110100100111101000101000000111011000011011110001111111011110101001;
#1 $display("%b", po);
# 1  pi=207'b000110001000101011010100110001100001101010111100001111011011001101011110000101010110101110000011101011010001110111110010000111111101000011101111100010011101000100100101101000011110001001101011100011100011011;
#1 $display("%b", po);
# 1  pi=207'b100011100001100101110110101111110010011111000100000101011001101010101001011011100110011010011000100000010111010000010001001000111100011101111110100110111101000010000011011100010100101000110011110000010000100;
#1 $display("%b", po);
# 1  pi=207'b101001000100111111110000010011011111011011000100011101100001000100111011110011100110111100101001111100111001011101110000010111110010111110111111011110111011100100110100101011110100011110101101000101001101111;
#1 $display("%b", po);
# 1  pi=207'b001110011000100001011111010100110110000011110000010100010110000100100001000011101110110111011010001110111001001100110100101011111010011001101010011101001000011001101111101010010111011101111100101010100100001;
#1 $display("%b", po);
# 1  pi=207'b001001000000100011001101010011111011001010100100010100011110000100011111000011011100001100000001100000100001010101011100110000100111110101001011110110011111111000011001101100101001101001111001001001001100010;
#1 $display("%b", po);
# 1  pi=207'b001100110101001111010011100111010001001010011011100010000000001110110010000111111010101000010001110100000111101110100011110110011000010010111010010100111010110000000110110111001110011010110011011001001110010;
#1 $display("%b", po);
# 1  pi=207'b001000100101000000101001110111001100110011001100011000101111000010010100110001000110110010101101001011001100111001100000000001010110110010101100101111100111101000000001101101111010100001100000100110001000000;
#1 $display("%b", po);
# 1  pi=207'b010001001101000001111011010010100001001111110010110100101010010100000110100100110110011111010011001000110111000010101110111100011010001011101100010101101000110010011100010011111001110001011100110100000010110;
#1 $display("%b", po);
# 1  pi=207'b011010000001010111001010111101110011000110010101110001000011000010010101111001100011001010010000101100100101100110100111111111001110100010110001010001001000100000001111101100001101011110100010000101001000110;
#1 $display("%b", po);
# 1  pi=207'b001110001000011010000010110010001000100010010001111101101011011010100100100100001110011000101101000000110010000000010000111111101010101011101111100101001000011111001110100101011110111011000001100011111100011;
#1 $display("%b", po);
# 1  pi=207'b010110000111111001000010001011101100101101001101011101001111001011100101000110001001101111110101101001101101111101111101110100101110011010011111010101100101000110000100100011000111000011101010100101000000001;
#1 $display("%b", po);
# 1  pi=207'b011000010100010110010111010010010011100011011100110000111011110001101110100111001001100000110111000111100010110001111000000000110000111001011100001101010000100110001111000001101101101010100010000010010000110;
#1 $display("%b", po);
# 1  pi=207'b011100001011100001010110100111110101000001110110010011000001000000011100100111011100000000011100001001111010011101111101010110101011100111011111000110110100001100001101111000010010111011010100001101111010011;
#1 $display("%b", po);
# 1  pi=207'b010100001101000100101000000011100000111101001010111100001110010101100100001010011101100101000100101100101100101101111010101011011101111100101111110000010100100010100110111010110101101110110001010110100000110;
#1 $display("%b", po);
# 1  pi=207'b000000100011101011101011011110110100100001000101001010110011100100000001101100000101001001100100111001000011001000110110110000101010111100010000011101010001101101110101001100000011010001100010001100011010110;
#1 $display("%b", po);
# 1  pi=207'b100011011000001011001101100010101010010100010101101100110010001110110111110111111001001001010001000000001100100100100010101100110101001100001001100010111110000001100101000110010011011101010111110000000111000;
#1 $display("%b", po);
# 1  pi=207'b000111111100010000011000111110111000111001010001101011010101100111010110001101100111010011110111010100011100001010111010110000011000011100101111010011000100000001110101001011010100011100101110000111000111110;
#1 $display("%b", po);
# 1  pi=207'b100100111000110010101001001101001100001101010000111011000000010110000011111101110111101001100110001011010010000110001100011101111110100001011010100111101110001001101100101000010010011000001110111100011111001;
#1 $display("%b", po);
# 1  pi=207'b000011000101001000110111110001110010101001101110111101100001011100110101100001110000001111011110111101111011101100111101100010101000110110100000001110110001001101111000011110010000101111001101011110000010111;
#1 $display("%b", po);
# 1  pi=207'b111001000000110001111111010001010111010000101011111001100000111111111000110001100011001010101011001110001110010000000101010110111111111100001011101100011101110101001100100101110010100011110000000100101101111;
#1 $display("%b", po);
# 1  pi=207'b100000100101110101111101101011010011100100101110100010000001111110000100111011110011011010001011000000110010000110110111101001110100000011100101110101101111011010011011100111010111001111011010111011101101011;
#1 $display("%b", po);
# 1  pi=207'b111101100001111010000111100000111100101011000110000011011111101101100010100011000100110001000010011100001011101000100001110011110001101101110110100101011101011000000001101000110010101111110110000101011111100;
#1 $display("%b", po);
# 1  pi=207'b110010001111111100000010000011101100011111010111111110110011101011110111110011001101100001111011101001001010011110101011000010111100111000001111010010001100000100111011111101011101100001101100001100110100011;
#1 $display("%b", po);
# 1  pi=207'b111000111010000110101011010010100100111111011100100110101011100001011010110001101000001011100111011101000110010000101111001100100001111111101010010110100000010100011101100001100101001000100110001011111100111;
#1 $display("%b", po);
# 1  pi=207'b111010100110101001010100110001000111001000010110111000110000010001100110000010110001011010001101001001100011001011000110010011010100000010101111011110110111111101100101010111101001110000111010001100111010001;
#1 $display("%b", po);
# 1  pi=207'b100110010001011111100100111010110010100010011010011111001110100001010011000011001011000010110011010111111101111000010100000001110110001110011111011110000000101000101001000001100011011001000110001011000000111;
#1 $display("%b", po);
# 1  pi=207'b010100001100011000010110010000100010010011001010010011000000011001101111011100111011110111001100000011110111010001000101110110011010110001110001000001111011001001010001011111111101110110110001001000110111011;
#1 $display("%b", po);
# 1  pi=207'b101111110100010111101100111010010110100100010010011001011000101001001010101011100010000101001111111001111111000001101011000111010010111011010000010010001000001011000010001101110001101011001001010111001000100;
#1 $display("%b", po);
# 1  pi=207'b101001001110011101110011000000100101100011101000101101011100100101110100110110010000110111110011011101100001111000100001001111010001000011000001001010010010101010111000010110001101010110001100011000101111111;
#1 $display("%b", po);
# 1  pi=207'b011011001011111101110100001011100010011001000010011001010010100101101001000100011111011011101011110011001100011010001000111101001010110001011001101011101010101111000011111111111110110111000110111110101111001;
#1 $display("%b", po);
# 1  pi=207'b111100110110101100100110101010011000100110001110110010011111100110110010101011111011011001011110011011101011001110100101111000011010011000101101001001101000101111101110010001100101000011001010001000111011001;
#1 $display("%b", po);
# 1  pi=207'b001101010001001111011100000010111100000010010110000111011101000111001011110000111000000111100111110111101010011000000000000100100111101100001000111000101111011110100111111001001100000011101000001010111011010;
#1 $display("%b", po);
# 1  pi=207'b101000010101110110111101110100110001111010010100111101111100111000011011100111111001110111100101100000001010101000110011101110011011100101111100110010011000000111110111011101000111011001011011000011000111011;
#1 $display("%b", po);
# 1  pi=207'b010111010001110101100111100011100100111110111001000111111110101111110001000001101000001011000101101010000101000000000111011010001111001100111100001100001000011101000000110001011001100000100110111010100001100;
#1 $display("%b", po);
# 1  pi=207'b001001110100100110110000010100001111101111001100000010100100101000101001101101001010111100101110001110101011011110111111000011100100100011011001111101111011001000000110110001001111110110010011110101010101000;
#1 $display("%b", po);
# 1  pi=207'b010010000101011111001111010001010111110110110010000101101100010110101100000100110011001111111100011101111100011001000101100000000010011010100001111000001000001000011111100100011101010001001011100000101101110;
#1 $display("%b", po);
# 1  pi=207'b111110101101000101010100110110111001001101110100111000101011100100101000111011011010010011000001110001100101001110100101000001001111101010001101110000111000011010100111100001001101011001100011101100010011111;
#1 $display("%b", po);
# 1  pi=207'b110010010100001110001100100010001110000010111101010011000100101100001101100001100101010010110011011111100100110010100110111110010010100110011100010001001010001001011101111001011000011001101001011000011010001;
#1 $display("%b", po);
# 1  pi=207'b010100100101101111101111000110101110000010110101110011011011011101110111101100011111111000100101111010101011101100011011110011101100110011100110000101111010010101100110010001011010111100101010100110000110110;
#1 $display("%b", po);
# 1  pi=207'b100010001010101110001110100010111110011100001100110110011110010111100101111011000001011100000101100011011011000111101001010001110001001101110010110110101101000001010001000111101000111010110100010000010100011;
#1 $display("%b", po);
# 1  pi=207'b110110001101011100101101000111111001110011011101001010100100010101010111111111111011001001001101011011110010110001100011000101011001010011100101111101001010001101100110110101111000101000101111010100100110000;
#1 $display("%b", po);
# 1  pi=207'b110100101010000110101001010010010101101111000011101010000011101001100111110000101110110010101010111101101010110110100111001100011010110101011101000001011110100001101010010101011000010110111011100010100011101;
#1 $display("%b", po);
# 1  pi=207'b101100111011011100111111110000010110101111110001110101001011001001010011001100111111110000101101000000000010111101011101101101110001011111011000001000000111100101110010100000101111110010101010000100011011000;
#1 $display("%b", po);
# 1  pi=207'b001011001010001000001001101101100000110101100100110010010000010001010110111100100110011000011110011010000001011010011101011010010010100101010010011101100001010101010110110001000111100101000100101110100000011;
#1 $display("%b", po);
# 1  pi=207'b111011111110001111100101100001000101001001000011111100111111011000101010101001111011001000110001010001110001000000101101110100110001100010001110101101110001010101011011000000001001010100001010111110001110011;
#1 $display("%b", po);
# 1  pi=207'b001011000000110010000110101111111000010011101100100001101111100110111000010111011000100011111111111100010010010100010011111110111100011010100110100101101000000110001110101001111001100011000001110001101011010;
#1 $display("%b", po);
# 1  pi=207'b000001100110101000110101100101000001110010111010100110011011110001100001101101000111111100111110001100000010011101101001011110000001101011100001101101110111001111101110100000111100111101010100101000011101101;
#1 $display("%b", po);
# 1  pi=207'b001010111100110010100000111011100011011101000101010000011001100101100100001000000100001011010011100001001110111111001010100001110001010001101000010111101001001110000100111000001010011101000000100011010001000;
#1 $display("%b", po);
# 1  pi=207'b110111011010100111110101110011011010100010100111111100000001011001111110010011101010010101110100000000101001101101100010011011101010111011100011011100011011111111010010101011010101111100010101100001011010100;
#1 $display("%b", po);
# 1  pi=207'b001010110101010000100001000000100111011010010100001010001010001010000000111110010100001101001001110100110001101110010010100011010111110010110101011011100110010010000001000111101111011101100110101100100010010;
#1 $display("%b", po);
# 1  pi=207'b011110000111111110111110000101001110001001111101010010110110000101011100110100111110111101111111001000101101110111100100101000011001100011000000100011100010011011010111010001011111011011110101001011101010000;
#1 $display("%b", po);
# 1  pi=207'b000000001011110001000100011101010101111100011001110101100100001100101110001000000100000010111011011110101100110011010011101000001111100111010111001011011001011000101000010101101110110110001010101101101111101;
#1 $display("%b", po);
# 1  pi=207'b110001011001001010111000000110010000001011110000101011001010000111001110000000110110101000010011000001100001110100100011101110100000001000000010001000001100100001000110010110111101111101011010101010011011000;
#1 $display("%b", po);
# 1  pi=207'b011001000110000111011000000111100100011110111101010111010010010110000011100110001101000000001011100010110101100100001011100100001100010010100101011001101100110010010110000110001011110100101101100110011010100;
#1 $display("%b", po);
# 1  pi=207'b000100101101111000110000010100010011001101000000000011001111100110111110111101111100100110110011011100000000011001001010111010101000111010011101011100100100100111011100100010011101111000111000001110011010111;
#1 $display("%b", po);
# 1  pi=207'b011100001001111110101010001001011111100000001000111101011101001101000100001100101100000001001101010000111111010111000110101100010011100001111000011101100000011111001100001000000111010111111010010010101000111;
#1 $display("%b", po);
# 1  pi=207'b000001011110010010010100000111011111000110110000011010001010111010001010101100100111000011010011001111000000110010001011100000001010000111000110100010000101001011111111101100001101111010101001010010001011001;
#1 $display("%b", po);
# 1  pi=207'b100011101001011011111110011010101000101011110000100101111000011010010110101011100000000101100101100010001000110011100101110000101011010111110101000010010000000110100100000001110111000010000111110001001011010;
#1 $display("%b", po);
# 1  pi=207'b111111010000100010001010100001110010000000110100010001100000111100010011110100110011100100110110000010111010111011000011101110011110110010110000010100001011011110101100101101000100011000111110001100010101011;
#1 $display("%b", po);
# 1  pi=207'b111011000001011110101010000110001001010000010000111001101011000100110111110011100111110100101010100011100010100110110111000101011001011110001001000010011101000011110011111111011110111100110101000001111001010;
#1 $display("%b", po);
# 1  pi=207'b011001101010100111011010110110101010000011010010000011010101100110100000101001100000110011100001110100101100110111110000000001000101010110110101010001111100100000111100100000110001000110110101011010100011011;
#1 $display("%b", po);
# 1  pi=207'b000011111100000001001111001001101001111000111111000100101010100010100111001010000000011011100110010000010110111000001111110001111110011101111001011001001101001101001011101110110010110000001110110000011100100;
#1 $display("%b", po);
# 1  pi=207'b101011100100111100100100010000010101010001110001010001011011000011000100110000011001110000010001000001101010101001100101100111101100001000101100001101110011101000101110101000100110001010011000011010110110100;
#1 $display("%b", po);
# 1  pi=207'b110010100100010101001011111011101111010100101000011101101100011111110000101000011011000100101111010011010101001011001110000100100101101111000111111000111111100111110000011101110110011111000111010000101111001;
#1 $display("%b", po);
# 1  pi=207'b011111000010011010010110110101101011000011011110010110000110101100000010101101110100100001110111100001000100111101010000000011100011100101110110101110101011011010100001100111010111111111101100100111011000000;
#1 $display("%b", po);
# 1  pi=207'b001101010010110111110010001011100000001000100110010110000110011010101010110101011000001010000000101110000100100111100100011101010001101000111001000000111111000101111111100111111000010011110000000110111010000;
#1 $display("%b", po);
# 1  pi=207'b100011101111010101101011011110010000001101010011111000001000010011001000100100001001110111100011100000001011010010110001001111101000010110100100000101100110011101110111000010000111110110111100010000011100100;
#1 $display("%b", po);
# 1  pi=207'b010001001010111100010000111100000010101101101011111110100101001011110110001111110101010100100101111010001011101111100000000000100100100010001100110111100011110100110111111101110101000011010010010101001101010;
#1 $display("%b", po);
# 1  pi=207'b000100011010010101100010000001100111111100011011000011110111111011001111100110111000000111111010100000110001111110111001111101111101100000011110111000010111011011010011111010011011110111110001001111100111111;
#1 $display("%b", po);
# 1  pi=207'b100000101111111110100100100101011001011001101001111111111110110111001011010101111000110001011001111101101000101101010101110000001010111011011101011011111110001001011001111001001001110111010000010010001001001;
#1 $display("%b", po);
# 1  pi=207'b100110010001010010110110101101011001101110100101000101010010101011101110111001010001001110110100110000000101010001011100101100101000011010100111110111110001000100011010101100101111001000001010011011010110100;
#1 $display("%b", po);
# 1  pi=207'b101011010001100000111001010001100010001111111000101110100000101011001101101100000001000110101010101101000100010011100011100001110001000101011000111111000010000111101101001000000001100000111000100101111100001;
#1 $display("%b", po);
# 1  pi=207'b111010101110110100100100011110100000011111001111110011100110101011110111101111101001101110010100001101000110110000010001011011010011111010010010100000111100001100011000100100001000100001110001111101001111000;
#1 $display("%b", po);
# 1  pi=207'b110110101101111001011010110001110110001100011100010100001001010010011010001100110111011010001101010011110110111011001001111110000111111000000111000010001001000100100011100000010010011111001001010010101111100;
#1 $display("%b", po);
# 1  pi=207'b110110111011110110001110110110111100010100100001001101000100101001000111111010100101100001000001010101111011101000110010001100010100111100111100010000110001101110111010001110001010100111010101001101011010100;
#1 $display("%b", po);
# 1  pi=207'b111000010111010000110111001010000001001110101111111000101110110111100001000111110101001111010011010100110110010001010000110001111001110011011100001010010011010100100110111101101011111100001110111010010111110;
#1 $display("%b", po);
# 1  pi=207'b100000100111001101010101001101011101101000111101010100010001011100101010010100011101011110001011100001010011111101101110000011100010100000010111111011111001001101010010011001000111111000011110010111010001101;
#1 $display("%b", po);
# 1  pi=207'b010010000110110111101100001001010011111100000101110100111101111110000101000101001010010010000110011011001011000101110001111011100111101001010100110001110100101101110000100011001000101101011001011101110110011;
#1 $display("%b", po);
# 1  pi=207'b000100101000111011000000000000101000011011000001100010000100100110010010000101010101000000010010001111010111100000001011011001111110000011000000100100001011111101011001001110110011000010101100010100100001111;
#1 $display("%b", po);
# 1  pi=207'b110001101001101111011011001010000111111101000010000011000001100111110111101100000111001001100011000100110001001010111010111010011011010001001010011111100100110101001011000111110010111110000000100010011000101;
#1 $display("%b", po);
# 1  pi=207'b110001101011011001001110101000100100100000011010100011001111110110000100001110111101101010111100001110110000111010110100100101010010001101000001100001100001000010000110100111110000111010111010011010000001101;
#1 $display("%b", po);
# 1  pi=207'b011101101010111001001011010100010110110101101011011110010100011111010010111000110110011011110010101110011111000100100011010101000101000010010111100010000011000011110111011011001110000111001101100101001110101;
#1 $display("%b", po);
# 1  pi=207'b001000011100011011111010010000110001010111100011001100000111011001110001100110001000110011000000111010101111100111101011011100000101011100100010100101000000101111111000011110101100010000011010111101100110110;
#1 $display("%b", po);
# 1  pi=207'b000110000111001110110000100100010110001000010000010010110010101110110110001111111111000011111101010100101001010110010110011101010011110101101101010010001000101111000110010011011000110101010000110110010011000;
#1 $display("%b", po);
# 1  pi=207'b101110100110101110100001110010110011101100011110100001110101100101110001010100100010010001000111111010101101001111000000100010101010001001011011011110100001010011110111101110110100000001000001011100110010101;
#1 $display("%b", po);
# 1  pi=207'b111001011111011111110010100011010001101011001001011001101101000110001000010101110101111100101000000010011110001010111101111001101010101000000010000011110000010100101001010000101011010111101010101100100110000;
#1 $display("%b", po);
# 1  pi=207'b111110000000010011111110111100001101100011101101010110001010010101010000000001110111110010110100111000011111001011011010101001100010100110101110100010111111101010111110100011000010110000111110100100001011100;
#1 $display("%b", po);
# 1  pi=207'b000111101101110101111100101101011000001001111010001010011110110010001100011010111001101000011110000110101010001011100000000000110001110010000011000110001101111001100010001010111110110101000100001000110010110;
#1 $display("%b", po);
# 1  pi=207'b100000011001111110111101001111110110100110011110111110110000000000101000001010011110111100110100110011101101001100110010010001001001100111010011000110111110101101100010101110101100011011110110001111101010010;
#1 $display("%b", po);
# 1  pi=207'b011110000110101010101011000001001000110001100101010011100101111111000000011110111111110111011010000010011100001000001001110110010101100111001011111011010000000101010011001100001001001100101111011101011100001;
#1 $display("%b", po);
# 1  pi=207'b011000110111000110101001101010100110001100101111110011001001111010101110000111000000010011111101000000101100111110111001001000001000101011111111001100000011111100100000111011110100010001000001100111111010010;
#1 $display("%b", po);
# 1  pi=207'b100111100010111011010001111111111100011000010111110110000100010110101001111100010110110100100101011011110011000010001000001100101101000101100000011110100100101101001101100101110110111110101010101010000110001;
#1 $display("%b", po);
# 1  pi=207'b011010011111001100100001111000000110110000100010001010011111000111100111100110111100001101101100010111011100011111100010111111101011010100101001001001100110001111101110111111011111011101100111000001010000011;
#1 $display("%b", po);
# 1  pi=207'b101000001000011000010101011111000001111101111001110100000000011011010100001101110000010001100011010100100100001111010011001100100110010110010001101111101100010011100011010100110111110011000010101110010011011;
#1 $display("%b", po);
# 1  pi=207'b001010100110110101100011001010110110101001100111010010001000010100010110111001110000100101010000110001100001001000101110101010010010100111001101100000001010001000100001111011101000001000100100001000000000100;
#1 $display("%b", po);
# 1  pi=207'b011011110110111100001010100111100110101001110011000011101010111000101101011000010000100001110000001011101011111001000011100100100000000001011001101100010011100010010111001010000011111100101110001000001100111;
#1 $display("%b", po);
# 1  pi=207'b011100000110001110110101001101111101101011111001010011111010010010001011010010111010101011000010110000100010101101111110100110110011010100001011010011010000000110011101111001110110010111001111111010000110000;
#1 $display("%b", po);
# 1  pi=207'b001100000010000111000001011111111001000000111100100000011111000110111100010001100100011010100001101011100110001101101000000001001010001011110011010110100100101010101001100000001001011111101111111000001000001;
#1 $display("%b", po);
# 1  pi=207'b000011101110111001001110110110100101110010111011101010010000011010110101010011001100011100000111000011000101110110011010011001101100111011111100001101110010011110011111110111110001101111111101001001101111011;
#1 $display("%b", po);
# 1  pi=207'b110101110110000101111111000110010100100011000101001100011000000110110101111100000100100010101001100011101110100110000101101010111111110111011011101001001010011001111010111011111011110100110101000100111101100;
#1 $display("%b", po);
# 1  pi=207'b001100110000001011110101110000100011100111100110100001011110111010100010010100101011100001011111110000111010111110011011111110111010010101110000111110001111100001110001110100011100001110010111101000011110001;
#1 $display("%b", po);
# 1  pi=207'b100100010010100110111011100111110011010110100011001001011011100110111011110001110001010110111000100010010100010001010010010011011100110100100000000110111110010000000110011101110101100011011111111111010001010;
#1 $display("%b", po);
# 1  pi=207'b100110110010100110010011111110011001000100010100001001111011100110000111101011010101100111011011100111010000110111110111111011011110010110111101000110100110110101100111001110011001101110010100100110110110100;
#1 $display("%b", po);
# 1  pi=207'b010010101010111100010000111010011101101000110011101001011110001100111100001010000000000011100100110000011011111101000110111011010001100110000001000111010001111100100111110111101101110001010101000001001101011;
#1 $display("%b", po);
# 1  pi=207'b101100000111110100011001000111100001000111110111101011010110110001100100011100000101010100101001000010111011100101000100110110111111011010110110100011100011000111000011011000001010101000011010010100110111111;
#1 $display("%b", po);
# 1  pi=207'b011101110101111000001110000101010011011000111100010010100100001010010110110011000101010100001100000100101000110010111011111001110011001011000100100001110101111100101011011111000110111101001100000011110000000;
#1 $display("%b", po);
# 1  pi=207'b100001111000001101101001010110001110111101111101101111100101010111001011111000100010011010010100101100010001001000100110110010101010100000000011001101110111100000101010001110001100101010001110111100010000000;
#1 $display("%b", po);
# 1  pi=207'b010010110000100100010111011111000110111101110100100010010001000001100001011000101010000010010001100000100111110110110110011001010010000001000001111001011011101011110001101110001101100000000001000100011011001;
#1 $display("%b", po);
# 1  pi=207'b101000100100110001100000101101100010110101000100000010000101011011110010000100000010101110110000110001010110011001011110100011001110000111011001010110101100101110011110010101110010000110001000011001010011110;
#1 $display("%b", po);
# 1  pi=207'b100011100001111110001110000101110000000001011011101111000010100011110100011101000001000111011100001000110010011011110000100000100110110010000111110010110011111100001000100001000011011010011010100111011010100;
#1 $display("%b", po);
# 1  pi=207'b100010100111011011111100011001101000110011101001001010101100111000100011110101011010000111001010010111000001000000100001111111100100101110011111000010111101011100111011101110110001111000101010101010011111011;
#1 $display("%b", po);
# 1  pi=207'b101011100010001011110100001010011011100101011011100010001001000000101001011100101100111100100110111011001100101010000100000011011000011010100110111100010100000010000111110000100100000111111110110001001000100;
#1 $display("%b", po);
# 1  pi=207'b111000000110111010100110010100010111110110001100101011001110011001101101001011000110100011011101001111011010110011100000010100011100111010000110100101100000101111110110110011110100010010001100000000100001001;
#1 $display("%b", po);
# 1  pi=207'b110111011011011010100010000011111101011011111001110110011001111010101010011011100000111111000110010100101110101001011100111110001100111000001111010001011110001101001100110101110100001001101111001110110010010;
#1 $display("%b", po);
# 1  pi=207'b101000100110011001011000100110111000111100001000011111110110000110101010001011111010110100001111000111101001001101110101001111001110111101011011101100111101010110000110000100011100000011000111011001011110000;
#1 $display("%b", po);
# 1  pi=207'b001011111101000000110110100111010100100100000100000100110100110010001010001100110101011011000010011100000000100001101100010101010110011111110000000010110100110010011111111101011111010000101101000101011000100;
#1 $display("%b", po);
# 1  pi=207'b000100101010111001001010000101001101011111001101101000011110111100011010110110100110010111101001000101101100010001100011001101111110110100011011011010110101010011001101100010011001111011100111001101011101011;
#1 $display("%b", po);
# 1  pi=207'b100110010100010110101110000100011110111110101101110011111100001010101000101010110000001010011111100001010010111100011101111110101000000001000011000000100011100001001010101011010010100001101010001101111101001;
#1 $display("%b", po);
# 1  pi=207'b100111010000100000010000000010101100010101111010000011111010111000001111101111010100011111100111110100101010011111101111100000100011001011010100011010001010001010001101000111000011110111101001101001010111111;
#1 $display("%b", po);
# 1  pi=207'b001100110111111010100101110111100110101000011111010010111101111001110001111001010001100011000000011101001100110010100000100111110010010100010101001010011111000000101101010111001110011000110000010001010011011;
#1 $display("%b", po);
# 1  pi=207'b011001100101000011001101110001110011111001001001001000100111011000011100010100001010000010101111010101101100010111001011000011001101000011000110001010110101010010011011111000101110000100101111100111111101100;
#1 $display("%b", po);
# 1  pi=207'b100010000101001001010111010100110110110010101101110011011111100100001010111001001011001010110001101001010001100001001110111000110010100101011110000010001101010011000001010011010001100011000001010000101010101;
#1 $display("%b", po);
# 1  pi=207'b110001000111001011001100001010001101111101111101011010100110111001111000111100011101000101100011000000001001001101000010011111111111100100001010010011010000000000111001010010000101110101000001011101001010100;
#1 $display("%b", po);
# 1  pi=207'b100010101010100100010110000110001010111101011101010011100011110100001000111010100101011100111101011000100100101010101011001001000000000111110001100100101100101100001010100010110100011011111101101000010110110;
#1 $display("%b", po);
# 1  pi=207'b010001010111011100100001100101101100000010100010110011111000001100100011011111110000011111100101100010000110000011110000111110110010101000110010100100110011001011010111111110111110010101101010101100100010001;
#1 $display("%b", po);
# 1  pi=207'b100111010010010101110010100011000001011011100100001101010110110101101111101000111110111011001001001100100000001111011110010000000100011110011011001011000000001100110111001011110110100100010011010010001101001;
#1 $display("%b", po);
# 1  pi=207'b101110001101001001010010010111101001111011001100010110001111110110000110101100111110001110000101100110100000101011111110011011010010101110001000100100001000011010111001101011000000001010010101110010100101001;
#1 $display("%b", po);
# 1  pi=207'b110010001101010101101110010110010111100010010111111111010101010011111101010101001010111110010000000111011101101111100111010001101000011100000010000100111100011011001100110111101111010101010100110110000111011;
#1 $display("%b", po);
# 1  pi=207'b101010001011010010100100101010000111010100001100001010110110010001100011110001110100001110100011111011010110011001100000101111011000000101000011100010001111010110001001011000000100011010110100011010001001101;
#1 $display("%b", po);
# 1  pi=207'b000111100011111101001000111100101110111100111111100100010010111101111110101110111110010100000101001011001010011001101100000000101100101000110100001111000100101100110101100110010100011111010111000100001101010;
#1 $display("%b", po);
# 1  pi=207'b111110111100111011101111100001110111010000110101001011100011000000000000111111011001000000100110011000011010110100110101111110010101011101001100001110001011100001010011100101111100000000100100000001000001010;
#1 $display("%b", po);
# 1  pi=207'b000110101010100010111111111010011110100111001010110010101001010101111000110111111101110011010001011111001101101100101100010011101011010101010100111000001100101000011111110111110010100011100000110000011001100;
#1 $display("%b", po);
# 1  pi=207'b100110011010110011100000111001011110110100000001001110110110010001011010100001001110011100011001001001000000011000011100010001110101010100110101100001100111100010001011101111000101011100110001000000101001011;
#1 $display("%b", po);
# 1  pi=207'b010011101000011000101100110000101001010000010011001000000111100100010100101011010010100111000010100101011101111000011110000001011010001101100010111011110100101010101001100000011010000000001011100110011111101;
#1 $display("%b", po);
# 1  pi=207'b000110101001101010111101001110000110101110110001101010000001011110000000110111110011000000111010001010001001001100111111110000011000011011010000000110001000001000101110010101111001010010111100100111111110000;
#1 $display("%b", po);
# 1  pi=207'b000001111110100000001011110000100000000100010100000000111111001111100100110111011110101110100101100101010000011111001000000000000111100010000001000010110101101011100111010000000100101110100011101110000001000;
#1 $display("%b", po);
# 1  pi=207'b000100100100001101100110011101101001000010000110111011011010010011101111011010100001111011000011101010110010000101011010010011111110101011001010100011100111001101000110100011000001100000011100110010110110101;
#1 $display("%b", po);
# 1  pi=207'b011110010000011010001111010010000010101010000100001100011111111001111100101101000011100101010111110001011001001011010111011001111010010000111101000010000111101111010010101110101010010011011100111001100100101;
#1 $display("%b", po);
# 1  pi=207'b110000110100011100101101000010000110110111000111110111111000000101011000011000011111011010011110101100100000011110111101110111001111011010001100001011001111000110111101010001110000000010111011000100010001001;
#1 $display("%b", po);
# 1  pi=207'b001101000101101110101101110001111011100000110011011110011111100101010110011010110011000010011001001001100010011101100011110110101110010000011111100110011111001111000101010110011011001111010001101111110111111;
#1 $display("%b", po);
# 1  pi=207'b100100111110001001001010110010000001101111101011011010001111111001000101001111001111000001111010001101111111111100100010101011010100010100100101010010010111010111111101001110110000001001110000010000101101101;
#1 $display("%b", po);
# 1  pi=207'b010010010110110101001110000000001110001111011010011110101000001001000100111111111110001011011010010111010101111001100010011100111101101111100000001010101101110100100001001001100100111001100111010000000010001;
#1 $display("%b", po);
# 1  pi=207'b110101001110010000110000001101001011000000101100011101101101111100001010011001010110011101111111101000110011001111000010010111110001111001100010101110100110111011101100010101110011101010011101001010110100100;
#1 $display("%b", po);
# 1  pi=207'b001011110010010011101110100111011111001001001111110111100010101111011001011011011100100110010010001011011000111000111110010011110000011010111001010110011101101011010001000011001010100111101100110000010001110;
#1 $display("%b", po);
# 1  pi=207'b110000110000101110101000111100110001001001101110000010001101110000011011111000001100001000101010011001111101100100001110011101011001011010110101110110101010100000010111111011100000101111100010011100001101111;
#1 $display("%b", po);
# 1  pi=207'b000110000000111001000110110110110011000011101001011111110011101010101011110100101111011110101110000001000001011000011111100001100100110000111100100000011111101101100011101011111010101101011101001011001011101;
#1 $display("%b", po);
# 1  pi=207'b101000100101111000011001110000001010101101110110100110101100101000101100110110011111110101010100011001000111001001011100011110001000111111111001101100001110111110000000110100100110101111001010001011101011010;
#1 $display("%b", po);
# 1  pi=207'b010100011001001001000010101111000111100000011100000000000101110001010010001000111110000101111001001101011101100101100101100110111111011100011111111101011101111000011001001010010101001010011101010101010100101;
#1 $display("%b", po);
# 1  pi=207'b011100001000100100010100010100101010111100010001110100110100010111111011001011001011111010100110111010000010110011000100110100100100110000101110010111100010010010100010011010001001001101010110110010010010000;
#1 $display("%b", po);
# 1  pi=207'b001000010011000110001011111111010101100101110010111011001111000011001111100111000011100101000010010011000000101011100111100000010101101100010011110011010011000111110000010111000111000100110011101001001011110;
#1 $display("%b", po);
# 1  pi=207'b001010001100101000110101010101011011111001100100101000100010111110010101101010000000000110111111000111000011011110000100001011011101111111010110110011100110010111110001001100101000110101001100000010110101001;
#1 $display("%b", po);
# 1  pi=207'b101000100001001110100111111001010011110110110000001111011111101001101101010001011000000011010011001011100011111011101010111010010101100100110001010011001111010000000110011111011010001100001111100110011010111;
#1 $display("%b", po);
# 1  pi=207'b111000010100000100001111010101100110100100000011010100111011100011111000100110110011010101001000000100000000010001010011110011001001100010110101001011011000000010000100110000010110111110100011111111011101010;
#1 $display("%b", po);
# 1  pi=207'b001010011010010110110001001010101010000101011110011010111110111110110100011001010100010001010001010011000111111111111000001100100011101101100010010100000100000100111010101000010100101110110111001010100000110;
#1 $display("%b", po);
# 1  pi=207'b110001011010101010111001110000100111111010010110111000000001001011000000100011110011100111000011110000000111101000011001001111100011010000111100000001111011111000101010000011011111100011001110000111000100000;
#1 $display("%b", po);
# 1  pi=207'b110110011111110100011010011101111100111100111000101111100000100101100101101011111101011001101000101010111111101011001111110011101110001110000010100000110110010101110110000011011000100101010001000011011110010;
#1 $display("%b", po);
# 1  pi=207'b110101010000010000101011101011100110011000011001001100001011010001100000101101011101001111101110001110100100000001011111001100101100101011100001101100000010011011110011101010111110001010100100001001110101010;
#1 $display("%b", po);
# 1  pi=207'b001001010101111000011000000111100000001111100010100110111000111111011101000010100110001001101101001001000111110110001110100110000101111101000010001111010111010110010001001110101100101100111101011000101111010;
#1 $display("%b", po);
# 1  pi=207'b011011010100000011011100111011000111111010100110000010100011101110000100110000000010110010101110001011110111000011011011111010011011110010011000001110110011110111011100011011001001100001011110011101111111101;
#1 $display("%b", po);
# 1  pi=207'b110100010000110110100010010111000110011011110101100011111100111000101110100101100111010010001110011100111111101101011000010100111001011101101111010001000001110110101010100000111100110100111011010001111110111;
#1 $display("%b", po);
# 1  pi=207'b100110011010000111101010100100110000111101101111111000010111111101110110011110110010101110010001011010101010101110011101101110011110111011101111110100110001001111110111101101010111110111111100010111010001010;
#1 $display("%b", po);
# 1  pi=207'b011001001101010011100101011101000101111100101010011000001100100111100100011101001100000001101011010100101011010100011110000001010000000100100110001100001011101111111011010000000110011100000100101001001011111;
#1 $display("%b", po);
# 1  pi=207'b001001001101100111110110111010000110011000001110111010111000001000111010101010100000100000111101111010100001110100001000001001010001001000100010011110000100101011111101101000101010111110000101111001111001011;
#1 $display("%b", po);
# 1  pi=207'b111110111011010111100010010111111100000101100111001000100101101110001110101011110110100011100001101110011001111100010010100101001101101100111101101000011001000111101010101001101000011100001101010101110000101;
#1 $display("%b", po);
# 1  pi=207'b101011111010001111101100111111101101000110111011111111001010100011110000000110111100000000101010111100110111101010101101111000010011010011010100010100110001110111001111011111100001101011011001011000001100000;
#1 $display("%b", po);
# 1  pi=207'b011101101101011111100011000101110001010110000101100010111100110010111101110010001101010110011011011110010101100110111010100011110101111110000101100110000010111110100011101110110000110100110000100000100101010;
#1 $display("%b", po);
# 1  pi=207'b100100101000110110110001011011001101101110010000010111000011101011100110111011100010000100010101001100011000010000010010010000011001110100010111101101111110011000011110000011000000101001011000101010001001011;
#1 $display("%b", po);
# 1  pi=207'b100000001001110101100110101010001111110100101010101011111001100101111010110011100000101000111010010100100100111001000110101001101010000001110001001111100111111010001001101011110001111100100110011100101000010;
#1 $display("%b", po);
# 1  pi=207'b101100110000100111001100100100110101100011110001011100000010101100100111101111001101100100001011100011111110000111001100010001011101110000111000111000110011000100010000010011011110111001110110011010000111001;
#1 $display("%b", po);
# 1  pi=207'b010011011010011010100010010010001001010011000100010111110111101101000111110111101101011101110110111100101001110101100100011111000011110000111101010101101010011001111110110101101110010111100101101111011110010;
#1 $display("%b", po);
# 1  pi=207'b001110000111001111110000111001010110101001000110110110011010011001111111111000011111101111010001010101100100011011010000101111010010110010110000101101010101010101100100100101001011000011110101100110101010000;
#1 $display("%b", po);
# 1  pi=207'b000001000111011110111001100001101010000101100001110011000011111010000110111111101101001011100001111111001111100111100010110100111001010111100010110111000001111010001010101011100111001000111011100110000111110;
#1 $display("%b", po);
# 1  pi=207'b001000011101100100000011000001111101001111011101100000110100110110000101111000111010011010110000011100111011011011001100000000111010110110001010000110011001101001111011110011001011110101010100110111100100111;
#1 $display("%b", po);
# 1  pi=207'b110001110111001101011101001100111000010011111000000111101011000111111010001110010000000010110000100001101110010110010111000111100110110110011001011111110100011001111000000100010000111000010111110110101010111;
#1 $display("%b", po);
# 1  pi=207'b011110001011000010111110101000101100100001110111101100001111010011000111100111011100011001110010111010100100001101110010110001000000000100011110111011101011000101110111001000011110101101111111011110010100011;
#1 $display("%b", po);
# 1  pi=207'b001001110101010000010001010110100011100101101010010100001110100101101011001101011111000100011110001100100100011101000110011111110101111011101010111111010010010010111010001000101101001001000011101001000110111;
#1 $display("%b", po);
# 1  pi=207'b011111010101101000110101010100100010100010010111101101110000111000000000010101111001101000100001111000011111100011010110011100000111000100010011111101100001100100010010000100000010100001001100001001110101111;
#1 $display("%b", po);
# 1  pi=207'b000010001001101111001011100010011101010101111001101101100100101011111101101011011100010111110001000110001011110011010101101100011010110011000011011110110111001001101001001010011000111011100000010011011100110;
#1 $display("%b", po);
# 1  pi=207'b010001001101010111011110111000100011110000001110100011100111100110101010100110111110101001010001100000101011110011101000111000000100111100100100110001000110011100000110100110111111111110111111100000000000101;
#1 $display("%b", po);
# 1  pi=207'b011011001011110110111100100001110110111101011111010110010100101010001011010000100001111010101011001000001110011001000000100110010011011111100011100011100100001000110111011000010110000000000010010010000101100;
#1 $display("%b", po);
# 1  pi=207'b100001000011111011101100100010101111000111001100100011000000101101010000010001100110100101000000011001000001110111001111111110111001010011111010101001010010111111101000010000011101000000111001100010010010000;
#1 $display("%b", po);
# 1  pi=207'b011010010111101111101111111110111101110001011111101011110011110100110011100101010010100010001000011100101011100111011101100000011011101011100001101000010110001010110000111100011101100111111111011001001000100;
#1 $display("%b", po);
# 1  pi=207'b000111011010000001110100000011010111100100001111101110010010000101001000010001001100110001000001100001101000000110010111011110001001010100100000101000100101111110100000001111011011101111110010111010110000110;
#1 $display("%b", po);
# 1  pi=207'b101000010010011110110110000100111010101111100011110101010101001101101110000110111000010111101000010010101001011110010001100001100111001011010100111100001100010101000010101000000110100010010101011100011010000;
#1 $display("%b", po);
# 1  pi=207'b110000011101000000100110110111100001000110101111001001001011101000001010111011111100101001000011101011101110110000011101110111011011110101101010100101110001100000110110010000011001111101000010010001000011010;
#1 $display("%b", po);
# 1  pi=207'b100011000000011111110111111110010001010011111001101001110111011000010111011100011010111001000001100100111110110001101001000110101010110011001100100100000010011011100001101000000001101111000101111101111000101;
#1 $display("%b", po);
# 1  pi=207'b010011101010011110001000001101011010111110001010101111110011110001000100111000101000111110101111101000010011000111111100110000100110100000010101000111100001101000010111110010110110111010010001111110100100010;
#1 $display("%b", po);
# 1  pi=207'b011000111010011111000010010000011110100001100111110111101100000001100101000010100101111011111001100011110010101001000000101001010101010011101111011100010010111101111100100110101010000000110000000101010000001;
#1 $display("%b", po);
# 1  pi=207'b000111101000100110110000000000111011010000010001110110110101011011101011000010010011100010010100101011011100101010111001001101100001100001000001111100000000110100011010001010100001010101001110101011101101110;
#1 $display("%b", po);
# 1  pi=207'b100001110010111101101101111111110101111011110010000011011110000100001101110011110101010010101111000111111110000010010101110000010111011000011111011101111011100011110010101101000001100101111111010000011101110;
#1 $display("%b", po);
# 1  pi=207'b100000101001101100111111111000100001101010100010100000100111101101010110101001110110001101001010110110111100011100100000010111011000111010000110011111001011101010101101110001101110000110110101001000011100101;
#1 $display("%b", po);
# 1  pi=207'b001000001110100011010100000110100010101000100110000011011101000001010010111011111110100010110111010000010111001111011000100011000110110100111010011000001001110100101010110001001011010001111000011011001000101;
#1 $display("%b", po);
# 1  pi=207'b100101011011010010011001010000001010110100110110111010010010111001011100111110010001101000100011100001110110010101101010011110011000100100010011111001110100101111011001101001010011110101110000010000000010010;
#1 $display("%b", po);
# 1  pi=207'b101101110101101111001111110111100001001010011011010001101110110010010011110100001000001110011111100101110000010111100101110100010000011110011100101001001000001011001000000011111111001101100110100001010111000;
#1 $display("%b", po);
# 1  pi=207'b100111110101010001000101011001001001100010100100011111110010111111111010011011011100110000100100011101001010001110001100110011101000111110011100101100011001100001000101101111011101010101010010101001000100010;
#1 $display("%b", po);
# 1  pi=207'b100100011110000001000001000101011001101100010000011011000010100100000001101000000011011111110101110101110000001111110000010101000100011001110101110111010000111011101100000011000010111111100100000101010100011;
#1 $display("%b", po);
# 1  pi=207'b000000111100000100100101101101100101100101011110101110110111111100111000001101100001001011000101100011100000101100110001011101011011100001010111101001111000101110111111100000010010011000110110001101111000010;
#1 $display("%b", po);
# 1  pi=207'b011100011001011111011010000100001100110000110010001111010100011111010101111010000111101001101000111111001001000001011011000000111010100001010010110001110111111010000100110101101001011000011100111110101000101;
#1 $display("%b", po);
# 1  pi=207'b110111101001111011010110010100011011000011011110001101010010100100010101010011101101110100000010010101110100101110110110010101110000110100011000111111010010011010000010000000000100100011101100000001110111000;
#1 $display("%b", po);
# 1  pi=207'b010010111101100110100000101011000011110100101110111001011001001010101110000010110001011010011000010101100100111110111001111000001111110100011110011100101000010000110001101000110110001011000000010111110101101;
#1 $display("%b", po);
# 1  pi=207'b100101111110100100001110110000011101011110001000101011011001000111111000000110111011010110001001110111011111110000111010010100110010110101000000011000010000001101001011100000000111010111110110100100100111110;
#1 $display("%b", po);
# 1  pi=207'b000001101111110001100011101001010101101101011110111011011010010000010000010001010100111111110111011010111100110010000001010101011100100000100010110001110010010001101000011100010101110101001001100010010001001;
#1 $display("%b", po);
# 1  pi=207'b110111111101000111111101000001000110100010010001001001101100001110010011110000111011110110111111001001110111100000011001011100100011011100001010010111001001110101011000110101110111011010010101100100001000110;
#1 $display("%b", po);
# 1  pi=207'b001011101000011111001101110111011011000001011000111111110101111011110000010110110001100101001001110100010000100110111110100110110001000110011010001111000101001011100111010010101110110010001111010101011000100;
#1 $display("%b", po);
# 1  pi=207'b001010011111111100001111010110001000001100001010111011010110010101001110111110111100011011110111110011101010110101100101101000101110011011010010101101010111011111101111100111111001101100111110001011110100001;
#1 $display("%b", po);
# 1  pi=207'b110100101001101011111000101001000001010011111110111100000110011111011001001101001011011001100000001000101000101111111010000000111011100011001110110111011100100101010000011111100010010101010101110110110011111;
#1 $display("%b", po);
# 1  pi=207'b110011101000010000111111100001110101011011010100110000101010100111011100111110011111010100110010010100101100011001011101101101010010011100101011111001010100110101111101001110100011011000110100010011010011111;
#1 $display("%b", po);
# 1  pi=207'b011011110011101110001000000010111110101100001000111000101101000011010010111001011110101000000100111010001010110101010101110111101111011100010000101000011010010100111010101100010000001011010011111000011100101;
#1 $display("%b", po);
# 1  pi=207'b110110100111000000000101110101101101101110001011110100101010101001001111111101110011100000101001101111100001011101111101101100010001100001010000100110100001100110011010100001100111111000111010101100111101000;
#1 $display("%b", po);
# 1  pi=207'b010010001110101100001100001000011101011100000000111001111010111010000110000000100001111011110100011001010001011101000010110011101011100100101001111111111100101011110100010000110000001010000000011010101101100;
#1 $display("%b", po);
# 1  pi=207'b110001111100110000110111110111101111100110011100101101111101110111011101001001001000010100000100011000010000001001011000101110010111111101000111010010011101010011110011110000010111100100010111110011111000111;
#1 $display("%b", po);
# 1  pi=207'b101000110101101000101110001000011100100000001100111000101100111000010000101000111001101111111100101101011111001001101100010110011011000110110001111000000000110100010000000110100101001110101010101001001110111;
#1 $display("%b", po);
# 1  pi=207'b010110000110101010111010011101100101001100101010010001101011110010101100101101010100101110100100111000001011001000010110111101011111010100001001100000001011110010000010100001011001110101101000010011011010111;
#1 $display("%b", po);
# 1  pi=207'b110010000101000001101110010110110111001001111101000101110110101110010011110001111000001000101001110110111110011011010010000001110100100111101010111101101010000101101110100001010001001011010101101001010101010;
#1 $display("%b", po);
# 1  pi=207'b000111111110100011100110010110101000110101101010000110010011110101100101011000001010010001111000000010010011100100011110010001101001100010111010101100101000001110110101000000000011100111101010100101001001110;
#1 $display("%b", po);
# 1  pi=207'b111111101110000111000011001010111000010000111100111111111011010001111001101110110101010101110100111110100011111100011110110110111110010001000110001110000010100010110011110110100010101100010111100010100000000;
#1 $display("%b", po);
# 1  pi=207'b110100000101100100110011010000110111010100111111001111101110100011111000010111111110101101111010000010011100011011001101110111010101010011110000000110011000010010011110000101111100010000100111100111110111001;
#1 $display("%b", po);
# 1  pi=207'b011110010000000011101110000100111101001101101101001010000001111000001001101111000100101101001011010110011000010001100110011011000110101100011101001010111010010100010110110101000101011011000011011011001000101;
#1 $display("%b", po);
# 1  pi=207'b010001011010100111111011110100100110010001001100011010111010111101100011001111001000111011010100001111111110001000111001001111010011001101110101011011111011010100110110110110010100100001010001110011111101110;
#1 $display("%b", po);
# 1  pi=207'b110111010011111001110111011010110010100010010100001010011111111001010100001100100110010101111000000010100011110100110001001001000000110010100000110000011010001000100001000110001101111111110000110010000000100;
#1 $display("%b", po);
# 1  pi=207'b001100011100011110101000010101010101011011100010110010000110101110000001000111101111000101111110101000111111000000100001100000011110010010110111100001011100100000101111101011101111111110000100111100110011011;
#1 $display("%b", po);
# 1  pi=207'b100100011010010111101100110100000110011101111010000011011001000110001011111100001011011100100110001101110001000011101000011011011110100111101111000101111011011111000000100100011101001001100110111010011011011;
#1 $display("%b", po);
# 1  pi=207'b101010100101010101110111100101011100101110010111001111101001010010100000011100100000100100101001101110100010111011011100101011101100110110110100000100010101001101100010101000000010100000011011110101010001001;
#1 $display("%b", po);
# 1  pi=207'b011101100011011000011011110100101100100000010111110110111010000011101000000001000000100111110110101100101110110111110010101001110101111110001001101011111001001101010010101000110101011101001001100110000001010;
#1 $display("%b", po);
# 1  pi=207'b101101111100111011000111011101000011111001000111000010000000110101010111100111110101000011001010110111000101010101100110101001011001100100000111001110001100111101000010011011001111111010001010010001001100001;
#1 $display("%b", po);
# 1  pi=207'b001000000000110101011000011111011000011110101110011100100111101001111110000011000111111011110101000111110011010111111010111110011100011110110100100100111000100000001010110111100110001001011000000100110001101;
#1 $display("%b", po);
# 1  pi=207'b110110100110001001101010000100000100011111101110000111110111000010111011000001001011101000111000101101011111000100000100110110101110111110010011110010101010010011000100101001000011011000011110010011000101011;
#1 $display("%b", po);
# 1  pi=207'b011111000001000000010100101111010110010000110011111110001101010000011001111110010111011011100110000100000110110010100011101110111101010110000100011010000000100111100111111011011101001010101100001011101110000;
#1 $display("%b", po);
# 1  pi=207'b110101100111100100011001010100010001010010000010101110011101110001101110001110101011100001100000111110101001100111001100100111110011111011011111110101000010011010111101100010111101111010100100100001101111111;
#1 $display("%b", po);
# 1  pi=207'b111010100110101111101110000011100111110100110010111101001001101011100001111110101000100000000011000011101011111111101100110100101100000100011011000100111011001010100000100101100100000111100101010100101100000;
#1 $display("%b", po);
# 1  pi=207'b100111000010010111110111100000100000011011100101010010100011000100100100101101011010101110000100111111001110011111000001010011110110000101111001101010001001110001011011000011001001010111001011001101011011101;
#1 $display("%b", po);
# 1  pi=207'b110100000000101010101000111110000000001010111000001010001010001100100111100100000000111101001100111001111110100100000110110111110100001111010100101000111010100011100111000101010011111110001100011110010100101;
#1 $display("%b", po);
# 1  pi=207'b111100010010011001100011010111010110110001101100101110100011011010100110111111100001010101011000000000011100101111011011100001101111000011110001011111101110101000100100001100111100010101101010011100111110000;
#1 $display("%b", po);
# 1  pi=207'b010001111110101111011101010111101001010100010001010001110001010111111101010010001110001010011010001011010110111010001111101001110110011001010001010111000101100100000100100110000101000111100000001011110011111;
#1 $display("%b", po);
# 1  pi=207'b000101011010100011001111000011000100110000011011111011000100101011011111101100110001011110111100011100001001111010101011110000111111100110001010100101011010110101110000101011100010010010111111110110100111001;
#1 $display("%b", po);
# 1  pi=207'b100100011110011110000010000100001101100001001000111000011110001011011110110100001110010011011110011101001010001000001101100011101001010101010000000010100100010010010100011110111011110110100100001010001001010;
#1 $display("%b", po);
# 1  pi=207'b010101110010001101100100011000100101001000110011100001001101001001000110100100001010101101101100100101111101010011010100100011101100111101000010110100001000100101011111000001101100000011111000100100011100100;
#1 $display("%b", po);
# 1  pi=207'b111110111001111111000001000010011111100001111100010011100111000001111011110001110110000011100111010100110010001101011000100110010101000100100011101101000000011001010001010101001100000000101011100001110001000;
#1 $display("%b", po);
# 1  pi=207'b110110010110101100100101011010111111100000000001100101010010110110110001100101010110100110110111010001000101001010000111000010110001110110010101101001010011111011101111011100000110101001000001111110001010100;
#1 $display("%b", po);
# 1  pi=207'b110101110111000001100000110111010110001000100000010011111001011110110100100010110000000100000000110101111010101101101101111000000010011011011001000111010101001110101011101101110110101101110001010110010011110;
#1 $display("%b", po);
# 1  pi=207'b011110010101101000010111110111000101011011110101010110000000110011110010100011001101001011100011111101001000010101100011010101111000110100111010111110101010111011000101111111001010100010000010110110100011000;
#1 $display("%b", po);
# 1  pi=207'b100110001101010101110010110101010000011010101011000110110111001110111011110011010100101101010110000111101110110111000001111110101000101101101111101011010110000011000101000001111111101011011011101011000110000;
#1 $display("%b", po);
# 1  pi=207'b001000111100000101101001011011001101100011110011001110011000100110000001100100011111010001011010100110001001101101111000110100000010010110101000100110011001011000110100110011001010010000011100011111000001001;
#1 $display("%b", po);
# 1  pi=207'b011100110010000100100011111100100010011000010011110011100010011110001000010000110100000110101111101111010101011010001010100101111011101000101101100000010101110101100010111001010111100110101000101100010100000;
#1 $display("%b", po);
# 1  pi=207'b111011101010000111010010101010101001110100011101100111110111111010100011101011100001100100011001011001011011001011111010000100101010111010010001111101110010010100110001111101010010110000110010111000110101111;
#1 $display("%b", po);
# 1  pi=207'b001101001100100011011111001011000000100100001111101100110100101010111110011111111001011000000010010001010011011011000001010011111010110000000111101010001111100001011010011100111110100100010110100101101111011;
#1 $display("%b", po);
# 1  pi=207'b000010101110110011111000111111001000010011111000001110101100001011000000111010110011011101010110100101111101011011000010000101010110000000011011110010110100001100000101100100101000010111001011011101001110101;
#1 $display("%b", po);
# 1  pi=207'b000011100101010010101110001100001001011000111000111111010001101101100110010110000100001110100110001110010010101111101001010001100100010100100010100000000010011010101111101100011010011110110111001010000001110;
#1 $display("%b", po);
# 1  pi=207'b010010001110011011011010101010111011011010000000000111100001110001101010100010100011011100010100001110011101111001011110101110110011110110000011111100001010101101111000100111010111111010000001001111110100011;
#1 $display("%b", po);
# 1  pi=207'b010011011010111001100010100101110100000001100011001010100101000000010111111101111110100001010110111101000111101100001011010000111000001101111000010111010110000001111010111101110110111111010111110101101000001;
#1 $display("%b", po);
# 1  pi=207'b011100010100101101101011011101010110101110100110001110000001111011001101100100010111100001111111011011010011010100011001100011101011010111000110011101111011101101110101011111000100001100000101111000110001000;
#1 $display("%b", po);
# 1  pi=207'b110110000001111110100100000101100101011000000001010110100100011011101010111100110110100001100001100011111110111110100001000010111001010011001111010111110100111001110000010100111110111011010000100010001111100;
#1 $display("%b", po);
# 1  pi=207'b001110111101010001111000100111100010001011011001010010001100101100100111001010011111000001101111100111110001111111101111000110010101111010011101101011010101011110010100001111000001100111001110011000011011101;
#1 $display("%b", po);
# 1  pi=207'b100111110110000000011011111000111011100111101100000011110100111011011000101101001111011001000000111000110011100101101100000011000001010111011010010001100001101110100110111011000011111010100101001101101101001;
#1 $display("%b", po);
# 1  pi=207'b111010101101101010000000110000100000000000101011001011110110100100100111100011111011001001001101000110011011111111101001001110111011000001101010010101100011001010011001011111001100001111001011100000111011110;
#1 $display("%b", po);
# 1  pi=207'b000101010011010111001111000010011100110110010011010101101001000111100100001111101100110000110011111100111010001100000010101100100111100011110100001101001100100101111000111001111010111100101110111000011100101;
#1 $display("%b", po);
# 1  pi=207'b100011111100000100101010110110011001110001000001111110010110101000001111110000110011001110100010100010011010010110011101110101111001101000100011101101100101100000110100110111011011000101101010101000010001110;
#1 $display("%b", po);
# 1  pi=207'b110111000101010100101111101000001101001000100001010010100011110000111101011000011100100011000010110011000100110011101110101001110010010010101111101011110110110111110011110001010111101001011001001010111111001;
#1 $display("%b", po);
# 1  pi=207'b001001001101011001010100100010011110000000110100101111111110100111010111000000011101100111101011100001101110011110100100111100000010000100100000011011110110010000101101010011100000011111001101001101011110010;
#1 $display("%b", po);
# 1  pi=207'b110100010101010011011010000010001001000010100011110000000110101110011001000000011011110110000010100100101110100010101100110001000000000101000100101010110011100000000101110010000111110011001110001100011111010;
#1 $display("%b", po);
# 1  pi=207'b110011101100000000100001110011111100101001011100101100111011110100100110010010101111011000011011111000001100101110101101001100101000011111001101001010000111101111111001011011000001010101100001010110000101110;
#1 $display("%b", po);
# 1  pi=207'b100000000011001011100000100111010110101001111110010100111010001010100010101010010110101100111011101111000111001010110000101111011110101000110001010000000000110100000001000001011100001100000110010110011010000;
#1 $display("%b", po);
# 1  pi=207'b111011011101110001111110000100111011011101001110000101010010000101000110101100001101100011101011101010110100110111101001011111001000100000011000101011000000101001010100111010100100001001000101110000001001000;
#1 $display("%b", po);
# 1  pi=207'b011111011100100110010110101100100100011110100100001101011011100101001111001010010100000010011001110010000001011010111101100101111100000000111001111001000101111100101111010010010110001101110010011111101110011;
#1 $display("%b", po);
# 1  pi=207'b000101110001100000101110000010111110011011001101110100111011110000111101110000001011110111110111011110100100110010100110101000011111111011011010001111010101100110011011110111101111010111001001010010010000111;
#1 $display("%b", po);
# 1  pi=207'b001000100010000000011110010100110001100010111001011001101011011100111111000010011001111101010010110111010111011101110000010011100011111110000011001011001101000011110010110011011111110110100011101101110110110;
#1 $display("%b", po);
# 1  pi=207'b100011110011001100110101000110110011101001110000111110111101011110011010101100101001101000100100111101100001001000111010000100010110110111101111010000100100011010111010000010100001101011011101110111100010111;
#1 $display("%b", po);
# 1  pi=207'b001101110111110000111001100111110010010101000111010011011110110111101011011101100010110101011101000111111001011101001010000111110100001011001100110111101000000011010100111000001011001101100011010000111011000;
#1 $display("%b", po);
# 1  pi=207'b011110011011011100110010010110101000111010010111010001100111100011100101100011100011000000101010010010010000111100000110111101011001000011100000101010010111110011001110001000000111100001100010010110010001000;
#1 $display("%b", po);
# 1  pi=207'b001101101010001100000001111101110010111000111101001011100110100010010010100100001101101000000101011100001101001100001100011011011110010001111011111000010010101100110011110001010011011011101000100011000000011;
#1 $display("%b", po);
# 1  pi=207'b011100000000111010011010100001110100001011111110010101001111100001101110001101100110110110000010010010111011100101011001111000010111111001001111100010010011101001011101010100011101111001000010110111101001101;
#1 $display("%b", po);
# 1  pi=207'b011001100011011111011101101111110101110001110011000000000110111111000001100111000100101011011111110101011010010101010111101001111001010110111110000011001100101010010111111100111100010010001110100111001001001;
#1 $display("%b", po);
# 1  pi=207'b001101001100110111101100100111011000011110101011011111000010101011011111001000110010010001111110111110011011111010100111111100101110001011101101001011101001000010100000111000000110101000001110000100100000110;
#1 $display("%b", po);
# 1  pi=207'b101100000000111110110110111010011010100110111110000110110001011101001101101001001001001111111111010100101100100000111001110101110101111110011001010000100101010010011101011000010011010000000100011010011100100;
#1 $display("%b", po);
# 1  pi=207'b110100101101101000111011110110101000100010101011000011110011010111101001111001000011101011001000100001010110110010111001001100011111111000001001111010110010000101001011001101001011000010011010011001111010000;
#1 $display("%b", po);
# 1  pi=207'b111010100101000010111110001000101101011101001011001100101011000111010100111010010110011000100000110011101111101010010110101011110100000111011101100010111101111111111110010010011001000100000110111110101110101;
#1 $display("%b", po);
# 1  pi=207'b001010111100111011101100111000110011101010010010111010010000001111001011010110100011110101010000000001110101110111100011011011101111100010001110111111110000001011101011110100101000101101110010010101100011001;
#1 $display("%b", po);
# 1  pi=207'b100100000000110000111110101100000101011000010000110101010111010000110110110101111000011000110000101010010100110101010101100011100100010110000110111010101110010101010011010001011011010000010010101011101110001;
#1 $display("%b", po);
# 1  pi=207'b000000001011101010111000101010011101010111010011100110111000001110101101101000000001010001000011101100001101110011111110110111001011101000001100011011110100000001000110101100111100001100011001110001010111001;
#1 $display("%b", po);
# 1  pi=207'b000100111010011000001011101000000101000001010010101001110011001001100011100011001001011100110001010010010000011010110010011111100010010100111110101101110010001011010011110100111010100001010000001110001011001;
#1 $display("%b", po);
# 1  pi=207'b101101101100111011011111001111000100010001110100001011001110010110010101100111000111010110010111110010011110110101110010011010100001000100011110010001111000001101010011111100101101000000001111110011101001111;
#1 $display("%b", po);
# 1  pi=207'b000000011001100000011000001110011101111100111001111001101101110110001101011000110101111001100110110001110111110100110101110101110000011000011100001011011001001010011000001100001011110101000000111011001000000;
#1 $display("%b", po);
# 1  pi=207'b001001010101110001011110000100110000110000110011011011101101011000111110011110000110100001110011111011000001011001110000101000000101010011001100000011010110101111101000010011000011101000011101000011111110101;
#1 $display("%b", po);
# 1  pi=207'b001101110101010111000111100011000100101111100111110011111000010101101010011011011011100010001101100111100111010111100100001110101010111100011111110111100101100100000010111011011011000111010000100010111101000;
#1 $display("%b", po);
# 1  pi=207'b110110101011010110100000011101110011111111011101100001111000111010111111011010001101000100010011011111001100110010010111101010011111111101101111111101011011101111111011111000010011100101111100100100000111111;
#1 $display("%b", po);
# 1  pi=207'b011011101100010001110000110000000110100001011001110000110010101000010101100010110000000111100100110101110000111100010011000100000000101001110011101011010010011110010001111001111000111010111011110001111001001;
#1 $display("%b", po);
# 1  pi=207'b100010101111100010101001011011101010001110001111011111011100011101100100010001000111000111011011111000110101110110001100100000000111011001010101110111011010101010001011110110010001111101110011001111011101100;
#1 $display("%b", po);
# 1  pi=207'b010101100110111111101000100011001100001111001101111111100000110010101101001000000111001001100110101111011101010101001011010011010111000100011101100101001000010110000000000101100011011011010000001000011000010;
#1 $display("%b", po);
# 1  pi=207'b100001101100100011011001011010110000010100100011011101011101111100001000010101011101110000100011111110000101101000001001101010001001001011001001111110111111100100000101010000111000101000110010000110100001111;
#1 $display("%b", po);
# 1  pi=207'b011110111010110010011000100111001111101011010110100100100110100110010010001011101111101111010110110011000010101100011111001000101111111011101001000011000000010010100010101111011011111100101100111000110100111;
#1 $display("%b", po);
# 1  pi=207'b110101010011111110100100001000100101001100101011101011101101111001101001110000000100110111100011011111101111101011010110001000000110100110000110101100100100000110101001110001000001100000100101111100011010001;
#1 $display("%b", po);
# 1  pi=207'b011010010100010000000011011110010111110011000000011010010010100100000111110001010000101000101010011011000000011000100010000011011111100001010111001011010001101101010101100111100111101000010001001001001101111;
#1 $display("%b", po);
# 1  pi=207'b010100110111010101110111100011101110101111001110110100000111001000011000111101001111011011011100101010011000011111100101110101001010011111100111111101011001101111010001011011101110001110011100101010111001001;
#1 $display("%b", po);
# 1  pi=207'b110011111011011110010011100100110011111000100001110001000110011010011100011001110111100100100000000011011111000011001111100100110001101000100010110011011001000001111111000101011101000001001001111011100101111;
#1 $display("%b", po);
# 1  pi=207'b100000100010111100111010111111110100010001101011010111011111011101111110100000111001110011110001111110000010010100110101100001111100100101001001010000110111010111110010001100110100001110110011010111001011011;
#1 $display("%b", po);
# 1  pi=207'b111000010101110100001110101101111011101100110011001000110001001010110010101111000100100110110101011100001101010010010001000011101011010011100100001000010110100010100111101010010001010101000000010001010100100;
#1 $display("%b", po);
# 1  pi=207'b001101110000011000100001110110111001100111011111100011111111111011111111111111111000100011001001100011010000010100010110101101010001100011000011110000101100001000111010000101000100010101111001000101000110010;
#1 $display("%b", po);
# 1  pi=207'b101010100100100010111111100010100100010110111010001010111001101111110011011110000001010000000111101000111110011110011000100111001011000100011011101110100000011001010000111000111001010001110100111111111111111;
#1 $display("%b", po);
# 1  pi=207'b101101111101110110110000100111011011110110111001100011001101101001110010000010111010101000001111111011110101111011100000101010001001110110000110101100101101000111010010000111000101000000001001001110111111111;
#1 $display("%b", po);
# 1  pi=207'b111101011001101111001001101000011111001101110111110100110110011111100110000000101011100001011011110101101111100001001010100011011100011000100100111100101111110010001010111000111111111001000001000100011110000;
#1 $display("%b", po);
# 1  pi=207'b110001110011100100000110011010110100110010100101110111011011011101101010000010001011011001100101000001100111000001110110101010010100110101000001100011011010001011000101000010101111101001010001001011101001100;
#1 $display("%b", po);
# 1  pi=207'b110100110111111111001010000001010110101101001001111010100110100100111110111101010000100001100000000001001011110010000000100010010111100011001101110110100110001100010001111000010101101011111001000110011010111;
#1 $display("%b", po);
# 1  pi=207'b011100101111101110101111101010000110010100011111111111111000110101100101101000101100000100000001100111000101101101010011000011000101101101000001110010001000110101010110010001010000110000001100101001100000111;
#1 $display("%b", po);
# 1  pi=207'b000100001001110110010010011101111000110000011111011100010111010010000110101010110111010001000110001111101010001001011000011000111001000010111001101010010000110001011111100011001101100110000001111111110111000;
#1 $display("%b", po);
# 1  pi=207'b000010111111010100010000101110000011000010101111001010100101000111001011010100101010110011100001011100011010111110010101111110001011000011010011101111110111000111010001111010011010100110001001001101111000001;
#1 $display("%b", po);
# 1  pi=207'b111010010110001010100000011111110001010011101110110100011010010001010101111001010011100100010000101010000101101000110000011100001001111011111110010001011011100011011111100010100100001000101100011010000111101;
#1 $display("%b", po);
# 1  pi=207'b101001100111011100011111100101111101100101001100101000001001101001000010111010001100010001101010111100101110011011101111001010011010010111100001101011000001000111110100001111011011110010000111101011111001001;
#1 $display("%b", po);
# 1  pi=207'b011101000000101101111000011100011001111110001100000010111110000101000011001110011011111011111111001111000011111101000000000111000111101001010000101000001100011000011001111000100000111110110010101011111101111;
#1 $display("%b", po);
# 1  pi=207'b011111010011101001111011011000101010110110111001001001100111111001010011111101000001100111110000110001000101011101101110011011101110010000100010101010100001101111110101001100010101110110000110000011100000100;
#1 $display("%b", po);
# 1  pi=207'b000000110001110101010111000010001110101000110010100001111101110010111100100101110100001101111000000111111011101000111111011010010110010100011011000101001111111111100101011010101000001010100101100011010011101;
#1 $display("%b", po);
# 1  pi=207'b001000001101000001111001100100111000011010111001110000011001111010111100110001001001010101100111110011010001011011110001011011010001011100001111110001100100100011110111011110110011011011111101101100100011010;
#1 $display("%b", po);
# 1  pi=207'b011010001101000100100110010011000111001100001000101111000100110010111100110000001100100000000000010111000011101110000001000000010010001011010111101101110010010100111110111010001101000010111010011001100100000;
#1 $display("%b", po);
# 1  pi=207'b011101100011010111100011100100001001001110110100110111001010111110000100110110101001110000111100111100000000001011101110100001101111110011011100101010000011101100010001001100111011001111111011000010110011111;
#1 $display("%b", po);
# 1  pi=207'b011001110001110001110000000111010101001100001010000000100111011011010110101101110001011100000000100111010101011001100000101100101100001111101111110101010100110111110001001101110001110000111001111001011100001;
#1 $display("%b", po);
# 1  pi=207'b010110010011101111110110110111010111010011101011110011111111000100000000101101001111001111100001010110010110011101011111010111010111001000100110111110010010000000011100010000100001110001100000110100101111010;
#1 $display("%b", po);
# 1  pi=207'b010100001111011101111100101100111111010001110101000010111101110110100101100101111110000110000101110110011001000111100000101111110010100100101001011111110100011101011100100011000101111010000011100101111001111;
#1 $display("%b", po);
# 1  pi=207'b000000101111110000011010011010000111111110110110011101010000011110110110100110011011110101001001001001001100101101100000001000000101011111011000110001100001110001110010000000111100110010110010100100110011011;
#1 $display("%b", po);
# 1  pi=207'b111111010011100101110001111101110010011001100010001010100011101100011010100110001011100001001110111110110010000101001010011100111011100101101100100111011111101001011111101001010000111011000101011000110001010;
#1 $display("%b", po);
# 1  pi=207'b011110111010110100011001111101100011001100110100000001100100110001010110100001111100100111110101100001000000001100011010001101001011001101011001111111010010111101010010010000100100101110110110001111001100111;
#1 $display("%b", po);
# 1  pi=207'b001000100000100000101001101110011100110011001011010000010100100111111101011001100110010001110110000000110000010010100001100110100000011100100011111100010101000001011101011001100110010000110001111110001000001;
#1 $display("%b", po);
# 1  pi=207'b010110001100000100011111101011110011010011001010101111110101010011110110000001011110101111010010110100111110011011110110100011111101001001010011001111011001001010110000010010000000100011000101110110110101001;
#1 $display("%b", po);
# 1  pi=207'b110000110010010111111011100111101011010100111101111100010011101100101100101111100110101110010111000001011110100001101101010100100000101000010111011100110101001101011101000010100110000010110000011111000011101;
#1 $display("%b", po);
# 1  pi=207'b101111001001110111001000000111010101101001000110110100100001101110001010011100100000111101101110111110000101101000011111101001111001100000101001011110101110100001100011101110110011101011010101110001110010110;
#1 $display("%b", po);
# 1  pi=207'b010000010101100011111001001010011110101011000101110011100111110111101101000000011101110010101011011111000101101010011001000011101011101101010010010101011111001000001110110100111011000011011100011011000110010;
#1 $display("%b", po);
# 1  pi=207'b100110111111110110011000110100000010111111000111110001100011101001001110011000111111111110010011001010001010110011101111110011100010001101000011101110001011000011001001110110010010101111000100010100100010001;
#1 $display("%b", po);
# 1  pi=207'b101111011000001010000100111011001110001101010000100100010101111101110000110011001000111010000100101110110110101011100111000111010000011100100000000110111000100010110101111010000100000101001101100000001011111;
#1 $display("%b", po);
# 1  pi=207'b001110011100100111110110001011010001111001111100111100000110011001001010000110100111110000110010011100010010110001000110110011000101110000101111001010000001011010000010011001010010111000010100010101110101010;
#1 $display("%b", po);
# 1  pi=207'b100111000100011101011001111100111001111101100101010010010001110010110011011110110111101100001000111001101101001011011101010001110000001100001100010000100101101101011001000101010100110110101010000001010011100;
#1 $display("%b", po);
# 1  pi=207'b000011010001111010001010111111101010010110010110010001111001111111111010111101011010011100001000011100101101110100111001001011110101010101010101111011110111010010011100100000011100110000001100100001100111100;
#1 $display("%b", po);
# 1  pi=207'b101010111010001001110011100011011010110110110111010110101000110110100110011111010110001001111100100111100110001001011110110101111101000010001010100110100100000110111011100011001100000100010011011111000101110;
#1 $display("%b", po);
# 1  pi=207'b101111011011110110111111101001001111111110111110010111000010011100101011101100110111011000101101100110111000001011111111100110011110010111111001101110110101000110111111000010011011001100111100110001111011011;
#1 $display("%b", po);
# 1  pi=207'b101010010011011111101000010111011000110011011110110001101010010110011000000110100111101101001011011010110011001111010000001011100000100011111011110010001000011000011011000110101011011101110101101101101110011;
#1 $display("%b", po);
# 1  pi=207'b011001000101000110100000001110111100000000100101011001101010000111111001111111010011000110001001110000011001000001101010001110001011110110111110111101110000100011111010110100100111110110010111111111110011110;
#1 $display("%b", po);
# 1  pi=207'b001100001101111001011111110111011001001100011110101001011100111111000001100100101011011110000010000111001001011001000101111010111001100010110111010011010011100000000100100000101001001000101110111111101100000;
#1 $display("%b", po);
# 1  pi=207'b110000000110000100100101101101100110101110111111110010011100000110101110011011101010101011110000101001000111010100001001110100101001110111100001110100000110100000001001101111110100000001011000000000010001101;
#1 $display("%b", po);
# 1  pi=207'b110000101100010101101101000001000111001111001111010111011010001000111000001011011010011010100111010110011010000110101100000000001001111011101000010011011010010110110000001100010101000010111111000101100110010;
#1 $display("%b", po);
# 1  pi=207'b110010010000010110110100001010110110011000011010010110100101111001110010000010011100010001100010010111010111100101110101001101101110100110010010110000101101011011111101111010110101101101110111011001011110010;
#1 $display("%b", po);
# 1  pi=207'b111001010100001111010010010000100110000111001010011110110001110001010100001110110011011001100011010011010001001101100100001110001100001011010100010001000010110000001100101010111000001000111000000100011001110;
#1 $display("%b", po);
# 1  pi=207'b110000111001001111101010100101000010110111010011001111111100011000110011010101100011010111000000111011010101100100001010110110101111111100110001001100101001000001011100000011101110010001110010010001010111010;
#1 $display("%b", po);
# 1  pi=207'b010110001011101010101000100100111100110001110011110110001100010001100010000001000011001111110011111011101110101001110010011100101100000110010100101000101101101000000000001001110010110100101110001001101001010;
#1 $display("%b", po);
# 1  pi=207'b100011110011011011010001101011111000110100110001110001100011011001011110100001001000111010011110111101100110010001010110101100110110011000001111110100011010111010110001111010111001010011110010000000000011110;
#1 $display("%b", po);
# 1  pi=207'b011111011100111011111100011010111000101111011011101010100000001001000101000001010110011011010101000111011101111000101010111001100000000001010001010100010111001000101111001001101000111110101100010100111110011;
#1 $display("%b", po);
# 1  pi=207'b101101101010110001110000111000000001000100001000101100011111100101011001000011110101001111000001100100100010001110011011100001010010010000011000010111110101100010001001100011100111010110011100111100101101110;
#1 $display("%b", po);
# 1  pi=207'b001010001001111101100010010100011010011000011101011110010111100101010001101011001010010011100001100101000110110001110011110001101010001010101000000001010111011111111001111011011100101110101101100001100000001;
#1 $display("%b", po);
# 1  pi=207'b111011010110011000011001000000110101111000110010010100110000000101110010011000011001111111011101100011101010011111000110111010010011011111101011010001001001101010100011001100011101011011110001110110001111000;
#1 $display("%b", po);
# 1  pi=207'b100010110101010100001001100100010000001001011110110011100011100001111111001011011111000101011111100111101001010101000001110101110010111101100100110101100001010100000101001010110100000010000110000111000111000;
#1 $display("%b", po);
# 1  pi=207'b000100100110011010111100000100000111101100111101111111010000000011111000101010111000111111101100101110010100001010011000000110100101010010000100111110111110110110010100000011000011010010010010000000100001011;
#1 $display("%b", po);
# 1  pi=207'b001111010110000110010100100011001101111011010111001101001001110000110010001000001010111110100001011100110100101010011011101010000110000110001010000111101000001010010101000111100100110100011101011111010111000;
#1 $display("%b", po);
# 1  pi=207'b110000000000110101101000001010001000000100000011101111111001111101100011001000011110100000010101011010110110111111000011100011001111001111100111000110010010000101110010110111100010111111011110000100010110110;
#1 $display("%b", po);
# 1  pi=207'b011101111010100000110111100001111100001000001000001011100010011000110011111011000101011011011110010110110111110000010010011111100111100100110010100111011010111000111010010101000100111111011000111011100001101;
#1 $display("%b", po);
# 1  pi=207'b101101101100011000100000000101010001100010010101100110100011000001100011101111111110001110101100100100000000110100111011001011001000100010110010111100001000110000111011010010110100011100001101110001010001010;
#1 $display("%b", po);
# 1  pi=207'b101010011110110010111011011011010110110101001011001111110011011100010011010101011100100001010101100111100010011110000110111000011111011001001111001111010111110000101011111011100110011101111110111101100001100;
#1 $display("%b", po);
# 1  pi=207'b100101010110110110011001101000000010000111101101101101111001111010010101011110100111010010111000101011110101001001000111100011010010001010000011000010001100000001110101001011011110001010110101010010001100100;
#1 $display("%b", po);
# 1  pi=207'b111011010101100001010100111001100101000001111011011100001110011111111010100100101001001001011101101000110000000010001011001101010111001100000010011111110101010000010011011101001110001010000111100101111001010;
#1 $display("%b", po);
# 1  pi=207'b101101000111111100111111011001010010101110011110011100010101110000101011000110101001001011110010101001110011000111111100110100010011101011101000000110000101100001011001010110110101101100001010101001111111010;
#1 $display("%b", po);
# 1  pi=207'b110000100001001000110000000110011001000001010001101010011101100010100001111001110001100010100100001001001110001001000111001111110000100111010101001011000001010000001010010010001101011001011011111001110110001;
#1 $display("%b", po);
# 1  pi=207'b100111011001011011010000010000011100010010000100100100011110110000011110110101001110111110001101000000111111000101000001111111111010110011001011110100100111010110101100101101100010000110000101000000101110101;
#1 $display("%b", po);
# 1  pi=207'b001000100011100011001011110000101010100011011110010101111100110010110110111011111111110010001011001111001000100001001101100001011110100100010110111001000011000110100010110101100010000111111001001110000100111;
#1 $display("%b", po);
# 1  pi=207'b011010111100110110111011011100001100100001101011101010111110111110110100100000000001100001000000000000101111000001000011111100101011110110100011001110111100001111101110000010101100101011001000100100010100011;
#1 $display("%b", po);
# 1  pi=207'b001001100001011001001101100110110000110011001001100001000010100000100000101010100010101111010101101100010010001001111001001011011111111100111010011001011000110011000000101111110000000001110001000111001100011;
#1 $display("%b", po);
# 1  pi=207'b001101110101011100011100110100100010000010010111110100011010111000001011011001011011111111000011110010001001011010010001001100100101100110000011101100101111100101010101111000011101001000001011010110010111101;
#1 $display("%b", po);
# 1  pi=207'b101110100001101100000111001011000101000000010100011111001000100000011000101001011111110100000101100101100010001111000000110001010111011101111101111101110011100011101110111001110101101010111110000110000111110;
#1 $display("%b", po);
# 1  pi=207'b100101110000100110101000101000110101101001001001110011110110001001011000011001011001111000111111111111100010111010110101010101010100001111101110011010111110111110000000110001010101100000110100011001111110110;
#1 $display("%b", po);
# 1  pi=207'b110000111000101101011101011011000100011000001000000111101001000010101011110010100111110001010101000101111011111001101000100100110011010110100110000010101000110011110000010010001110111001100111010111101011111;
#1 $display("%b", po);
# 1  pi=207'b110001101001100001100100110110100101001101010011010000110111000111111000101000001100001111111100000110100001011010111100110101100011010111111101010010011111110011101000010001000101010100001100000011010110101;
#1 $display("%b", po);
# 1  pi=207'b100000000010000110111101100100010011101000011111010001011111111010101011100110010010010111110100111011111001000101100010100101001010110111000101001011001000010110000101100010000011100100110010111000000100100;
#1 $display("%b", po);
# 1  pi=207'b111110001110101110010001000100001010110000101011111110010001101001111111111010000100011010101100111011011001100110101111111000110110001101110011010110000001010010101110000011010100101000111011001001000111110;
#1 $display("%b", po);
# 1  pi=207'b101101101111100101001111000101111000110011000011111110000001101101011001111111011101001011010001001001011111110000110111111110110001101100100011010100111011000000000001110001011000000110001010100110000111001;
#1 $display("%b", po);
# 1  pi=207'b101100001101000001000110110110010101000101101000000100110101001010011111011010000001011010111101101010110100011000011000101000111100101101010100010100101100110011000111110011101011111010110100001011011010110;
#1 $display("%b", po);
# 1  pi=207'b110111111100001100111011010010011001010110011001101111001001000010100010010000111001101000101111111111001011101110000010011001101100100100101110001011111111100000110101111010100111101000101111101101111011101;
#1 $display("%b", po);
# 1  pi=207'b001001101001110000101101111000110100100100101111100001101000000101010011011100010100101011010100000101110011110101011110101100111111101110100000100011000010010101111011110001100100111110101101110001111001010;
#1 $display("%b", po);
# 1  pi=207'b010110001101001110101101110101010000101110001110001110010010011111001110011011100010111000110001010100000010100000111100100101010001101000101101000011100101110010100011100111001101110011010110000010011100001;
#1 $display("%b", po);
# 1  pi=207'b111111001001001011011011001110101110100111100010101010010011111110001110100001010100111000101101010101110110101010001010011010111000100000111111100100010100110111000010111011110000001011010100011000010001100;
#1 $display("%b", po);
# 1  pi=207'b010000100000111101001010011111100101110011001011110101011111011110111010111001110010110111010001110000101000111000100001101011000111010100001011000100100100010011010001011101100000000000010000110000101011100;
#1 $display("%b", po);
# 1  pi=207'b001101110111101110110100010000110011101101011100010101110101101000010010001001011101111110010100001100011010000100011000001010110000001011001010011001000010111011100110101000010111001100100100110100001111110;
#1 $display("%b", po);
# 1  pi=207'b000111001000001110101000100010000000100000001011000101001011001100010100010011100111101111100110110011100001101011000001101001100001001110010000011110110111110010001011100110110110110100110100001100111110001;
#1 $display("%b", po);
# 1  pi=207'b000101101000001011011010110010001001001011110011001001000101100010111001011001110101000100011110010010010011110100001101001000011100110100010001001011001011011111100111110110001100100100110111111100111111111;
#1 $display("%b", po);
# 1  pi=207'b100001100111011111011100010110100100000110100000100001001011110011000001111101111100000001100110110100111010010010000110000000111100000010101100110011111110110010001101010000010001101110001011011001010001101;
#1 $display("%b", po);
# 1  pi=207'b011110011101011110110101110111011110101111100000110101000111001111001010010010111101101110001101010100100011001111110110100011011101101110111001000000100111010011000011110100101101000110111111011011101110110;
#1 $display("%b", po);
# 1  pi=207'b110001000010010100000101110110010111101000110011111001100001000110000001011000111010110110001010010110111001111110000000001000110001101010110111100011010011010100110100001100111011000111101010000111000101110;
#1 $display("%b", po);
# 1  pi=207'b110001100010110000101100100011111101001010010001110001110101100111000011010100111111111101000100100100000111111001111110100110100011100101011110001101110100010010101011001111101011100110110101011010011010010;
#1 $display("%b", po);
# 1  pi=207'b001101101110011001010111101110100010010001111101101101110100110100101111110000100001101001111101001000110011000101001111100110001111010010101000001101110100110101110001111001101101011011000101100101100111110;
#1 $display("%b", po);
# 1  pi=207'b101110000100010110110101011011101010101000010100111011001111111010000000111110100110010101101001101110000101110110111000101001000110011101001111111010011100111011110111001101111000100001100111010100100100101;
#1 $display("%b", po);
# 1  pi=207'b000100110101100110010111100011001000111110001010101110001000111011011001001100010000110100010100110001100010110010111111110000110110001101100101101101001011010001001010001111001011010010010011100111010110110;
#1 $display("%b", po);
# 1  pi=207'b101001101000011110110001110111000100111101111110100000111001010010000011111100000101111110000010011000000111110110010111111001111110111101010011010010100011101110101000011110011110010101101010000111111010011;
#1 $display("%b", po);
# 1  pi=207'b001100011110111110011100011000111100011101100000110111111100100100111001101101100010001001111000110110100011100100010000010110111000110001001010011111010000100101100001111111010001111111010001011110001011001;
#1 $display("%b", po);
# 1  pi=207'b000101011010001001001111100010011010101101011111010100110001100100011100100100111000110010011000110001000111001110111011011111010110100011100001010100011110101010000000111110101111100111000111111101111011011;
#1 $display("%b", po);
# 1  pi=207'b101011100011101001010100100111011110110101010100000100010001001100000111110001011110100100101111011111001011010101010100011111110101110001111001011110111000001111110100010100101110001101011101101100100111011;
#1 $display("%b", po);
# 1  pi=207'b011000000100010101001011001010100010100001101000101111001000011000110001111010101011100001101110000111110011010000100011011100000110010001010000101101110110011010100111100100010110100011111010011001000010001;
#1 $display("%b", po);
# 1  pi=207'b001111110011101100001110100011001001100001011011110010100100011010111010011110010101011111001101000001010111000101011101101001101000000010000101100111011100010101100001110100111000110011000001111111011110001;
#1 $display("%b", po);
# 1  pi=207'b101011010000100010010110101100111010011100011111100110010100001000110101010001010111100011111100010010011000111110111110001000000011010010111100100110001100110001100001111100011010110101000001000011001000000;
#1 $display("%b", po);
# 1  pi=207'b010010101100110010111110111001010100001001100000011000010100001001001111110101111010101100111010101011001111000101001011011001111010101010001001010111101110000000111011001111100011001101110000111111110001000;
#1 $display("%b", po);
# 1  pi=207'b100101100001111000001101010000100010110011010101001100010011001111101010101101010110100101100000010110011001001110110011011111101011111101011110110000001001011101111010101000000010111100100011100011101110110;
#1 $display("%b", po);
# 1  pi=207'b100101101010111000100000011101000110011011011110101101101100100010101011111010100011001011001000101101011111100011011100101101011000100101000101110110010000110010100111001111110011110101011101111010011110011;
#1 $display("%b", po);
# 1  pi=207'b011010001010100100000000111010001100110001011011001100110011111100001100010100010000011010100011111111101011010110111101100110011011101101111101000010001011111110111000101101001001100010000101111110001100001;
#1 $display("%b", po);
# 1  pi=207'b011110000100100000100100010101001011101101100010111110011101010101001000001111111001001100101010100101110110100011100011011010010010010000100100111011100010001011111010000011000000110110011110010101101011111;
#1 $display("%b", po);
# 1  pi=207'b111101011111011010000011011110111010010110000100111100100111111011101111110011011111110101001000010101110001001111111100111110100101111101100011101001100101110010110001000001111101100110011001100111010110000;
#1 $display("%b", po);
# 1  pi=207'b101101000010000011001110000001110111100111100010010011011000000010001010010010100111001111001101101011110111101111001001110101010011000011101001100110101101111101011100000001100101000000111001001111100101100;
#1 $display("%b", po);
# 1  pi=207'b011011110101000110010110110001000110110010001111001110001000100000000111001010100101101100000110100101001110111010101001110011001111110010010000100010010001111100100101001100001110000101111001101111110001000;
#1 $display("%b", po);
# 1  pi=207'b111100011111111011100011110100100110100000110000001011101000001110111011010000100010100010110000000111000111000000111100111110110100110001110001010110110111010010100101111011001111000100011111001100110100010;
#1 $display("%b", po);
# 1  pi=207'b101010111010010101100000001000111001000000110011001011100110001001101000100110101100000010111100110000111111111101011000000011100000111110101011101000000110111001011010010100101100111111011010000100100111010;
#1 $display("%b", po);
# 1  pi=207'b001011101011010111100010010000111000010101010000110011011100101101011000100101100011100011010001010101101100011001100011110110000001111000110111000001001001011110101000010011001010101110100010000110100100011;
#1 $display("%b", po);
# 1  pi=207'b000010110011001110110011010001000000101100110011011101101010101101101010011100101001010111011001101001000011001011100011011000100100101010101001001010110010111001100100011000011011101100000000111011001111110;
#1 $display("%b", po);
# 1  pi=207'b011011101001101000101011010110001001010000000010110011010111011100011101010000111010011010001011010101110101100001111110110011110010011001010100110101110011000010001011111010011010001011111001101101010100100;
#1 $display("%b", po);
# 1  pi=207'b100001001111011001110011000101110110110010010000111010010111111001101111001111101010010111100101011010100001101011110001000100000000011100110001010110001100011010010010000000001011101001000001111101101101111;
#1 $display("%b", po);
# 1  pi=207'b011001111110110100011011010011110011100111110011111101000010111010000100101001100101100010100011000011000101110100100000001110001010101011001110100010000111010100111010111100011101011010101110100100110001101;
#1 $display("%b", po);
# 1  pi=207'b001100010010101010000101000011110111101100011100100100110110111011001110101110001100001100011111100000000100101100100101001011111111110011111000000101100101001001111110011110111100000000111111101111010000010;
#1 $display("%b", po);
# 1  pi=207'b010000111101001011110001000010001111111101010000000010001100011010001011011001110011111100111111101011011011011100011100100101111011110110101110100011100011101100000110001110100011101100101011101100000110010;
#1 $display("%b", po);
# 1  pi=207'b001000101101110111000111101001111100101101001011011111010011000110001110011011101111110100011000101000110000110001001100111000000100100011111011100011000000001001100100000001110001100001011110110010111000000;
#1 $display("%b", po);
# 1  pi=207'b001011111100001011110111000111101111010110001101110100110000111111111001000010011000010001110001101100000100101100110111001101010011001000101010001010010000000001110111000111110100000110111100010110000001011;
#1 $display("%b", po);
# 1  pi=207'b010001001110100000010110010010100001000000101000011100101101011100100000011101010010000000101110001001000100001111001111010001101101000101010100110111110010001001100000111000100001000101111011100110101101101;
#1 $display("%b", po);
# 1  pi=207'b100001000001000010111101010111000010011010101001010111100011000110010101111000111100000001101111100010001111111101011111011101101001001000110110001101101000110010111101000101101010001011001001101001001110001;
#1 $display("%b", po);
# 1  pi=207'b111111111000111111110110100001011101111011011111001010010011101100011011000101101001011101111010111110100111001111101110011110101110100111101000100100001001001001100011010000000110000110101101100101101000000;
#1 $display("%b", po);
# 1  pi=207'b100100010010001000101000001110000100010100000001101010100100110100100010000011001011100001001000010111011011100111011001110001101010101111111110110111001101111001110110000101001100010111100111010111110011100;
#1 $display("%b", po);
# 1  pi=207'b110000010010001001111110000011100011011010110001110110001101011011111000001011110110110111110111110010000110110010011101100111110111110110000100100101110001011001000011100001100000001111001000101110101110001;
#1 $display("%b", po);
# 1  pi=207'b111110110110010010001001110001101010100101110011000000100101000011011110100110000111100111010100010101100010100010001111001000010110010010100100101000011010110010111000101010000000111100001000110011110110110;
#1 $display("%b", po);
# 1  pi=207'b110110101001100000001111001111110101101010101000101110001101011000001000011000111000001101110000101100010010000000001001110011011010100101111001111011111011000110100010000100101010011111110111010100000110000;
#1 $display("%b", po);
# 1  pi=207'b011110101111101011001100001111110011011000111111110101100010001110000100111001110000100010011111101111010000100010101001000011011111000000001110010101000111010000111110000100001110000101010111101010001110110;
#1 $display("%b", po);
# 1  pi=207'b111011111111001011000000010001010110100010010111111100100100010000111101011101101011011001000101011010000000111100111010100000001100100011000111001101101101110110110111010100101000111100111110000010100110001;
#1 $display("%b", po);
# 1  pi=207'b111011100101010110000010001010010100110011100010001011001000000101001001101011011000001010011110101000001011001011100000101101110010110110100100011111001111010111001111100111110011100111110000011000110000001;
#1 $display("%b", po);
# 1  pi=207'b000010100111001011101011010111001100110111010100011101111001010100011111110110111111010101100111010010100110100011011001010011010010001010011010110101010011110100101000110100000000100000000010011011000001111;
#1 $display("%b", po);
# 1  pi=207'b110110100110111011101011111110000001010101001000100001110000100110011011011100001011111010100010111110010111100011100100001011100110110110010000111110011101111110100110111001010010100111111100100101111010101;
#1 $display("%b", po);
# 1  pi=207'b010010101001101101100001010110000010100100101110001110100101110101110000000001111110101001111101100110010111100000001100111100010001100010011000110110111110011000011100101010101100001101101101111010101101001;
#1 $display("%b", po);
# 1  pi=207'b101011000001110101001010100110100000010011101010000100101111010010111001100000001010001001101000001110001011100101110010101011110101000111110001001000101001000101101111001111001011101010011011010100001111101;
#1 $display("%b", po);
# 1  pi=207'b011101001000000000001010101111001101110111000100110110100111101011101101111011100100011100011100001010101101100011011000011011001000010011001001000110000001010101100100100110111110010101001001001010111100011;
#1 $display("%b", po);
# 1  pi=207'b000010000000110111011111001100010001000100001111011100000000001000001111100001100001000111111001111001101011101110010101100111110010100000100001101010001100100001010000110111111001100101011110111001011110011;
#1 $display("%b", po);
# 1  pi=207'b010100000011001110111001001011101011111101101010110011101110111001000001100011101101111100011011001001011001100001110001010001001011110100001001010110000111111100010011010011011101111001110101011110011101000;
#1 $display("%b", po);
# 1  pi=207'b011101001100011001010111001010101011011101110101100100011110111111011101101101100101100101101000101010010001011000100111000010001000011001111101100001111001111111001100110101001010010011011110001101010101110;
#1 $display("%b", po);
# 1  pi=207'b001110110110111011110111000100111001110010010011001100101010001001111001111101010010011110011111001010001000000111001100100000100111011101000100110110011011101001110001000100010110011001010111100011001011100;
#1 $display("%b", po);
# 1  pi=207'b100000110010010000011101011111000010110000010001110000011001111111010001101101000010010100101011100100111000101001000100101101000001011110100110110100001000010101000100110111110001011101010001110010110110000;
#1 $display("%b", po);
# 1  pi=207'b111000110100010000111100111000001101100100110011100110000000010110111011110101011001101101011101100000110101101000001010101111000010010101100100100001000100000111101011110110111101100111100000010000110000111;
#1 $display("%b", po);
# 1  pi=207'b110011100000000101010111111011001001111100010100110101110010011011101110110101001110011010100000010001111010000001000011111110101001100110110110100000110110100110000001010001011011001011000010110000000110001;
#1 $display("%b", po);
# 1  pi=207'b001110001010010010100111001101010001000111111110101110101001100100000101000110010110111000010110110010100000100001111001110001011001101010011000100101000100001011000010101100111111110110110010110111101001111;
#1 $display("%b", po);
# 1  pi=207'b000011100100011110000000001001111010100110111110011101000010000101110011111110101110011010011011011010011100010110101011000010110010111001100100100001101100001000001010001011010000100011110101100001000001110;
#1 $display("%b", po);
# 1  pi=207'b101100111101111011101001001000011001110000000100100110100001101001111001010101100011001011011000010001101000011010010110010100010010010110111100100000101100010000000000011101101100010110110011000001111000000;
#1 $display("%b", po);
# 1  pi=207'b011011111011101000101111101100010011100111011010011111101110101111010001101011010010011100000001011011110111000100100000001100100101100101110111010111101101101010100011000111000100101111110011111101101001001;
#1 $display("%b", po);
# 1  pi=207'b001111010000000110010011011100010001011110011101110010110001001001101001111110110100001011010001101110101100000010100111110101011101101001001011101111000001011001001011111101110010111111101110000011010000011;
#1 $display("%b", po);
# 1  pi=207'b111110101011111110100010001111101001000110000001011110001100100111011100011101110010101011110001001010101111001010100110001010111011100100011001101100000101100011001100001101010110100111100000100001110001101;
#1 $display("%b", po);
# 1  pi=207'b101110111000100011000011001000100111000100000111010101010111011101010100001101100000000011001011000010001010111100000001111010010000001011100111011001010000001111110001010100011000010011000000000010000101110;
#1 $display("%b", po);
# 1  pi=207'b000110101000001001001110100010100100010101011011100110111101011110100011010100000111000000110100010010111110010011001100001010011110000010010111010101111011111110010000001001011111101000100000100101010101111;
#1 $display("%b", po);
# 1  pi=207'b101100111101010001101100011000000100101100000111000001110100010000110010111010011000111000001000111101001111000001010000000000010000011000101000101100011110110101010001111010010011010110101011100100101110000;
#1 $display("%b", po);
# 1  pi=207'b010110110101010110010110110001000000001100011011000001110010011000111111001010000011100110000100010001110100011110010001100111000111001111110111010011110100101011010111010001010101001101000000000000001001000;
#1 $display("%b", po);
# 1  pi=207'b001010110111101110011011001010100110010010000001001011001100101011011011011001110000011000001011101100011111110010110101101010010000110100010010001111111001100111000001000010101011111010000101000010000001110;
#1 $display("%b", po);
# 1  pi=207'b001010000101001010100100111111010101010100101100100101001000110001110111101100100101011101010010100101000100010001010111110111000111011101100011111010010101110111011111010110001011011001100011001111011111000;
#1 $display("%b", po);
# 1  pi=207'b011111111100000101101001000111011101101101111010101010100111100011100110110001011110000010010010001100001000100111000100000010100101110011010111010010001011110010010100111001011011000100101000010111011111011;
#1 $display("%b", po);
# 1  pi=207'b001000110101110000010010001110000111011100100001011111000011011100001010001001000100101101001111001011110101011111101010110010011000101010100011100011111010001111100110100010111100110110101001010000101110101;
#1 $display("%b", po);
# 1  pi=207'b010011000111110011111111000010100111001000001100100001111010100100011101011010000111110001001000010100010001110101000110010010100001000111000100000101111111111100111000010001001101110110110000100110010100110;
#1 $display("%b", po);
# 1  pi=207'b100010111111001010010100000011111000100101000101110000110010011010111101000000010000010000110001011010100000110110111010000111011010000010101010000100001100111100000100111100000101011001011110011011011101011;
#1 $display("%b", po);
# 1  pi=207'b000000010011010101101010000000100001110011010100001000110001101001000100010000010100001110101110101000100001011111001101110111001100010100010111101000101011110101011101001000101011010011011100000001010100110;
#1 $display("%b", po);
# 1  pi=207'b100011110110101011111101110000011101011010011100000010101000010101011000101100010100101001010111000110110000110011101110110100100001111101010111111000011000100110010111100011011000000111001001110001111111101;
#1 $display("%b", po);
# 1  pi=207'b011011001110001011110000111010111001001000101000101010101101010110010010100110100111010110001001001100111000000010011110011111010000000110010000001100011111001011100010101111110010111000100111100010000011111;
#1 $display("%b", po);
# 1  pi=207'b001010111111101010100001001100010000001110101000110011101001010100001111100100001111100100101011010010111110100101100100111110101110100101110101100110111001011011111011100100011001001000011001001111111111011;
#1 $display("%b", po);
# 1  pi=207'b110110001011010010001100101101110001001011000001100111001010111000100101100111011110001101000100011100101110001010111111111001000000001111010000011110101000100011101011101100100110001101000010010011110011001;
#1 $display("%b", po);
# 1  pi=207'b101001010111000111100010111101010100001000000100001010111111010111101100101010110010010001110101010011011011111010011000110001111101100000000000110110011100001100100100111110110100111111000001000101110011010;
#1 $display("%b", po);
# 1  pi=207'b101111001111110011001011100000000110001001010100000110111110000001110100010000010011100001011111010011010000001100000010101010011101010111111010110010100011101100111101111010111001001100111101111001000100011;
#1 $display("%b", po);
# 1  pi=207'b010010111110010100011101111101100101111010111011101100011101000000111000100010110001100101011001100001000100001110101001000110110110011011000101101011111110100101000101001101011010000110010110111010011000011;
#1 $display("%b", po);
# 1  pi=207'b001000011110100001000001101011100111011000111000011010000111010010010001011100001001000000001000111110000001011011001111101100011111110110110011110000111001010001000000110011010011101001001101111111000101101;
#1 $display("%b", po);
# 1  pi=207'b101111001101110000100001011000111110000100111111000101101001100110111010110111001001101000100110100110101000011100011111100001011110101011101110110000011011010100001101011000100011100100000001010111000011111;
#1 $display("%b", po);
# 1  pi=207'b111000101001111010101101000111000101111110110010110101011110100101101100110011001101101001110101110001011010010000000010001110010010011101001101101101010111100011011001110110001100011110000101101011011000000;
#1 $display("%b", po);
# 1  pi=207'b111100110110100010000111100001001110100011000100001000111101011011000000001110000011111111100100110100010111011111011101011000110100100101000000110001001111011101101111011100010010100011101010010111100001000;
#1 $display("%b", po);
# 1  pi=207'b011010001101001101110111101000001000001010111101011111010001100110000101101111110101011111111110010110110101101011100010010100011001000010101100001101010011000111010101111001011011110111001101000010010011010;
#1 $display("%b", po);
# 1  pi=207'b101101111101001110111010000110011110000111111001111001111011100011100000100010000101011111111100111001001100010100111001100010001000000001110001000101101110001010100001110011100111111011011010001111000010000;
#1 $display("%b", po);
# 1  pi=207'b000000100100000111110001100001011101110001110010000000010001101000011110001101100001111011100111001101011001101100010110111111011111001010000011100101011110011011010011111010100110010100100110001001000101111;
#1 $display("%b", po);
# 1  pi=207'b111001010111110110111110111001010101011001011100011101101111110100010111010011100000011010001111011011111000100011111111111101111111100001100111001101000001100100111101111110101101100001111011101010000000011;
#1 $display("%b", po);
# 1  pi=207'b011000000011001101010001000001010010110110110101000101100100111111000010110011111100010100101110101011100101101111101010011011001000011111100001111010110101010010110001110111010001111101100111010010011100101;
#1 $display("%b", po);
# 1  pi=207'b010010001011100101101110010001000100110000111101001111000111001110100101011011110000100011100011100100101110000111000011101101100111011010111011010010000001010000100110010110001011110000100100111011110100001;
#1 $display("%b", po);
# 1  pi=207'b110001011100001011100100110011101001011111011110001101011100101000110010101000001000110100111000001011100111101111011110110001001110011000000101011010111001000100011011111000011011001000000101001001011001010;
#1 $display("%b", po);
# 1  pi=207'b111111100000110111000111010011101011100110110001001100011111100110010100000000100001000001011001000111000101010111101011010010100001101001001110011011001001111100110111011010010100101110011111011101111101010;
#1 $display("%b", po);
# 1  pi=207'b011001011101111010110010111101101110000111010011110000011100010110111100100000011110111001011000110011011010001111011001101111110011010001010111110001001010010001001011110000110110011111010000111101011111111;
#1 $display("%b", po);
# 1  pi=207'b010011011100110010011100011010010011101111000001110010111100001011001100110101001000010010001101011000111100110100100111111110001011000110101010110100100000011110001111000010001110110000000011110110111011111;
#1 $display("%b", po);
# 1  pi=207'b110100000000110100100011000011110100110100010000001110000001000000100011010010100011110010010110110011101011110101111001001001111010101111010111001010100000110001101101001101110011000000000100110100001001101;
#1 $display("%b", po);
# 1  pi=207'b101110001110010101010111011011001110000101110100110001111001001001010000011101011000000011111100111111010101001001110000101110000110010010011110100100100001111110100011111111010110111010010010000110110100001;
#1 $display("%b", po);
# 1  pi=207'b010001100111010011111010000100001011010000101111010111001100100101011111010101110110111010010000111110010111001000000100101001100101001011000100001000011110111001111010001110000011001101010000101000011110000;
#1 $display("%b", po);
# 1  pi=207'b110011101110110010111010001011010000000101001001011110011111101100111000010100100011110110110011001101010000111100100101100000011101011000101000100111010110100110100110001100111000001101101111100001111100010;
#1 $display("%b", po);
# 1  pi=207'b011011011101000101010000000111100111010001111000100000010110111000111011010101101100011111111000000011000000001010111011111110101101010000111000011100001010101100001011001011110110001001100101101101010000001;
#1 $display("%b", po);
# 1  pi=207'b100100000100100010111100100111110111011000111001011001100010010010111101100100101100001011111010001010001000011001111110000100101101001110001100101101000001100010011001101101011111010001001000101011100000010;
#1 $display("%b", po);
# 1  pi=207'b011111011101111101010101001010100011010111000011101101010110101110101101101100100111011010111010011101111000000000010001111011101001110010010100011111101110010110110011100010110001101111000110000110000100101;
#1 $display("%b", po);
# 1  pi=207'b000110111001100010110111110010101010100001101001001010110101011001001100111001011100010110101001001000100101001001101011100010000110010111011101000001110001011101100010111010001010001000101010101111011001001;
#1 $display("%b", po);
# 1  pi=207'b010100011010000101000001011111111001000000000000111000000110100110111010001100011011001010010001100010010111111011011010001000011100101011010010000111010011000000000100010100001000100000000001100000001010000;
#1 $display("%b", po);
# 1  pi=207'b010111111010110100101110011011011101100100000101111010100011000100111101110100010001010101010001000010111000111110001111001110001010111011101000100010101111101100000100000001001011001110101111011011011110001;
#1 $display("%b", po);
# 1  pi=207'b111010101110011111100000000001011010011000111001010011011001100110001001101111011011010010010001010001010101111111111010101010000011001100010000011000011011100010000010100101100001011110110010000111100000100;
#1 $display("%b", po);
# 1  pi=207'b110010010101001010110000101101100101000100000110111100000101000011010100100001111100101011100000010101111111010111110001111001101100011000001110101101101101001111110010100011001111110101100010000111010111010;
#1 $display("%b", po);
# 1  pi=207'b100011110110111000001110111010110111010000000010101111001110001010110111101000000000011011010001110010000000101010010101111100110111010010001011110001100000111101001100010110110011101010111010111110011100000;
#1 $display("%b", po);
# 1  pi=207'b100001000011011101111110111000000111011101100001101010010100101001110000001011011011010110100110010011001100110110000111101101100110011101000000010110101001100011001110111001100000100001011000110101100101101;
#1 $display("%b", po);
# 1  pi=207'b110101011001100001101011110010101011000000100111010000000100110000110001001001010011111010110100011000000111001011111111000000111010110001110011000111000111101111110010110011001100101100110101000000111110100;
#1 $display("%b", po);
# 1  pi=207'b111011010111111101110011001100101011101001101011101110000100110010001000100101110001111100000100110111010101111100101010010000010110100010000011011100111001100000100010101010011011100011111000110100100000110;
#1 $display("%b", po);
# 1  pi=207'b000110011111001000110001111010100000000001101110000111111010101001101100111111000000001110000001101010101110101110110011011001101111000000001010110101001001010000001001000110001101000111000101001010011011100;
#1 $display("%b", po);
# 1  pi=207'b100111011110001011110101010010011100111011100010101001000010100000010001011000000100101010110111001110100001100100100111100111101011010101111111100101000101010110010011010100100101010010000101010111111100000;
#1 $display("%b", po);
# 1  pi=207'b011100010111111001111011010100001010110101000100101000000100110111110010000100010111001000101010110011111101101100011011110001101010010101100101100101001010011011000001001100001010111111000011101111100011110;
#1 $display("%b", po);
# 1  pi=207'b111010011110100000010100011001011011000000111010111100111111010010111101001011100010101110110011010100111111101100110010101001011101111010011110011000000100001001101000010011111101010101000101111100001101111;
#1 $display("%b", po);
# 1  pi=207'b000000101101100010101110101000100101111010101110010100100011110110111111110110011001101110011011001000000010100100001000011100011110111011001011101011110010001110110100111100100000101011000100100010101110110;
#1 $display("%b", po);
# 1  pi=207'b001101100011111001000110111000110010011000100101110000101000000001101110101100110101111001111011010101001100011110001001010110001110100101101001001101001001011001010000001100101100100010111100100111001110100;
#1 $display("%b", po);
# 1  pi=207'b101010100100011010111111100111111000110111111000111001010011001001010101010000000101011011100111101111000001001110001010110000110001110011011101101110100011110101101111110100001011111110000110111110000111111;
#1 $display("%b", po);
# 1  pi=207'b010010100011000000000010010001101011110100011111010111110101000001111011110011001100011011110010011100101110000011011111000010000111110011110100101101000111100101101001011011001111000001111000100110011011110;
#1 $display("%b", po);
# 1  pi=207'b011001101101101011101100101010100000100000001111000011100100000010111010011101111110001110000110101001001100001010001010001110000011111000100100001110110001010000001100110101110101110001010110011110100111001;
#1 $display("%b", po);
# 1  pi=207'b101000000010111000111101110111101001011001100001110010000110011111000010010100011111001110101111111011000101011011011001010100011110011111000101011110101100001001101110011011111111000101000001110101000110111;
#1 $display("%b", po);
# 1  pi=207'b101100101000011101100001110000011110101000110110110011110001110001011100010111101011100001011011111111011101001111000111110011010101010011010111000000110010101000111100100100001000010000100000100101001110001;
#1 $display("%b", po);
# 1  pi=207'b101101100100100100001111100001001000000111011110010100101011111000111101011000011001100110011111110011011110101111010000101110101011001010110111000111010000000111000101111110110010011011010011000101101001100;
#1 $display("%b", po);
# 1  pi=207'b101001001100011000010010011111111100100111011001011001011111101001100100000001011001011010110110001000011010100101101101000110000001000011101100011110000100111011101101011101000101010111110010011100001101110;
#1 $display("%b", po);
# 1  pi=207'b100100100101110010111110100011110100000111111011110110100101111111000010011000000011110001001110010100100011111000011110010100001001101111011100100001100101000011110010000000110001000110010010010111111010100;
#1 $display("%b", po);
# 1  pi=207'b001100001000000000000001001001000000111000001110010100000111111011100001001111101111100110010110110111011011110001000111101010010110110111100110100011010110101111011111001100101000001000110010010100010111100;
#1 $display("%b", po);
# 1  pi=207'b111010010100011001100101000110001000010111101100000100110000111111100001001110011110011111110001111110001010011111010111011101001111111011100101111010001010111001001100100110100101101111101100000101111111000;
#1 $display("%b", po);
# 1  pi=207'b001010111000110110000000011000110110010001000100110110110001000010100110000100100010100011010101011100100100010111101000001110010100110011001100111011101000000100101110101010101110101000101101010100111100110;
#1 $display("%b", po);
# 1  pi=207'b100011010001111101001011010101110100100000101111011011100100000011110110111010001000011000100101100001001011000011001000001010011110011011100011101010000000001100001010101111010000010011110100111101100100110;
#1 $display("%b", po);
# 1  pi=207'b100101010110000010011010110010010100111110001100011101011111100101011011011000010001110010011110000110101100111010000000011001100100110001010101011001101010000111110001000100000101000001011000110011011011011;
#1 $display("%b", po);
# 1  pi=207'b100111100110101010010101011111011011001011000010011110010010110010110110001001111011110100111000001101010101001010111100110000110111000111101000011010110110001001110000001000001001000110001110101010111011100;
#1 $display("%b", po);
# 1  pi=207'b010100111011000111111111010100101010011101010000110000000101001000100111110100011111101000010100111110111111001110101011110100000110110100001111000001000001010011100111100010011111110100011100011001101101101;
#1 $display("%b", po);
# 1  pi=207'b001011111000001011000001100111101000110000011100011111101011000011000000010100110110001110011000110010110011111010110011001011110110100011101010111011011000101000001110011011010010101000110111110011110000101;
#1 $display("%b", po);
# 1  pi=207'b000001000011000011011100101001111110110011000101100000011100110000011010000001101010011001000010101011010000110101001111111000110110011000000000011101000000011101101111010100110110010000011000110010010010001;
#1 $display("%b", po);
# 1  pi=207'b111100000100001111011010001110010100100010010101110110101101010100000011110110111001000011100111001101111011101001111000110100101110001100100111100100101101000010001111110011011101010011011100101110000010100;
#1 $display("%b", po);
# 1  pi=207'b110110110000110000100001000010001111001001000101101011100111110100000100011010101000010100110010001011010010111101101101000110111010101110000111101100100110111110111110010010001110001110000110011010111001001;
#1 $display("%b", po);
# 1  pi=207'b000000000110011101011101001100110101011100110110011100110000010001100100011101100101010000111000101110100010101010100001111111101111110010110100110011111100101111010101011111101111010101111011111001010011010;
#1 $display("%b", po);
# 1  pi=207'b011111111001101111001100110100000111110110100101011001010001100001001001110000010010000110001110001111110001011101111000011100100011001001001101101011011111110111111001110101010101011001101010010111110110110;
#1 $display("%b", po);
# 1  pi=207'b100011110110000100100000111110100100110101010111001001010001101110101101011101101110011101001100001001111011010011011001001001001101001111001111101011001010000001011100011001101101010111000101000000001011110;
#1 $display("%b", po);
# 1  pi=207'b110010010000011000000110001010001001011110110011000010110000001101010000010000110111011011101011001001001000101011111011111001111110110111000010011111111010111110101100001101010101111010111010111011101010000;
#1 $display("%b", po);
# 1  pi=207'b101001011000110011011111111000100111000111110111000000011110001101001001110001100001100000101101111101001000100010101111000001001000011000001110011110010101001111100001110111010101011110110110010011001101011;
#1 $display("%b", po);
# 1  pi=207'b011100010100110100011101010100100100001101000110110100010011001011001100000101100101101001000111100001000010111110111110111011011011010001001000100000111001011100001110111010011001011010001101110110011011011;
#1 $display("%b", po);
# 1  pi=207'b111110100000000010110000010010101101011001111001001110001011110001000001011001000100100111001010000111001011011110110001000111100111010111111100100101001000010110101100001111001111110011111101000101010111111;
#1 $display("%b", po);
# 1  pi=207'b010011110100001101100000100000000101111000101111111001100111011101111001000100100101110010100000010101001111011011010111011100001101111001101010001010000100001101011101000000110100010010010110001011000000101;
#1 $display("%b", po);
# 1  pi=207'b100010110001000010000001000100011100101010110101000001100000100101010111110111011001101001100000000110000110001101100110110001111010011001000001101110001101010001000100011110011000101000011110000001100110101;
#1 $display("%b", po);
# 1  pi=207'b011011100010110001010010000101111011010110100000010011010111011111000010010000001001101011110100110001000101011101100001101001101011110111011111011101101000000100101101001011111011000010010110100001111101010;
#1 $display("%b", po);
# 1  pi=207'b110111110011110110101101110001111011101001010000111110100110011010101111110001101000100000000111100111001110010010000001101100011111001101011011010101110111010011111001100101110000011001011100110111110111011;
#1 $display("%b", po);
# 1  pi=207'b101010100111011111011000010011110000010011110000101011010001001111000101000010000100000001011101011111000101011110000011101111010011000111001111001110100000110001111101010001001110000010110101111110001001101;
#1 $display("%b", po);
# 1  pi=207'b100110011010100010001010001011111111100110010101101101001000111010101000101111100111010011110101001001111111010111111100100101000011110001000001011101110101010010100111001011001001101110110001011110100010101;
#1 $display("%b", po);
# 1  pi=207'b111101011101110111110100111100001011100011001110001010010110001110110011110000001011111000111010111000010000101000111110101000000010001111110010111000101000101010000001001010111101001000010101110011110001101;
#1 $display("%b", po);
# 1  pi=207'b001101000101110011010010111000111111010101001000011000011011101100110101110001110100110001010001101001100110000111101100100101001010010110001001011100000001000010110010001001000111101000111111100100101100010;
#1 $display("%b", po);
# 1  pi=207'b000100010101000100100110110001101000111010111010001001101010111000001111101001011011010010000110111001001101010110011101010001111111011101010001010111000110001001111100000010101101111100111101111100100100111;
#1 $display("%b", po);
# 1  pi=207'b100011000010111111000000010010111101001100000100111110101001101111101110001010000101011111110010010110011010000011111100110001111110101010001001011101000001011001010011100000100011011010111110001000111101001;
#1 $display("%b", po);
# 1  pi=207'b010011110110011010110101100110111101111011001101101001011111101011001001100111010111101111000001100100111110011101000111101000000000101101101100010010100110110000110010101110001000111100111000010011111011100;
#1 $display("%b", po);
# 1  pi=207'b001111000001010101000101000011110010110000101000111111011110101001111110001110001000000001110000101111001101001001011100111101110011011110000111110010111010100111011011110001001110100010110011011101110100010;
#1 $display("%b", po);
# 1  pi=207'b111010000011010111111111101100000100000110101110100010110011001001111001101100010111010000110111001001101011000110011011110101111011100010001011000100100111100011110010100010111011000000010110110100000010011;
#1 $display("%b", po);
# 1  pi=207'b100000010110110001001001111101101010010010000100111100110000111100111011010100101011001100101001110001000010001011100110010000110101100101011000001010010010110010011001010010000100100101101010101010001111011;
#1 $display("%b", po);
# 1  pi=207'b111010011010110110101001100100100010000000111100001111000010001111101100110110000010001101100000101101010110110000010110110100001101111011000010110110110111011100011001110111010101111111110111110001110101010;
#1 $display("%b", po);
# 1  pi=207'b001011000110101011010000101001010110101011000000101000000001111101101111110001111111101001010100010010000010010001010111000100111100010110001000011110011011111011000011111110111000010111101111011111001011101;
#1 $display("%b", po);
# 1  pi=207'b000110010100001010001011011011101001110110011001111110011110000101111001001000010010011110100001101111110111110001111100011001010000110100011010000001101010101100001111010100001010100000101011101101011111101;
#1 $display("%b", po);
# 1  pi=207'b111001010000011111100101010101100001101000011000110101010100011101001100001011111111000110011111011110011001111111000001010110100101100000100101011111011111110111011101010111110110100001100110010010011010100;
#1 $display("%b", po);
# 1  pi=207'b110100100000101011100011111001110011110001011110010000100001111001011010000101110000110010001110100100010110101111010101010010001110101100111000110011011010001100000101110100000100111001111111011001110001101;
#1 $display("%b", po);
# 1  pi=207'b100110010011100111010101111000010111011110011000000011000001101001101000011101110100111011100111111011010101110110101101001100000010100110110010110111111101100001100110011111111001111110011011101101011100111;
#1 $display("%b", po);
# 1  pi=207'b110001100101100010110011100110000011110000000001110010111000101100011100101000001000110001101101001001001111001100000010010111001110010010101000010010001011001011111010111000001101110100010110110001111011100;
#1 $display("%b", po);
# 1  pi=207'b101011110001000001011101111100111010101111110110011111101001001000111110101011100101011011011110001101110000101101101011111100100001111110011000100011000110100101100110001001000010010001011101011101100010101;
#1 $display("%b", po);
# 1  pi=207'b010011111101110000010011011110011011010011110110100101110111100001111100001111110101100011101010101010001000111111101001011010000010101011110110000111100111100010001101010111100110111111110100010100000010011;
#1 $display("%b", po);
# 1  pi=207'b010000011101111110001110001101010111101010111001111001101110111110000010101000111010111001001010111100110010110000010100000101110010001000100101110110010000000100010110110111001110111010101011010100101000110;
#1 $display("%b", po);
# 1  pi=207'b111100100010101011011010110010011101100101110111000010110101100110100100101000100010000110111000001000011000100010101001101101110110111100100100001111010000000111100110000111110011000011000000001111000110111;
#1 $display("%b", po);
# 1  pi=207'b011100111101001010100110100001011001001110100011010100111110010111111100110001111011010010000110011111111001101001110101111010011010011110000000010010110001000111011101101100110101011011110011001110101101110;
#1 $display("%b", po);
# 1  pi=207'b110000000101101100101010111010111001011011001111111111100000111010010111000000101110100000000101000011110000111110111100010110101010001110111001000100101000000111011110001011010111011100000110001111101001001;
#1 $display("%b", po);
# 1  pi=207'b011100010101111101001011101010101001110010010001111011011000011110001111011011111010000111110101001111111011000101011001101010100111001100100001110111101101111011110100101110101100010111111100101000110100001;
#1 $display("%b", po);
# 1  pi=207'b111100100000100101000100000010101001010011111001101011110011101010111000011100001001001011011001011000110110100110110011110100010111010010111011011101011111001010000011000000000111111011000000100000010011111;
#1 $display("%b", po);
# 1  pi=207'b000111010100011000100001101010100011001100000110000001101011110001111001110100010000111111001111010101100100100000011111111011110110110110010000101110101011101001000110000100100101001000011101001001110011110;
#1 $display("%b", po);
# 1  pi=207'b100100001101010110010101100101111110000001011100000010101100101110100110011010110100101111110000110011101101010100100000111000101000010111100010010101010001110010111110001010111101011001111100001111101100100;
#1 $display("%b", po);
# 1  pi=207'b101110111111110100111101001110110110111110011111001010001001110000100011001100001010101010101101000000100111000001001011011001010001010000010010001010001101010001011000011001010010011010101001100111110010011;
#1 $display("%b", po);
# 1  pi=207'b011111001111000110011101010010010000001100110110111110101011001011011111110000100110101111111110110110100111100010101111000010100110100000101101101110110001000100011010111011101111100111001101101100011010011;
#1 $display("%b", po);
# 1  pi=207'b000001000011110000100001001111000010101110011111001000110110000010010011100000100101001111101000011110111111110101011010100001011101110111011111100001101111000001100011101011110101001111001000011010010111000;
#1 $display("%b", po);
# 1  pi=207'b000110111100110001111110101010011011100011001000001111001110001010010100111000110101101101000101101001000110100011101000010001100100000100010100100010101001000001011000000110110111000000001100110111110001000;
#1 $display("%b", po);
# 1  pi=207'b110010010111011100010110011100001111100011011100010101011001101010010101100000110100000011000111100100100010100101110101010100101011000101110101100101001110111111111011110010101100111010100111000110101000100;
#1 $display("%b", po);
# 1  pi=207'b101110001100100111001101100011100011101000110110010111011100001000001010001111100001100100001111001101100110001101101111100111010001010000000111011100100110101000001010011010111101100110001010001000100101001;
#1 $display("%b", po);
# 1  pi=207'b001101100001000000100110001010110011011111000110010111000011000101011000011010000010011101011101101010100110011011000011101000100000100111010110010001000000011100111100100011000000000000000000010111111011001;
#1 $display("%b", po);
# 1  pi=207'b101100010111011001100111010111000011010001011111111110010101001100100101111010100000010111000001000011100011110100111010110010011110100110011011110110000101000110100000110110011111011110100101010100010101001;
#1 $display("%b", po);
# 1  pi=207'b000000101111100000110101101111110110000000110111110111000010011110001111010010011100101111110101101111110000001110000110000000111001010111000110110100101001110110101010101101001001101101001100101011011011001;
#1 $display("%b", po);
# 1  pi=207'b110001010010011001010010010111110000010001000101000000001100011000111010001110100101100011000101101110110000001100001101101011100111111111001000011110110100110101110110000000000011000100110011101001110100111;
#1 $display("%b", po);
# 1  pi=207'b110110001111111011100000001011001011011101011100010011000101011111100111110100001000010011000111101011110000111000011100011010111001110001110101111000110101100111110000010011100011000011011111001011110010101;
#1 $display("%b", po);
# 1  pi=207'b101001001100100110111010101110111011011101100000010100011000010111111111100101001001100011110101001011101000101101100000100001011111100111000000001111001110011011110000101101010101001110111111101010111000110;
#1 $display("%b", po);
# 1  pi=207'b111110110101111001101111111000001001101100111011000110001111101000110001011101111000010000001010111110010010000100010111101011100010101010100110011011100001011111110101001110011011011111111011000100101011111;
#1 $display("%b", po);
# 1  pi=207'b111101001101101000110110111010001000111100001000111001000010010101011010101010110110001101111110101000111110101001110101000010000001110111010100000110110100011101100010001011100000000011101110111100100110001;
#1 $display("%b", po);
# 1  pi=207'b010100000010101101101010110000011010110011110101000011011100111010101010100000110001101001001101001001100001100111100111110101101000111110111110001110110110101010011001011000011110101101010000101010100110000;
#1 $display("%b", po);
# 1  pi=207'b100010001100101011110000001110011111010000100100000010101101000011010011001101000100101101100000111001110101011011100010010111010000110010100101011111000111011001011100001001000100010110010000101010000110011;
#1 $display("%b", po);
# 1  pi=207'b000001100000000010000010110100101101010001001000100100011111000101110011001001000001100100101111100010101101101100011000100011100001010000100110000000010111001010000101111000101101011001001001101101100101110;
#1 $display("%b", po);
# 1  pi=207'b001000011010000000100011010000100110101010010011001011101101011101110010010110001010110001101101011110101000101001010110011011110101111100000010010111000100001000101010101111111110010011011000000001001100011;
#1 $display("%b", po);
# 1  pi=207'b010010111111101110001100100101101011001000110011010101001010100100010010000111100001011000111111111000001111110000110111011100111000011101111110100110110111101010010101011000000100100111000010111100110111000;
#1 $display("%b", po);
# 1  pi=207'b111111110110000000111100010110000011110010110001111111011010000100011010011111110111001010111111001101000010000111110100000110011010001011111000111010001110011011001111111001100111010001111100001010110001110;
#1 $display("%b", po);
# 1  pi=207'b001111000010010000011011100001000010100010011111000011100101010101101100001100110001100000001011000000010000110100010101011001001011001010100110100000110101010101011100001111111011100110011001100111101000011;
#1 $display("%b", po);
# 1  pi=207'b101110111110010000111110000001000111110011001000100100110001110000111110010110100000111011000101101101011111000110000011110110100001000010001010101010011111110100100010110000001111011000000000110111001000100;
#1 $display("%b", po);
# 1  pi=207'b101111111100100111011010110011110000000001110000110110010110100101110111101100000100100100110001110101010111111111001001010111010011010000101111000111111110111111100100100100000101100101001100001011000000100;
#1 $display("%b", po);
# 1  pi=207'b000000111110000111000101001010111011110110110100001111011110110110101111101100101000100111001000111000101000010001110101001101110101011000010100111110101000000100011111111101110011011100111110101100100111000;
#1 $display("%b", po);
# 1  pi=207'b100110111011001111001000000010100000100101101110101101111110000010000101110101101100101010010010101100111000111101000100100111100000000011101100011000110000001100001001000011000001011010000011011001010001101;
#1 $display("%b", po);
# 1  pi=207'b111010100101001000001100010010011001110101100101101111001111100001000000000010001101010111110111000011101111010100001010101110001001110110111010110100111011011101101001110110011111110010110000000100101110010;
#1 $display("%b", po);
# 1  pi=207'b010100100101110010100110011111011101101011011001000001000110001011101001011101011001101000001001110000100010001010011111101000010010010010101100000101111100010111011100111001101001010001101010110111100111001;
#1 $display("%b", po);
# 1  pi=207'b011101111000011000111110001100010110000101100110111001101001000011111100110111010111100100100011110010100010010111011101101110110111011011001110001000110110011111011111000011111001110100110011000000100011101;
#1 $display("%b", po);
# 1  pi=207'b000110111011110100101001010000100111001101000111001101100001011101000011011100001100111011010001111011001110101000010000000010110000111001100011100111010000010101010001101010000011100110101010111110100110011;
#1 $display("%b", po);
# 1  pi=207'b011111111000010110111111101110100111100011111111000011011011011101100001100101101110111110000100010011110110001101011111011101110011100010101101011000001010000101110100100011011111011010101000101011011111001;
#1 $display("%b", po);
# 1  pi=207'b111100010110111110110111101000110001010010011011001000000110100111000111110010110100101010001010111000111000010011110010100001110010000111111100100011011010100110100001000101110111011000001001101010110100101;
#1 $display("%b", po);
# 1  pi=207'b101100010111110011011100011000110011010110010100001001111001011100100000001011100010101001000010000101110001011111010001011100011001000000011100000010001011000110100011010110100011010101100000110110000001001;
#1 $display("%b", po);
# 1  pi=207'b011001111011010101001010110001101111111111110100010101100011011111101100100100100001010101100011100000111001010100111111011100011010110111010011110111101010110010100011000011111101010100110100110101111110100;
#1 $display("%b", po);
# 1  pi=207'b000010100000001100110001011110010010011000010010111010010100100110011100010100100101000001101111010000010100011011001111000001011101010011000100011111001111010101101100110111111100010001001101010110110101110;
#1 $display("%b", po);
# 1  pi=207'b111011100110110111000100000101011101010010001001011100100110001111011001011000110100101111010000101111000100000001100001111100001000000101001011000111111010010000000100010111110010100001101011101101010100011;
#1 $display("%b", po);
# 1  pi=207'b000111111001000001000001001001011000111101111010111001101101110110011001100010001110110111001000101100010110111101100010000011100010100111101011110011011100001101110100000001101110100101001101110000010001100;
#1 $display("%b", po);
# 1  pi=207'b111101100010010011110000101010101110001011100000000101100001000100010100101111011001101101000001011100010101101100010111100011100100110111100111110010110000010110010101110010110000111010101110011011101100100;
#1 $display("%b", po);
# 1  pi=207'b001110100000011001001101100100100110001010110001111100100000111100010011001100001110010010011010111010101101110101001001011001110000101100100101000000001100111011110010000001001101111011101111000110010110011;
#1 $display("%b", po);
# 1  pi=207'b101001111110010011110111010001011010101111111101110111100111001101011110011011011010101110100110001000011100111001010100001111010001000110100101010100011111010101101000000001111001001100001111000111110011001;
#1 $display("%b", po);
# 1  pi=207'b000010010010100001000100101001110100110111000010011010011110010001011001110011010111011111000101111101011000111110000110101100011000101100001010000110101101000010100111001011001011000001001001001010001011011;
#1 $display("%b", po);
# 1  pi=207'b110100111110011111010011101110100100001001010101100111011110101001000110001101011101011111110110110111111000110111111001101001000001101011100001110010111010101001010011101100000111100111110101100000110101101;
#1 $display("%b", po);
# 1  pi=207'b100010110111000011000111001100001000010010000110110000000001011100001100011100111101101110000101110011000010111000001000011110111010101010110000111101110101110001000010111100001110000110100101011101011100010;
#1 $display("%b", po);
# 1  pi=207'b110001110011100010010101110000011100000100101001011010001011010011110111101110010011111010101100100000001010101011000011111110101010000110000111011000101111011100110101010010001010010101100100011011001000001;
#1 $display("%b", po);
# 1  pi=207'b000011101000000010110110101110100111010111010011011001110011000000111101010111011000001000010010001101010100011010000100000101001011001111011001010001100000100010110001101010011010101111011111010001111001010;
#1 $display("%b", po);
# 1  pi=207'b000011110011000001000011101011101000001111000111010100111000110010000010111110110101100001100111000010110101000111100001111100110100000111010001111010001110110110100010110101011101110001111001010000110111100;
#1 $display("%b", po);
# 1  pi=207'b110000010101111111111100001101011100100110010000111000101100100001001010101111111101011000100001111111110000100000010101001010111101111000101011100110000001011100101111110010001001111000101110101111101100010;
#1 $display("%b", po);
# 1  pi=207'b110001001001110100100111110001101001110011100111010011000111011010101001101000010001111111101101101011001011010011011000010011010001101101011100011100101010101011101110011110000010011111010000001010110010010;
#1 $display("%b", po);
# 1  pi=207'b100000011101011100001110110100011011111010010001001110111001101010010010100011001110010100110000001100010110010110000001011000101101111111001100111010110100000011001000010011010100101100001110111010010100110;
#1 $display("%b", po);
# 1  pi=207'b010011011111011011110001111101101100010110010100010001110100000101101100110110001100101101101000000111011110010010111100111001101111100010010100011010100101111000001101000000011000100100110000010010111000001;
#1 $display("%b", po);
# 1  pi=207'b100001011110111110100100110000111110110101100111111100110110000011111100001000101110111110110011000000101010001111111001101011110001111111011000001001010011101010110000000011100111011011101110110001010011110;
#1 $display("%b", po);
# 1  pi=207'b011000000000100011011011000101100000110110010011110100100000110110000100000010010010010000010000101000111011101010001001010111010001011111000100011010001100011110010111010001110001010110011100000110001011101;
#1 $display("%b", po);
# 1  pi=207'b001101101000100111010000100011111110010001000111001111001010011110100011011110100101001011011101000001110000101010001011010101010001100111100001110000110010010011100111010100111110011100001110111001101011000;
#1 $display("%b", po);
# 1  pi=207'b111001100110110011010100100111001110001000101110010011101110011011111101010100101001110110011010111110110110110010111100001010011001011010000111111110110111001000100010001001110111110001100001010011101110001;
#1 $display("%b", po);
# 1  pi=207'b001010001111101001011011110000001011000111001000010010100111011000100101010101101001110100011101001101000011001101111010011001101100001111101111101011101000100001000001100010111000000110101111110011010111100;
#1 $display("%b", po);
# 1  pi=207'b001011111110000111010110101000011011101101111010111111101010100100110101110001001010001011001110100101101111000100011101101110100011001101110100001100110100111100101000000110101000000110010100010011100000000;
#1 $display("%b", po);
# 1  pi=207'b111000011011101001011001001010001010010100001000011000000110011110101010100100000100000011110110100101101010000010011111000010011110011111000100100101101101001001010100101100110101000010101100101010010101100;
#1 $display("%b", po);
# 1  pi=207'b100001010001011110100011100000010011010001100100001100011101010011111101101010001110100101101001001110110110110100010011101101010010001100100100011111111111011010001111101100101110001011110111011110101111011;
#1 $display("%b", po);
# 1  pi=207'b011001111111000101110100101000111001110100111001010000110010100110010100101100000101110001111010110000101011100011010110000001001100101111011111111000110011010100000110110000001100011101100110000111011010001;
#1 $display("%b", po);
# 1  pi=207'b101000111100111011001101110011010000001101110001101111111100101101111001010100010010011000010110110001001110100110001000100011110001101111111010011011000111001011010011101110111101001101110011000110000011110;
#1 $display("%b", po);
# 1  pi=207'b111011011111011001001101101110000010001110100100000101100100111100000010100001110010010001010100011001010100001001010010101010100100110001110011100110110111100110001111110000100101110110111000111001001001100;
#1 $display("%b", po);
# 1  pi=207'b100101000111011001100010000100100110110100101101100100011110101110111011110101001100101110011010010101101111011010011010011111111111100001011100100100010101111001101100110010000111101110001110100111100001110;
#1 $display("%b", po);
# 1  pi=207'b011111111111001111100000001101000101111100001000010000001011100100010111100000011100001001101001111111011111100000000100000101011001110011111110010101000100100100010010010101101100101011111101110101001000110;
#1 $display("%b", po);
# 1  pi=207'b000011001101111110110011000110110000111011010100110001111100100010101101110001110001011010100000011001111100010100110110010010000010000011001010001001000100111110101110000011001011001011000101100110100101100;
#1 $display("%b", po);
# 1  pi=207'b110100001010111100001000010011001101000111111011101100111111000001111000011100010000110010110110000111101111101010000111111111010110011001010110000100111101000101001010100110101010001100001001101110011101000;
#1 $display("%b", po);
# 1  pi=207'b001110101100101101010110111011001110010001101011000100101111010000010110000111011110111001010000000010111011000010000101111011010110010101001110010111011110010101000010000000110000111000101101011000001111011;
#1 $display("%b", po);
# 1  pi=207'b011101111100101010010110011000000111001111011110010111000111011111000100011000010000101100001001100111111100111010000110111000000101010010001100000111100111001010001101000001110010111001001011001011100000101;
#1 $display("%b", po);
# 1  pi=207'b010110010110111000000000000110011100000101010101110101111100001100111010000111101011001001101011000001011001000101110011001100011001100111001000111010001110011101011110111100100110110010111101001110011001100;
#1 $display("%b", po);
# 1  pi=207'b001001010001001010001101000100001010011100010100011010000010000000111011011001101100010010101101110000000000110001000010010100110001011110001001100100000011000101111010011101100001011000010111101101100111100;
#1 $display("%b", po);
# 1  pi=207'b011110101010001000011100110000010110000011010001111000111011100011011101100111101001101010111001111010111111111101110110110000101110101111001111100001001000010100010010011011100011111100001000100000110010110;
#1 $display("%b", po);
# 1  pi=207'b101110001111011011001100010100101101001111011000100011111101110111111001110000010110111000111010010010011010111110110111110001010100100110110010111001110100001010010010010000001111001110101001011010111111001;
#1 $display("%b", po);
# 1  pi=207'b010110011001101010110100111000000011011001011000001010001101100010011100110001001110000001111111011001100000010101101111000010110000001111010011110110101100000111011101110010011010100100111011110001111011011;
#1 $display("%b", po);
# 1  pi=207'b000110101000010000101101110010110111100001000101101111000100000111010011010010111001001111011100000100101010011011010000010100110110011100010010101101001001101000101011111100101011000011011110101000100000111;
#1 $display("%b", po);
# 1  pi=207'b011010110100001000010000101010101101100001101101000001111100101110011000101100101100101101001110101111000111111111100111111000010101001011010000110101111010010000110010100111100001001010110000111110011010111;
#1 $display("%b", po);
# 1  pi=207'b111001101010111111000110100000110101101001110111110100011101110101110000101000010000110110010011011000001100111101100010001110101111111000111100011010001111010001110101110110101000111011101001011110110000101;
#1 $display("%b", po);
# 1  pi=207'b111010111101100000001000110100100101100010001111000001111101110010101110100101001011100011101010111011010001001000100100000001000111101011111100110000000101001101110101010001001011111110010001010111001111111;
#1 $display("%b", po);
# 1  pi=207'b110110111010101000010000010001111001000011100111111000111111010001001111101010001101010100110001000110111000100000011001110110101001011001010000010000100101010111111011111011000011110111010111011000001010010;
#1 $display("%b", po);
# 1  pi=207'b010011110001011101011111110100101111001000001000100011000111010011001000001100000000110110100000001011010010000000110110000011010110010110001101011000100001001000100110100100101111000111101111011000100011010;
#1 $display("%b", po);
# 1  pi=207'b101100100000011011111001110010101101010010010010001001111000110110111100100001111110011100010100011010000000101000001110011010111101101111011100011011110101101111111010001100011101001011101100000001101110100;
#1 $display("%b", po);
# 1  pi=207'b111001001111110101110110010110111100001000100010111100110100100110001010100001110001100011110110001100101111111111100001010100000011001011111011001110011110000100101111010111001010111011110101101101010011011;
#1 $display("%b", po);
# 1  pi=207'b000010101100100011001000111011101110101111110101000101110110111100000011110110100000110101000001110100101101100101011001110110111111011111010011001111000001111110010110101100100001101101100111010101011101101;
#1 $display("%b", po);
# 1  pi=207'b000000110010110111110100110011001101000110111000001110110100010110100000000000111101100001100001111101101011001101111111111111001111111011111000010000000001001001011110011010111111011101111010000011011110101;
#1 $display("%b", po);
# 1  pi=207'b001100011111000100010001110001011101011011100000010000001010111000110100111100010001101001010111000101101110110010001010110111000010110010100110010011101111000101010000010101011010101111101011100111011001101;
#1 $display("%b", po);
# 1  pi=207'b010011011001010100111100111110011000110011110100011011110011101000011101010001011011000100100101100010100101000010000100011000110000000010111111010111000011000010011000001011110010101111111100010010101100000;
#1 $display("%b", po);
# 1  pi=207'b110011000111001000001000011010100001110110110111110101100101101011011100001100101110000101001000001100111101010100000111011101010010111000100111010010001010000100111011110011110001001110001111100011100010111;
#1 $display("%b", po);
# 1  pi=207'b100111101100001000110011100010101010100011100011001111000101011011101010101000100011101010100101100111111111011010110000011101000111011111110011011110101011000011011111110110100101111010011001100100100000010;
#1 $display("%b", po);
# 1  pi=207'b111101101101111011011101001010110111000010010000100010000111110101101100101111100001001100101011111010010101110001010000110010010011010100001010000000010000000010110001011111001000011011010100111001101011110;
#1 $display("%b", po);
# 1  pi=207'b110111001100110111110010000110001001001001110010010001100001010101011110001111100110101100111110010111100001001110111111001101101110111000100000110110100110001111000001110101000101010110000001010100010111011;
#1 $display("%b", po);
# 1  pi=207'b101010001110101100111110001110110110001110000110111010011100110110100001011100010101011010010100111111101111110000010011101000000101111101101100010100100001010000110010011101111100101010001001010111100000011;
#1 $display("%b", po);
# 1  pi=207'b001101110110000001110111011100101010100010011001001010101110011010000010100110110001011000110101011100001100011110010011111000011001100101011100001000100100110000010000110110001010000100111101110101110100101;
#1 $display("%b", po);
# 1  pi=207'b101011000110000000010110110001110110110010111001100011010000010110011100101101001001001011001100111010000010101101000111101101011100101101101100110101000010000011000111010011011110001010011010011110011000010;
#1 $display("%b", po);
# 1  pi=207'b110100000101011001110111111000001001111101100101111000000100000001000110000101101000001001110110100110101110001000011111011111111000000010101011111111111100100110111011001100100100011011001010101000100010000;
#1 $display("%b", po);
# 1  pi=207'b000110001010011010110001011001100100001101000111011001110010101011101001000100101011100100111100111111100010000000001110100101110001110111110010101101100101010001010000000011111110111010000110001000000001100;
#1 $display("%b", po);
# 1  pi=207'b011110100111000101010000001000010110111011101010011100110101110000010010111110000110100100110111000100111010110101111110111101001010010101010100110110100110011011000001000101100110111010011000010010110000000;
#1 $display("%b", po);
# 1  pi=207'b101001100010111000111110001010000000101001011101011100001001110101000110001111101001010111110000001111111111010101011110000100011001011011110101000100001000000101010000010111111100101101010000100101001001001;
#1 $display("%b", po);
# 1  pi=207'b001111111000101110010001110000001111100001100011111011000001000010110111110101100100011111001000111001001100101100111001011101100110111111001100100000011001110111000110101010110010111000011101110001010011011;
#1 $display("%b", po);
# 1  pi=207'b111100110111101001111011100001001111011010000000001011100111110011111111110110101010010100110111000001111100000100001101011011010101100000011001011100011001100111111110110110010000010010101111101100100100011;
#1 $display("%b", po);
# 1  pi=207'b110100010100101001101100100011011111101101010111101010000010110110011010001001011001101001101100000111000110000101011111111101101100000000100001111101010100110110111011111010100110001111001001101101011100111;
#1 $display("%b", po);
# 1  pi=207'b001000111010010100011110000110110000001101000000010100111010001101111100100111110101001010110001101110111100000100111101110111110111110000100101011000110111011110000010100011111110111010011110100010110001011;
#1 $display("%b", po);
# 1  pi=207'b011000110011110000000100011011000110110010111100000000000000010010100110010011011101011111101000001010010011110100010010010010111000010111001000110100101110110101100001000010100111101011111010000011011001001;
#1 $display("%b", po);
# 1  pi=207'b000001100001010000010111101001000001000000001111000110011101000100000000100001111100000010100000110000110111100101001100000100110111101101001101100111111101001001011101100010010110101001001110111011100111100;
#1 $display("%b", po);
# 1  pi=207'b110110100110111000001110111100100110001010001011010001110011110110011110101101011000010100110110001011111111110010011111011000100110001111010010100100011010101000011000101001110100000101010011001010000100010;
#1 $display("%b", po);
# 1  pi=207'b010100001100001110111010011000011000000010000011101001100010001110110010000101011011010011110100010111110110110001101000110011000101110000000011001100010001001001001001010100010011101001011111100111101000011;
#1 $display("%b", po);
# 1  pi=207'b001010011001011000110111010100000011011111100000100101000001000011000010001111010001010100101110001111010001010101110000100101011010011001110001011111011111000111100100001010110010101100010001110001100001110;
#1 $display("%b", po);
# 1  pi=207'b001001110100001000001011110101010100100011001000110011110111110011011010010101011010000101110100010110101100101111101110011001011001110100111001000101011010010100000101000110100001100010110000101010011010010;
#1 $display("%b", po);
# 1  pi=207'b111100001000000001001100110100100011010001100001100110011101001101110111100001101000001100110011001110111010000000100100000100111101011001101010111000010101001111111101100101100110111100010110001001000001101;
#1 $display("%b", po);
# 1  pi=207'b111010010101000010110000100000111100101111001000010111000000000111100010000011111011001000011100110100101011100011101111000101011000100111011010010011100010010100110001110010101101110110100001010101001111010;
#1 $display("%b", po);
# 1  pi=207'b000110101111011100001001100011111101010011000001111011111101111111111100111111011001100001001000000000000000110010101001001001010000110100001100000101110100111111110110011110000000000001111011101000101111101;
#1 $display("%b", po);
# 1  pi=207'b111001000001001010101010010001100110100001100101100000101100011010111000000010110010010111011000000000110000011000111101001111010010001011000000001100010011111000100100100101110010010101010101010000000111010;
#1 $display("%b", po);
# 1  pi=207'b011100011111101100101000000101111100000110000000000000101001101000101010110111110000000100001011000011011010111100100101011000100111000000110010011111110010010111101101001011011000110011100111000110000101011;
#1 $display("%b", po);
# 1  pi=207'b001000100100101110110101011010110001111111111111100000111011101011100110101000110111010000100011101011101000101101111011111010101111010001110101100100000110110101011111001100101110111101001001101110101100011;
#1 $display("%b", po);
# 1  pi=207'b011011110000110000100010110101010000011010011100111111011100111110111011110111111010001011100100010001110101001010011101001101010010011101101001110000111110100111001100101101101000011111010110011110010101111;
#1 $display("%b", po);
# 1  pi=207'b110110111000000001111000011011101000111000010011010100111001110101101111101100111010100001111111001001010011001000001100101001100001011110111101011101100010001111001111001100100101011010001010110011110001101;
#1 $display("%b", po);
# 1  pi=207'b111111000110100100100000011010100100100011000111011010110011011010000100101101011000001101101111110101001010100011110100110111001100100101000011100011001001111010101010001110000001011110110101011111111000011;
#1 $display("%b", po);
# 1  pi=207'b110000011111100101101100101001100001010010111100101001110101011110010001111111011011011110010001000011101001101010010011011101000111110111000010110010111100110111011110011001100101001010000010111111111000000;
#1 $display("%b", po);
# 1  pi=207'b100100111010101110010111001110111010111000011011100001100110011110010011110011100100101100110111010011110011000011110010001000111010001100011100001011011000111111111010101101111100000010001101111010010101110;
#1 $display("%b", po);
# 1  pi=207'b100110010111011001001111110011111100000101000011011001110010010011000101110010000001111011001100000111010100101111101100110000110100101100100001011000101001110010110010011101111010011110010110010011000110110;
#1 $display("%b", po);
# 1  pi=207'b111010110010101000011110100011111110111000001110000101100010100110101010010011001110110100110010001011100111001110011110110100110100101110110000001001101100110101000010001110000001010100110000010001101101000;
#1 $display("%b", po);
# 1  pi=207'b101101000110100111000000101100010010010110110110101010101001100010011011001001111010100010101110111100011010100110101010100110000000110111010000110010000100110001111000011000101101000000000001100100000111101;
#1 $display("%b", po);
# 1  pi=207'b101110010110011100010011000100111011110011000010100000000010100011011011100000100101001111100100000011000010101010111100011001111111000101101010101011001101100110111100101101101100101101010000000010011001010;
#1 $display("%b", po);
# 1  pi=207'b101100001011001000101111001011010100100101101010010011100101110001111110010110100100100011111011101000000110100011111011110110101101100010000110011000100000000001010010000001100111100100001001010110001110000;
#1 $display("%b", po);
# 1  pi=207'b100001111010010011001011010100110010101001111111000101100111000101000000110010011010100100000000010011010111101000110100111111001000000101000000101110001011011100101010110101001111010100010001001110110110101;
#1 $display("%b", po);
# 1  pi=207'b000011100110101110000000000001001001011100001010000111111000100100010111111001000110101100100011001111010110101111101010000111100001101111110111001100010101111010100111100100000101000001010110011100101110100;
#1 $display("%b", po);
# 1  pi=207'b101110011110001100011001010010111100010001110110011101011001111110101111101010111011110010010111001110011110110000101110011111001110000111110101000010111011011111111101010111100100001111001011111001001111110;
#1 $display("%b", po);
# 1  pi=207'b111000111111110011000101100101000011010001010000100101001101000000000111010100101111000101110011110100100110110111110000010011001111110010011100011110100010010001000010100000110101111100001010111100001101010;
#1 $display("%b", po);
# 1  pi=207'b000101010011111101011000010111001110100111010000110001010111001100011011001100100110101011010110011101011011001011001111111000101010001011100010000110100011110001101101000011001010111000101111000111101001101;
#1 $display("%b", po);
# 1  pi=207'b010111000011111001011000101100010110111111101100110010010101101111000100000110111010110000110010010111010011011001110011001101001101000011001111110001010001100110001100001000111010010001000000101001001110111;
#1 $display("%b", po);
# 1  pi=207'b110101100011100001100101000011101100111111010111101111100000010110110100110010111000001101101011111010101011001111001000001100000010101111110111000111001111000000011100011100001110000101001011100001001101001;
#1 $display("%b", po);
# 1  pi=207'b011100111011101101110111101100111111100100100110100011010000000101001110010000001110110111101111001101111000100100110110010100111010111000100001100000100101111111001101101101000000001101001101100010100100010;
#1 $display("%b", po);
# 1  pi=207'b101111011010110111011010011000011100011111100000001011001011011010100011010100011001101101110010010101011111100111110010110100001101101001101011010100101000110010111000101111111111100110111000101110010011000;
#1 $display("%b", po);
# 1  pi=207'b001011101000011011111101110010111010110101100110000101000101010011101010100011100100110110000111001100110111011000100001110110101101100101000011011010010010111100001111001001111100110110011001100001000001000;
#1 $display("%b", po);
# 1  pi=207'b000001000010111110010001010001010010010011011001101000100100010110110111110101010111001011011000101101011101111000101100110011011101110000110100000111011111001001100001101100110000101101010001000111011000110;
#1 $display("%b", po);
# 1  pi=207'b001100010011111001111110011011100110011011010100101001010001000010001111000100101000111011001001100000011111111011000001100000100000100000000001011000011101101111010100100011101100111011010010000100001100110;
#1 $display("%b", po);
# 1  pi=207'b011000000110001001111011110001110010001101001000001100100000001000001011111010010100110110101011111100111011010110100111001100011001101011010001011101011111101001110000111101100001100100001001010010001111000;
#1 $display("%b", po);
# 1  pi=207'b101111001001010001000000011101110111010111011010000111000010110000010100010000111100111010001000010011100111110010101111110001111000110010111101010000100111011110000100101011111111010110111001010100100010100;
#1 $display("%b", po);
# 1  pi=207'b101011100111010110101101000010101111011001000111011000010011000111110111110000110011010010010100101101100000110101100101011000011010000010011101000100000010110001100111000010000101010010010000110001100111001;
#1 $display("%b", po);
# 1  pi=207'b011101110010100101111100001110001000110101100000011000000111011101111110110100100011101111011100011011001001101010111011001010001101100010010000111010110010101110111000111100110101001101111100000001010000110;
#1 $display("%b", po);
# 1  pi=207'b001001001010010000001110110000011010010110000110111010010000110111011110111111110100111101000001011100000100111011000111001100111100010010000111101011101010100100100011001000011101100100010100111100011100110;
#1 $display("%b", po);
# 1  pi=207'b101101001010000001111111111000011010001011101000001010000100110111000110001011011000101100101011011110101011000000101001100011101000110011101110000101100011010111101100011000101111110100011001001011101010110;
#1 $display("%b", po);
# 1  pi=207'b100111001111001011111001011000000100110111001001110101000101010100101111111001110100010011111010000011010001110000100011101011111010000111101010110100011010000101011001101011101000100111111110011101100100111;
#1 $display("%b", po);
# 1  pi=207'b010010000110100100010000010101001111111110011111001010100011011001111111110001011011101101011000110010001001111100100110011010000111001111000000001100010100010111110001001101001001110111011100010111110101101;
#1 $display("%b", po);
# 1  pi=207'b001010001110101101110010000101000111000110101100100101110101011001101001101100100000100100011110011010101000101110110011000011000011101100000101010000100001001011010110000010100111001111101001101000100111111;
#1 $display("%b", po);
# 1  pi=207'b001001001110000001110100111101100011011010010111110001000101111101011001111100011001001000000101000110100011100010010011111011111100100100000110000110011100010100100001111011111010010000111010111011110010011;
#1 $display("%b", po);
# 1  pi=207'b010100000101011101101111100001100100010110011101011100111101000010101001010100011011001011111010000101101100000001011001000100110101110111011001001011010010101000011011110111000110011010010000101000010000001;
#1 $display("%b", po);
# 1  pi=207'b101000011100001010000001111001001100000111111010010001111010011111011101011001011010110010001101010011100111110000001110111001100100011000011011101001010000101011011011000101100110101100100100111111111001111;
#1 $display("%b", po);
# 1  pi=207'b011010101110101111000100110111111010011001000000011110000011101001101010001010101011011111100111101000111000010100000000000010110001100100010010001111110101111001001100010011011100111110110010101001001100100;
#1 $display("%b", po);
# 1  pi=207'b010011111101010000101010100011010101011110001011110101110100100010010111010010101001100111000110110111100000001001111101001111101010001010011001101111011110100001011101110100000010111010101101000101110000000;
#1 $display("%b", po);
# 1  pi=207'b000111000110110011100010011010101100011111001110001000011101100001110101110001000001100100011001001001000111100111000111011001001110010000000001110011010010000100100111010011000100000000000110011001101110011;
#1 $display("%b", po);
# 1  pi=207'b010111001001101100000010010000000110001011010100010101101100010001010000111011111001011001111111011000010010010110001101101111011000101100110001101011000011110010010001001100010101010000000011100010001011000;
#1 $display("%b", po);
# 1  pi=207'b001001000001101000001011111111110001111001111001010011011001110011100000101110011010000011010001010111011101001010010011000010111111101000110000101110101100011110011111000101110010111110101111111000010101001;
#1 $display("%b", po);
# 1  pi=207'b001010101010100011101000000010110011000010110011000000000010101101101101000100011101011110101001111100111000100000011001001001010100111100001110110001000001100000010111000110111010101010011001010110001101111;
#1 $display("%b", po);
# 1  pi=207'b000110010100110100010110101100100011110111000001111000010010001001111111110000100110000110001101010000000001110110010000001010100111101100101100100000001110011111000101100001011011001011001000110101100100011;
#1 $display("%b", po);
# 1  pi=207'b101001001010101100011000110011100101011000010110011011101101101010100010010100101111010110000001110010000001111000100011001000001010010100001110101111110010001111100011011001001011100111100111011111101011000;
#1 $display("%b", po);
# 1  pi=207'b011111111011100110001001000110100110101110111100101001110100101001011010110101001100110001011011110000101010010001111100001110111001000010110111110001111000101000000000101001111100000101101001111111010101010;
#1 $display("%b", po);
# 1  pi=207'b110000000011001110110001101000110011010100011001110011101001110011101101010111001100000100101011000101110100100001010101010111010111000100011011000110100000101101111001101001110100111110101100110001111011011;
#1 $display("%b", po);
# 1  pi=207'b000111101011000011101001100110101111110110111001010010010001100111010001010011100110101110011110101101110111011110011010101010000110001000100100011010101000111010101001000010011110110010100110011000110111001;
#1 $display("%b", po);
# 1  pi=207'b111110100111111000010110110101010010111100101110000101010000000111110010000000010110101000000111111000101111011000101001111111001001010011110100010001001111101001001100001101100010000010011011001011110101111;
#1 $display("%b", po);
# 1  pi=207'b111000101000100011101100001001111000100010000101111111101000000010000100001011011100000111011011011000001001100000000011101001110100011110011010010010011100110010000111110100111101111101101000011111000011000;
#1 $display("%b", po);
# 1  pi=207'b011111010011001101001110111111111100100100100001110001111001100111100000010100111111101101001110111101010110110010101001101100011101111000000111001011001011000001101010001101000010010100000010010101001011110;
#1 $display("%b", po);
# 1  pi=207'b001011010101110111010011001110000000110101110100011101010100100110000101011011010010101100110111001001111100101010010101110111101001100000011110001111001001011011100101001011101101100110111010100010101101100;
#1 $display("%b", po);
# 1  pi=207'b011100000111001011101101111010111110000010011111111101011011100000011000110100001111011101100100100010111111011111000011100110101010010100100010011010011001100010110010010101000100110000010011100100011010111;
#1 $display("%b", po);
# 1  pi=207'b011011110101001110100000001111100010001010110101100000110111101000110011010000111001100011011010010111100011001010001000001010000010011011010000100110111100100011111111001011100101100010001111010100001011001;
#1 $display("%b", po);
# 1  pi=207'b101001111100010011111101011001110110000011100111011101101010110010011011000001110110101101111101101100011001011001111011000111100101011011111001100010001011011101110111111011000011110100011101101111001010100;
#1 $display("%b", po);
# 1  pi=207'b111111011001110111000101010110111010011111001011000110011111011100100010101011011000011110011000101101011101000001001101110011010100011100000010000110000001000001001100010010000110000000001011000110110101111;
#1 $display("%b", po);
# 1  pi=207'b001110010100011110101110110000010100111111111101011111010101111111010000000001100011011000010000000111011011110011001110010010110110110001001010001010010111001111001000001000010111100000011011111000010001111;
#1 $display("%b", po);
# 1  pi=207'b110001000101001100011010000110000010010010111000010010110011011111010101101011011001111110111101110111000010011001110101101101111111101110111101111000011001011100101101101100100001001011011101000010000101110;
#1 $display("%b", po);
# 1  pi=207'b110111101011101100011011110110010111010010010100101011010110001101100011001111010100101101100111001101001000000001010001100000100101001101100110101000110000010000110100110110010011100111101010011011001111111;
#1 $display("%b", po);
# 1  pi=207'b100110011110000011001000100010011101000000101001100100100011011111111011010000001100001110010011000001110111111011000000111000011111011110001101001001001001111001010000001010000010100111001110011011010101001;
#1 $display("%b", po);
# 1  pi=207'b100001011111011011001111101101100001000010010001001010000111011010011000101001011101101110100101101110110010001000001101111110110010110111011111101010000000110010000111101110101110010101100100101010011010001;
#1 $display("%b", po);
# 1  pi=207'b111010000011100111011101111101011010010111110100110101011110011000110110001000011111110100010110001111000101000000011101101101101001010110001010010111000100111000100011001110101011001011110101011001000101110;
#1 $display("%b", po);
# 1  pi=207'b010111001011010010011111111101011011110011101111011111011111101111011011100101111011101010001011011000010001101001001101110010001110101011101011111111000000010110101111111001010110100011010000011011011000110;
#1 $display("%b", po);
# 1  pi=207'b000001101011001001101101100101100100111010101001110100111000010111111010010010011110100001111100101011100110011011010100111001000101001111110101011000000010111100110100010011101101010011110011111101000000001;
#1 $display("%b", po);
# 1  pi=207'b100001111101110010010100100101110111000110110001101011001010110110111110100101010101110101111010010001110111010101000001000011011111101100010110110101011100111010001000111101100010101110001101111110011100101;
#1 $display("%b", po);
# 1  pi=207'b010000000001000111110011110111010100100010010101101100000011000000010110101001111000110011111011010101011110100000111100001100000010011001000010100010100001011101010101001010110110001000101100001110010111101;
#1 $display("%b", po);
# 1  pi=207'b111101101011010101101010111110001101000001000000001011111110110000111001100100110010000111101110100011010010100110110000110100010011011111000000101101110101110111111010010100111111000010111010001101011010010;
#1 $display("%b", po);
# 1  pi=207'b000011001010100111011000000010111011001100010010001000101100001110110100111001100100001011111001101011111000101101110100101111111100101101110001111101100110100111010101001111010110010000010001011010110111010;
#1 $display("%b", po);
# 1  pi=207'b101001100000100110101000011101001000110101000000000000110110101110111001011011010011101100011111001101101100101000100001111000110110101000010110000001011001010101111010100000101111110000011111110110000101111;
#1 $display("%b", po);
# 1  pi=207'b111000111001100100001011100000010100101011100010010010001000010000110001011001000001111110010011100100111110000011000011000110010001101100110010101000110110100010000100110000010101100101000010001010110100111;
#1 $display("%b", po);
# 1  pi=207'b001111111111000000110000000001010100111101000111110100000101011000100011001110111011110111000000000001011111110001100111010000001111111101000111101101010000111010101101100110010001011011101110110000010101111;
#1 $display("%b", po);
# 1  pi=207'b110101011101110100000110111001001111111110110101110100000101000111001111111010100110000100101101110011100001111000110111011001010000001110001110101101011111001110011100001111100011101110000010100111010111011;
#1 $display("%b", po);
# 1  pi=207'b100001111010100101111011001010110100001100000010100110010001011100000100000100101101110110101000111100001000000101000011111110001011000001100000000110110011101000000010101110000010111011110001000001000011101;
#1 $display("%b", po);
# 1  pi=207'b111101011111010100100011000110111101000010000101000111100010101111010111000011000001001111100010001001111011101001001011011100101000010010001000010111110101000011100101000000000010110011101101111001101111011;
#1 $display("%b", po);
# 1  pi=207'b001000110001110110000000010110110100110101011001100010011101101101110000110101011000110111101101010000010010010010010001111010001010110010011110010101010001010100101010000010000111011111000100010110011100111;
#1 $display("%b", po);
# 1  pi=207'b010101001101100111101001111011000010010110010100110000010010100100010010101111100100011000100101010100111010000000110011001011011111101100101100100100010111001001000000010001011010101110000111101101000101001;
#1 $display("%b", po);
# 1  pi=207'b110101110000010101111111100001000110110111011000110000110001000010111010010010010111101101001101010010111000111010101111011000011100111000101011001011011101100101110000110110100011011111010111010110111010000;
#1 $display("%b", po);
# 1  pi=207'b011010111100111001101000100011101100110000011001011110101010101011000101011110000101001010100011111110001101100101101011001010110101111000010000011100110010001100011110011100100101001011110111010101010101010;
#1 $display("%b", po);
# 1  pi=207'b111011011111110000111011100111101101111100011001111001101101001011000100101001011010111001101011010110010001110000110111001011101010001101100010000101001100010111100000010101110010000111101101011011101000111;
#1 $display("%b", po);
# 1  pi=207'b001101001100001111010011111001110011011001110010010011010110001100001001100000100111000000111100000111110101011100011110100111101110110101011111111001010101011001111111111011011111101010101101110101010101001;
#1 $display("%b", po);
# 1  pi=207'b001101100101000001100000010111110011101101111011101010110110100011010010100111011001000101101011111101010010111010001010100111100100010110010110101010111011100111110011111010000110010110010110001011101000000;
#1 $display("%b", po);
# 1  pi=207'b101000010110110110101101010011110000111111110101111100101110101001011001000010000111111100010011111101011101111010101000111111101010100101100010110111011100110110101111110001010110110010110000101011101001100;
#1 $display("%b", po);
# 1  pi=207'b100110100000011010110011001101011000110111101000100000011111001100110001110000010010010100011001100001100010100110111101110101100100110101100000011100011001110110110110000011101011100110110000001000001111010;
#1 $display("%b", po);
# 1  pi=207'b011100010101100110001110110001001001110011000001100101100110110110110011011011010010011000101011101110011011011001101000110001011001100000100010110001001010100010001001000110101101001100010110000111100101100;
#1 $display("%b", po);
# 1  pi=207'b111011111000100010101011000001011010000001001100010101110101110100111001000010000011101101101110110001100010110110011111000100101100001100101100110100000110101100010001001010111111001111111100000101001000111;
#1 $display("%b", po);
# 1  pi=207'b010010101100101000101100110110001000110010110111100000101011101110110011111100101100101010101001110110000110010010110110100111010110100110111100110010111101011111111101111011101010000000001001001100010011001;
#1 $display("%b", po);
# 1  pi=207'b000100100001000111111110011101100000111111011111011010011010111100011101110001111111010101010101100100000001011100001110010001100011111011011110011000100110011110100101110101001101110010001110001010000001000;
#1 $display("%b", po);
# 1  pi=207'b000010111010000001011010011011111011100000001101101001110101101001000001011001001101010100001100110100101100110010111100110001001100000111001011100100100011110001110011011001110001010100101101010101101000010;
#1 $display("%b", po);
# 1  pi=207'b111000010000101001100011100111101100101011000100011011111000010011010001011100101001000111100101001110100000111000001010010100010100011110111001001001011000000110111011110000101011001000101110010111001110011;
#1 $display("%b", po);
# 1  pi=207'b100000001101000111011011000011001011000101100011101011001000111010010101101010010011111111001010100111000000011000110111100011010000010001111011011000001100111000100011110110000100101100011001111010110010111;
#1 $display("%b", po);
# 1  pi=207'b010111110010110100111100100110010110001101011011101000010110110111001101001010001000101011000111111010111010011101011111000011001101100111101101111101001001001010001001010001110001000110001110001111000010101;
#1 $display("%b", po);
# 1  pi=207'b010011010001110101100010010001111110000110011001101110111000100010001011001101111101000001011000000111111110100010011000010110001111010110011111011111111011101010000010110100101100001110111111111101100000001;
#1 $display("%b", po);
# 1  pi=207'b011001110111100100011101110101101010111011110100010001111100101001101000011100111010011010101011100111011101110100100001101101011110110100101011111101010110011111000000000110110010001111110110000110001001000;
#1 $display("%b", po);
# 1  pi=207'b110101111010111010110010010101000100110110110000111110000101010001001010001011110011110011101111011011010000001110000010010000000000100000001101001001101000110010001001100010111100101010101111011101001100010;
#1 $display("%b", po);
# 1  pi=207'b100000011011110001110100000001101000100101001001111101001011011100101100011111001111111010100110001000111101010010000110010111110110010110110100110011011001000110100110011011100001010101011100110000110010101;
#1 $display("%b", po);
# 1  pi=207'b101011100110110011001110100000010100111100100111000000110110110110100100101110100001000111000000001010111111001000011010101011011101011100101000001001110011011100101001011110111110000100100010100001010011011;
#1 $display("%b", po);
# 1  pi=207'b011101011000001110010101100101101001110101101101110100110111010110110111101110110110001100010110001000010100000100101001101000010000111101000111000111101100011000000001001010100101101100101111110010010010001;
#1 $display("%b", po);
# 1  pi=207'b011000110101001101010000111010101110000001001110001100100100110010000010111011110010101001000000010001111100110010010001011000101011001001110010000111100010010011101010010010000100011110001000010000100100111;
#1 $display("%b", po);
# 1  pi=207'b010011011111000100001100011011111100110011011101111001101000001101100010011010100010110110000000101111100000010000100100000111111001100000011100001111101111100110011000111000000111110101101100011001101000100;
#1 $display("%b", po);
# 1  pi=207'b011000000010010111110111001110101000000100000001011001010001100010010011011000101110001101100111100100001001000000101100001101000111111001101000001000011100100101101001000011000001011000011000100101101100101;
#1 $display("%b", po);
# 1  pi=207'b001111001001111011101101011000010011001001010111011001100011111111011111100101011101101110000010001000101010000011001001000001001111110100001101101100100011100011011100000111000111101010001111100011010111000;
#1 $display("%b", po);
# 1  pi=207'b111011111110011011001111010010010010100011001000111000011010101000111000001111110011111111111111110101000101111111011111001111101100110000001011111000010100000110011011100001010101000110110001000001001010100;
#1 $display("%b", po);
# 1  pi=207'b010011000101111110010010110101111000100100101010001001001100101001001111101111001101010110000000100000001101100001010010000100000101101000001100111000001011110101100000110000111100101000101000011000001100000;
#1 $display("%b", po);
# 1  pi=207'b000001101011100111100110110011001101110001101101010001110000100001110101010001111010110100000001110101001101110110011101111100100101110110110101001110011111111100011101100101111001001111101011101100000101001;
#1 $display("%b", po);
# 1  pi=207'b011000011100100101001000101100011101001111000100000101000011000110110001110000111010110000010001111000000100000100101101001110000001111110110011001001010000100101110110010011011111011111000000111101101111001;
#1 $display("%b", po);
# 1  pi=207'b011000101111101000011010000111000001000100110111010111001111111000100101001110000111001001100101110100000100010001110100110100011100101111000111001000110110001101101111001100010111101000001011111100100100101;
#1 $display("%b", po);
# 1  pi=207'b000001111010111000001100101111000000100011010100010111101011011001100010011111001010100101100101100000101110000110001010100011110000011111111100000001101110011111001101101001001000111101100010000000001111100;
#1 $display("%b", po);
# 1  pi=207'b010000001100101111001111010101100010011001011100111010010000001011011001100110110011010011010010101111100111100001000011101011100110011001010011100100111000111001110111001001010110011001110000010101111001101;
#1 $display("%b", po);
# 1  pi=207'b100000011001110001000001010000010011110001100011011101011001000000001111101111101011010001111000011110111001011010101000001101100010000001101000000011001010001100011111011011111000010100010000101100111100011;
#1 $display("%b", po);
# 1  pi=207'b000000011000111011110011111000110100011011110110100111001011101111011001110001101111001001111001111101111101010110000000110000100110100001010100011011001010101110010111100101111110100001000100101011000101110;
#1 $display("%b", po);
# 1  pi=207'b010011100000000010010111011111011010100100000111001011000101000110010110000011000111100000000000101100010011011001001111010110101110100010010101001111111001101010101111101011110111111011000111111001100110111;
#1 $display("%b", po);
# 1  pi=207'b110110110100011010011001110111111001111010110111101111011011010110001100001010010010100001100111111111110011001011100001110000110010111000001011111000110001111110000000100110110000111100011100010001100010011;
#1 $display("%b", po);
# 1  pi=207'b011101001000111000010001001000011111110011011101001111100100100101011000110000010010101010100101011010101011101100101101110100111001000110110100111110101100110011010001000110101110101100011111010100110001011;
#1 $display("%b", po);
# 1  pi=207'b000011011001101000101111011011000000001001110100110001111011011101110110111001001110100111101010001110000101000001011001111110101111011110011110100110001110011010101001010101100001001010000001100101100010010;
#1 $display("%b", po);
# 1  pi=207'b111010000000110111101110000011000001011001000011010010000001001011101111101111110010010111101010101100001011111100011110110101001011110001000110101101011111111001100001000001111000110010111010010000100001011;
#1 $display("%b", po);
# 1  pi=207'b100011000110011010001101100001111011111110100011011100110001011001001100101100010001011111111100001101011111101011110101101000100101010110101011010011100101110010001011001000011110000011010010111110000010110;
#1 $display("%b", po);
# 1  pi=207'b101101111101101010010111011001010000010000101001111110000011000101101100110001001110111010000001111101110110000101111000110010100100010011011011011001000110100010001011110111011010111010000111100011011100101;
#1 $display("%b", po);
# 1  pi=207'b100111110011101000100100011100101110100100010010001101110100110001110010011110001101100000111101001011011101001111101100011001111110110001010100011100010010101111101000100110010011001101110001000010010101001;
#1 $display("%b", po);
# 1  pi=207'b000011111000010100001011001010000000000110111011110111010011100001010101011011010001110010000010110000000101010011000001000111100000110111010111000111001111000110001011111011101110001111010111011100001001010;
#1 $display("%b", po);
# 1  pi=207'b010100110101011110001111110001000011000111001001011111000100011110111001010001001010100111100100111101001110110101000110000110010101110110101101111001101001110111010000001111000001010111111001010000011011011;
#1 $display("%b", po);
# 1  pi=207'b011001011010010110011111001110111110110011110101101110010100101110101011111100100011001001100000010101101100000001111010101011001010100011110110110001111111111111100011001101100000100111000001100111011111110;
#1 $display("%b", po);
# 1  pi=207'b011001111110110100000011110100001001011010111110110010101010111101011011010001000011001001101000100011100000001100000000010110110010111111100000111010010110110000000110011001101000001100110001100111110111001;
#1 $display("%b", po);
# 1  pi=207'b100111011100011111100000100011001100010100111011110010001111110001011111101010101011111111010110010010111110110000101001110110100111100111011001110101001110001100111110001000010000011100000001110001010110110;
#1 $display("%b", po);
# 1  pi=207'b100010101101011010011001011011101010110001011101101001110011000111111010101000011001101000001011110101110001100101100000010011011100110010111101111100111011111101010101010101101111100111100100000001101000001;
#1 $display("%b", po);
# 1  pi=207'b000010111010111000001101001010011100110001011110110011100110111010000101010100100110110110110000010100100110110100010000000111111110011010001101111010101101101000001010010010010011101101010111000101011101110;
#1 $display("%b", po);
# 1  pi=207'b010100001111011110010100011011110101010001101111011111110111100000001101000010101011110010100101101101110010001110000101010011001100001101011010110111100100011111110111000010110000100101001110001101001010001;
#1 $display("%b", po);
# 1  pi=207'b101100110110001110000101110111111111100111000100011010101101001001101001110001111110101101010111100101100011101101000110111110001101011110000100001010110001101001111110101011011110001101000100110011000000011;
#1 $display("%b", po);
# 1  pi=207'b111010111111110011110000010110111110101100100111011010000010011010001000010010011110001001011100101011001000111000011011100000010000010000111011001011010011100111010111100110001001100011010001011101111001110;
#1 $display("%b", po);
# 1  pi=207'b111111100001011000111101110011010111110111110000110011111100110000110100001010111100110111111100101011101111000111000110010011101010101001111101010000001001011111110110101001001111101010010010100100000111100;
#1 $display("%b", po);
# 1  pi=207'b110000100010101101011001110000011111110011011001010111010110011001111100000010011111001010111101010101101000001100010000101111100001010100010000111110110011011010110011001000001100001111000010011010101010111;
#1 $display("%b", po);
# 1  pi=207'b100010011001101101011101010011100101110110010111010011010000001001000010010001111000011101101111011000100110100001001110100001100010100111000110000100110101111111010100001111100101000100100110111101000001101;
#1 $display("%b", po);
# 1  pi=207'b110111001001001101100111011001101100001101110111100010111101111111000000111110010101000100010110000100011000010010100000000100000010010110100101001110011101000111000010000110111001000110110001100011001001100;
#1 $display("%b", po);
# 1  pi=207'b010111000000000100100100010110101011001001011100110010001110001101001110000101111000011100000010111111010010111001000101001100110011110110101000100110010010110010001010000011011000010100010110111111100000011;
#1 $display("%b", po);
# 1  pi=207'b101110100000011110000010101011011001000100100011100101001111100100111111111011010001101111110011010010101010111001100010010000101001011101111010000010101100111000000010100001110111100101110101111011010101011;
#1 $display("%b", po);
# 1  pi=207'b100000101110100011100011100000001111010001110011010010100010000001000101100000010001100111101010100000001001110110010000110101110000101101100110000000000001011001110111101010101110101011011111111101011010100;
#1 $display("%b", po);
# 1  pi=207'b010011110100100100010101001110101000101101110111110001101100110001110010000100111010001001000101100111011001110101111011000000001011001011001001011000100101010000001010001101001100000111010001001011101101100;
#1 $display("%b", po);
# 1  pi=207'b111011000010000110011001100101101111110101001111110101010100101011011100101111011110101100101100101001111010101111100111000100000100000010010001101100111111011000100011001100011111100000111111010111001001111;
#1 $display("%b", po);
# 1  pi=207'b101110100110111101110100110100100100101111011110111001010001110111010101110001000010000111000110101100001010011001010010001110100111000010111001110100000100011011110111100110101011001100010100101010010100010;
#1 $display("%b", po);
# 1  pi=207'b110110110110010010010011110000010011010111100101010101011110000010101101111101101000111000101101111011000010010001010001101010101000001111111001111001000100110001100010010111110100000101001110000010111010110;
#1 $display("%b", po);
# 1  pi=207'b101000000011101101111010001101011010101011100111001010110010011100110100000110001101010011001001011111010010110100000110101011100000010101110000111101100100010001100001011010011010101011000011110011100010011;
#1 $display("%b", po);
# 1  pi=207'b101001001100010001011010111111101101011110011100011110001100000001100001101001000101111110100011111100100001110000111100100000111110101110011010011110000000101010110001011011001110010001111001011000000010000;
#1 $display("%b", po);
# 1  pi=207'b000011001011100110100010001010100001111011000100100100001100100111101011110101110000100101001000111011101111010110101100001100000100010010001011011010110011011100100100000100011011110011110100110111111000000;
#1 $display("%b", po);
# 1  pi=207'b000100100011100100010110111100100100101001001010110010000011001110001100100101110001010001100011010011100011101111100000110110110110001100000000111110001111001110000001101110010101101100001100010101101111011;
#1 $display("%b", po);
# 1  pi=207'b000011100000110101001011001101101111111100000101101100101100101110001001100101000101001010101011011101101011011011010010011000011011001010000000110100110111110001010100100101110111111011101111000001101100111;
#1 $display("%b", po);
# 1  pi=207'b000101010010001110000100000010111010011001010001111110001101010101100110101111100010011000010101101000111110100101001100010101101011100011010110110111000101101101101001111110011011000100000101000111100111101;
#1 $display("%b", po);
# 1  pi=207'b101010110111011100101010011001111011000110111111100000101111010010111010101111011100111110101011111001100110000000111000001011000000010110001100101011011100010001000110010110100011011100101101011101101110001;
#1 $display("%b", po);
# 1  pi=207'b100101000111111011111001100111000010101000011011110010110111000111001000101001111001011110101100110000110100111010111010011001000110010100101101010011010000000101000110001100011000111111110101011110011001101;
#1 $display("%b", po);
# 1  pi=207'b111010110010110000101101011001010010100011010111101101001110000001001101110010001000101011110001000110110000100101111101001100000110000001101110001011000001110111001010000000101101000000111101110100111011000;
#1 $display("%b", po);
# 1  pi=207'b001001001110101010001100100011010000101010101111111110000111000010110011011101101101010000111101111001100110110000000101101100110011000111010100001010111000101011100001011111010011100000011000110000000100011;
#1 $display("%b", po);
# 1  pi=207'b110100000010100100100100010101000001001110110010001111100110001001110100110101101110111011001100100001001011101101011011000111000001100010101111000100000100101000000001111001010010000001111111101110011100100;
#1 $display("%b", po);
# 1  pi=207'b000000111101110111100111101000111001000010111001101001001001100101000000110000101110000100001100100010000000111000000011011000000010010011000111010101010001000010010001011011110011101000100100110001011110000;
#1 $display("%b", po);
# 1  pi=207'b100000010111011100111101011010010010110100001001010110110101101111010010110111010100111011111111011000111100010100010000011000110001001010101110011100110001110111111000101101000111111110100011001110110101010;
#1 $display("%b", po);
# 1  pi=207'b000111110001101011001110111001000001100101100000011000010001010010110110101000111100100001100110000110111100010011010100110101111000100000101110011101110010011111000010010010001011011011111011110011011100110;
#1 $display("%b", po);
# 1  pi=207'b100100111101101101101111010011111000100100001101111011101111001011001100101011110001010010011001101101100100101010110001101001101001011101000110001110101010111001111111011011100100111101110111011011110110101;
#1 $display("%b", po);
# 1  pi=207'b111001111001000100100000101101110100010100000010001111100111011000000100110011110010001111111101101110011110010101001111100000110110011011001011100010110011000100110101100110000100110101100101101000110001010;
#1 $display("%b", po);
# 1  pi=207'b100011101010000001011101011010000000001100110110101100111100111000101010000101100000000001000110010100001101110110001101000101000110011111111111111101010111001011010110111010011010101000001001101111101011000;
#1 $display("%b", po);
# 1  pi=207'b000100001101110110011000001011000000101000111010111110110001000110110011001100111111011111110011100001110001101101000000101111100100000110011000111000001011101100010000011110100011000000011100111110000110011;
#1 $display("%b", po);
# 1  pi=207'b000000111101011111000001100010110101000010001110000001100111001100010100111100011010001110001010000010110110110001100100011100100111101100010111000101001000011011101010111110101010111010000001011011010011101;
#1 $display("%b", po);
# 1  pi=207'b101000011110110001110010000101101000100000110101000100010100011001110010111100001110000110110010001010011010001000011110000010111011001100011011111110111100100000010101001111011111011111001001111111010010000;
#1 $display("%b", po);
# 1  pi=207'b111000000111010100000111101010011101011001101111110100110011110010111001101110111101101001011001011010000001010011111100111010100110101100100001000011000111111100110001010001110010111011000110000101001000001;
#1 $display("%b", po);
# 1  pi=207'b001010110101100010001011111111011011011101111100101010011001111010101000001010000110000001000111011100110010010001011000101011010000001111001110001101000001100010001010110100001101110010010001011011001111001;
#1 $display("%b", po);
# 1  pi=207'b001010111010000111010111001011011001000101011111101100000101001110001101011111001111001011101000111001010110011100101010011001001110010000010101111111001000000010011001111110111111101101011111100111010100111;
#1 $display("%b", po);
# 1  pi=207'b010001000111101011000110111101001010001100101000010000000000101010011001010110101011110111100011010000111111111000111000011100000111100011101000101100101000001110001110011011101000000101100101000111111010001;
#1 $display("%b", po);
# 1  pi=207'b001100111110100111110101010110111000000010000001001110110001011011011100111010110101111001010100000101001011011000010011111101101001110011000010000101000110000000001000000001000001111111101111000100101010101;
#1 $display("%b", po);
# 1  pi=207'b001001010001101010010010110000100010010100111101001011000111011111101000110100010011100001000010111111110110110110110000011010110111010110011101111010011110011001011001110011100111100001111001101001111000111;
#1 $display("%b", po);
# 1  pi=207'b001101011110000110011001001110001001111110111100001011110111110101111100000010011111001110100101000010010100100101001010011000001001010000101001011110010111001011000011001110100001001110010000100000000111101;
#1 $display("%b", po);
# 1  pi=207'b001111100001100010100110001001001111110110000010000101011011111111001101000010010000010100110111010100001101000110100000100011110101001100110011101101110110110111000100010000110011101011111001010010100101010;
#1 $display("%b", po);
# 1  pi=207'b000110011111101000110001000111111111000001010011001101000010101010010111101010111000010100111010011001111100101100010001100110110111011100110111111011100100110000111111000011111000100000111010101010100001100;
#1 $display("%b", po);
# 1  pi=207'b111100001011000101101010000010110011000100011000111000100001101000110110010000000000111000011100100100100001110110101110011000111101011010100001110010111010111000000101110001111010000101111000101111100100111;
#1 $display("%b", po);
# 1  pi=207'b111001000010011111100111010001101111010111100100011011000010111100111000101110110110011100010101101101111110011100100011111000110001111100010111010010100010000010100000010001000111011101111101010110000101110;
#1 $display("%b", po);
# 1  pi=207'b110101110000101001111000010010111010001011010101100010010010011100010001001011101000101111111000001101100110011110001110011010001010010011100101000000000100011000110001000010000100000110110101111100111110110;
#1 $display("%b", po);
# 1  pi=207'b011100101100011110111110010000110000101110111000010000010010010000000100010101010001111101000111110110011001111010101001111110011101101011100010011100101011111100111000001100001010010011010011111001111111101;
#1 $display("%b", po);
# 1  pi=207'b000011100011101001010111011101111110101011110001001111110001110010111111110000010010010000000011010100101010100111001011001101011101010000111110000011011000011000100101011011111010011111001100010001111011110;
#1 $display("%b", po);
# 1  pi=207'b111100010010001101100110011101000000011100101000100000100010010011110001001100011100011100000100010111111000101111110100110110100000101011001011011011101001010110100100010100010101001001011100001010111111110;
#1 $display("%b", po);
# 1  pi=207'b111101100010110100110100101101010110011001101101000011100001101000101100100011101000110001010011110010010100010110111001011000010011000010001000110011011101011000101000001000010011101111000011110101100011100;
#1 $display("%b", po);
# 1  pi=207'b110111000111111010100110100101011100010000101001101101000100001101011111011000101000101111000010001010110001100001001001101010001011001111110001100101011110101101011100100111111111100101110010010111001110001;
#1 $display("%b", po);
# 1  pi=207'b000011111110010001101011011011000011010000001110111010011100110111011000010110011110000101110110010000110110111111010101011111111001101110010011100000010111111001001111011100111100111000000000011111001101110;
#1 $display("%b", po);
# 1  pi=207'b111100110010001111101100010110110101011011000001110000011010011000010000000010000111010100001101001011001110011001000000010001101100111111001011111001000010011101010011001010011010111110001011101001101100000;
#1 $display("%b", po);
# 1  pi=207'b000111000101001100010001001110111000100100011000010101110011000010000010001101110101101110111001011011000100010001111110111001000110001000011011011011000000110101111110100010000000011100110111110011110000000;
#1 $display("%b", po);
# 1  pi=207'b010001011010111001111001010110001101100111101010011101001101001011111100101001101010111010100011101101111010000010000101000100001000001011110000110110111001000101100100000111011111111101000000111101110010001;
#1 $display("%b", po);
# 1  pi=207'b100011101010100010110110001000011011000110110000001111111000101011001000000110100010000110101000110001101101010000111010111111001100110111010111110110001001000011100010100110011101111100111111001101101100110;
#1 $display("%b", po);
# 1  pi=207'b011010011101000010000101000101100111001110000101000010110111100010001000100110110000100101110000011010000111001101000001110010001011001100101101101100001010101101001110111110101011111011100111110000110010101;
#1 $display("%b", po);
# 1  pi=207'b111101010011000011110110010011110010100011011100101010001010010111110101111101000100100001010000010101101010111111110100010000100010010001001000000001100010001100101100000010001000011100101101010111010000100;
#1 $display("%b", po);
# 1  pi=207'b111011001011000011011100110011010001010111110101000000011001001001111110010010000110100001111000101011100001101000001001010000001000111000000110111011011101000100100101001110001011101010100001000010001100000;
#1 $display("%b", po);
# 1  pi=207'b100010111011011010011010101111011010010110001100000001010100111010001010000011000110001100110000000110000010010111011000101101001101101010100000011111111110011101111011011010110110100010011001011011101101000;
#1 $display("%b", po);
# 1  pi=207'b111100110111010010010111000110010000101011101101001110010001011001011011010001100010001011111010101101011110010101011111100110011010101011111000000110101111100110011110111000110111000010101011100001001011001;
#1 $display("%b", po);
# 1  pi=207'b000100010111110110111110000111011100111101110100101100110111101001101000001101100000100111111000101010001110001101010011001110111111110001100001111110011011110011100010110010101110100100101101100011111001000;
#1 $display("%b", po);
# 1  pi=207'b010100001110111110101101100000101010111100110011010111110010111110100111010101001100101111110010101101000101001001000011111101110000011000100100011010100111110110101011011100101011101101010001011011110100010;
#1 $display("%b", po);
# 1  pi=207'b110101001100011000110111110000000001000111001110110010001000001110010000001110110110001001010101100000000000011111111011000001111101000001111110001011100001010101001010010001101000101101101010111101000111010;
#1 $display("%b", po);
# 1  pi=207'b100001101100001101110001100011111111100100101011001111001101101010101110000011011110001011000101010011000000101010101011101100101010110110111001011000011001010000010001001011000111101101100110100001001011111;
#1 $display("%b", po);
# 1  pi=207'b010011100000000001011000101000010010100100000010000011011100100000001110000110110100110110010011011100101000010101101001111110101010010100010010100010011001110101101010111101111110110110010111111101000111101;
#1 $display("%b", po);
# 1  pi=207'b100110001000001111101111101000001011000100110011000011010100001010110011011010110010110010011010000111001011100111101001110100011111011101000101110110000110000010001010110011010100000000110000010001100100000;
#1 $display("%b", po);
# 1  pi=207'b010010000110110100100000011111110111001100010001110100111000101000001001100001101001100100101110000101011100011001001000010101110111011011100000111001000000111111110000100100100110010101111000011101011111010;
#1 $display("%b", po);
# 1  pi=207'b001000000001001001100101110010000010110101011001110000010010101101101001001110111111110001011010001000011101111110101001100011100001111010101011111011101011110011101111110000111011001001000100001001000000110;
#1 $display("%b", po);
# 1  pi=207'b100011100011011100011110011010101110101001101000011110110000101111101001001011110101101100100111010111000101010010011000010101011110100101101101011100000101011100100011001001100111010001011110001011111111001;
#1 $display("%b", po);
# 1  pi=207'b111101111000001110001110110111110110111101011110010010001011010110010010100001010111111111110110111110111001001000111000101011100001011011100010111101000000110100101101001110000111100000011100010101111110100;
#1 $display("%b", po);
# 1  pi=207'b001001010011110000110001101000111011101110101011101001101010110000101100000111010100000110011101101011011000001001010011100001000000010100100111111100101000011111101011010010110110001000011111011111111011010;
#1 $display("%b", po);
# 1  pi=207'b101001001011110100101000101000000010111001111010110111101100001011101101100101111111111000001010001001010101000111110111000010101101010001000000010111100111001100110101010010000000001011110111101101100011110;
#1 $display("%b", po);
# 1  pi=207'b011000001001101101111011101001110010101110110010010011111001011010101101111001101110000110011110010100010110000110110001010111100101101011000110001110100100001100001010001011010100100100101111001100001110110;
#1 $display("%b", po);
# 1  pi=207'b001010100101000001101101101101011000100110010111011100010011100000001110101001010100000100111010000010111001001101011100010111001101011100011011011011011101011011011010111001010100010010111101011101110000001;
#1 $display("%b", po);
# 1  pi=207'b100100010010001001110111000111111110110110010001111010000111011110100011111100100111111010011001001010111000010110110010101000100011010110001011011000011100010111110101011011000000000110011100111110111110010;
#1 $display("%b", po);
# 1  pi=207'b000101110001010011011001110011011110000101110010001001110001011100000010000100110110100100011010000100011000001010111001000001101000111001000100000000110101000100011110001011110000010011000100001100010000011;
#1 $display("%b", po);
# 1  pi=207'b111000001010010001000100010101001010011101110101011101100110100000100111001110111000110111101011010011000000110010010101111000011101111110111100111110000110101001100111001001010000111111100111010101110001011;
#1 $display("%b", po);
# 1  pi=207'b100101100101111100011000101100111111101110111100100001001000001101000100100011110100100111101100010110010111001101001110100010000010101110011011011101000011110110010011110100110001100100111110001111110010111;
#1 $display("%b", po);
# 1  pi=207'b100001001011001111011011010000010100001101100101110000101110011111001111011000010111110110110101110001010011100100110100000001101011001000010101111100011011000111010010101001110101001001010010011010010011110;
#1 $display("%b", po);
# 1  pi=207'b000101111101000010000010101111110010110100011001011010010010111101111101111100111000111001011111100101101010111110000011001100001010000110010010111000100011111100100111101100001110101001110010011100111011001;
#1 $display("%b", po);
# 1  pi=207'b001110001011101000001110100101111011001110110110101101111010111010010110111111000011110011100111011100111011001010000001001110100001011000101101001010101001010010000010001000110001111011110100111011110101110;
#1 $display("%b", po);
# 1  pi=207'b011010010111001011111110101001011000110000011101110011010011110111111110111001010101010000000001010110001011101110011011101010111111100101010101000100001001100001110111101000001010010011010110111000100010110;
#1 $display("%b", po);
# 1  pi=207'b000011010100111001101110111011110001011111100100011100001101000111000101111011100111111000101001110011111111101101111001110001101010000101111010111110010100011011101010101111011000011000110001011110000010010;
#1 $display("%b", po);
# 1  pi=207'b011101110011100101110101111010101000100001011100010010000100101110111101010011010100011110101011010011000000011111011101111100100001111010001100101100001100101011110011111110110101000000000010001111110110100;
#1 $display("%b", po);
# 1  pi=207'b111011110000000000111001101001111111111111011011000001000001000111001011001110111010011101101101100000000101111011000111001100110111010101110000110010101001100110100000111011100100110110010100110101001010011;
#1 $display("%b", po);
# 1  pi=207'b110100001011001101101110101011001110001111001101011010111110110010110100011100001010001111100100010111100010101001101111010100010001001000101101001101001101011011101111011000001011110111100111011000010111111;
#1 $display("%b", po);
# 1  pi=207'b000110001000100001011011001010100000001010100000010010000000111000010000011101011000111110101001011100100001100110011110010001111001110110111010101110010011000010101001111011111011010011111111011011111001010;
#1 $display("%b", po);
# 1  pi=207'b101001101000111101001111010111000101101110101110110101111010010100111011100111011010100101100011000111100000010000101100001100111000010111011001001100111001100110111010000000110010010101101011000100001001010;
#1 $display("%b", po);
# 1  pi=207'b001101111101101101101011111011001111101011100110011010101011101110111110001110101100001000110101010111111011001101110010010101111001111100010110101100100100111111000100101111001001010100010010000110000000000;
#1 $display("%b", po);
# 1  pi=207'b000011100010110001101111110011110001111111001010000001110110101000011011010001111000100010011000101110011111010100110101001111101001010001011110001100100000000110001110010000110001110110010101100111011000100;
#1 $display("%b", po);
# 1  pi=207'b111000110100100000011101100000011110001010010011010011001001001001000010110011111011010101110001010011010100100011111100111001110110101111100111111011011011110011101100101011011110011101000000101000111001000;
#1 $display("%b", po);
# 1  pi=207'b011111101011011001000110110000000000001000000010000010000010111101010001101111010110011000011101001110001101100100011001111110011001101001001100001001110001111011111000101000000110110110010011000001001101111;
#1 $display("%b", po);
# 1  pi=207'b100000001010001000010000111010110100111101011100111101101000000010111011100010000001011001010000001011011010011011001011111110111000100000001010001001101010000100110110001100110011111001101110011000111100110;
#1 $display("%b", po);
# 1  pi=207'b000011111111011110010101000100001100001001011110010110010001101000110101111101000110111111111011101100000100010010010101110010011011001100000000101011101011001001110010000110100000010100011011001110100000111;
#1 $display("%b", po);
# 1  pi=207'b100111111001000100110000111010110010000110111100100100011110101000001100101111011110001101101100110001000100011010011001100101001111101110011111111000011010001001101101100000100101111111100111011001100110000;
#1 $display("%b", po);
# 1  pi=207'b001100010010011110101100110000000000011101001110001001010110000001100111111110000011011101000011101000010011011011011100101010010111110111111000011001110011010101011001110111100100101101011101000101010001001;
#1 $display("%b", po);
# 1  pi=207'b001001101101101110010001001111010011101111000100111110000000110010100011010100100011010110111001010010000000000111011000010100011011100100000010000001111011100100111101100011111100001001101111000010000000010;
#1 $display("%b", po);
# 1  pi=207'b100101011110011011000011111000001011001111100000111000100111010111010000111010001000011011011000101100000011001001100001001111110010111101111010111110001001011010111010001111010010100100001101111011100001000;
#1 $display("%b", po);
# 1  pi=207'b001000010101011110110011011100010001010011111101101000010000000001001100000000111011011101000001001110101000111010000001010101001000011011111101000111011101101011101100011101100110000000011101001100011001100;
#1 $display("%b", po);
# 1  pi=207'b101100000111110101111101000011010110111000011010001111101011110100101101100001000110101001111101010110111100111001010011100011100001101110111111110001011110011111101000011001010110111111101110000110000011111;
#1 $display("%b", po);
# 1  pi=207'b000001011011001101011101010000011101100100110100011010000110110111010111010011011011011000001010010011001011100001100000011110000101010000010001000110110100101001100000110111001001101111001111110101001111110;
#1 $display("%b", po);
# 1  pi=207'b010111010100110100101101111000010111001000000000101011000111001110000010100111110000111000011011011011101110000110001010011101111110111101011011101101110000111100101111000100101101111000100011110110001100010;
#1 $display("%b", po);
# 1  pi=207'b010010111101101110110011111000000010011001111000110110000110110101110110111000100110100011100111101001111011010101100101001111000011100011111111001110100100111101000101001100101000110011101111110110101011101;
#1 $display("%b", po);
# 1  pi=207'b110101100100001001000101111100011101101110101001100101101010000110101101000111110111001001111000011101011001001011110101010101001011101011000110001011010000110110000100100010101010100011100000110110000110000;
#1 $display("%b", po);
# 1  pi=207'b001100011011101011000000110110010110100110110101101100011100001110001110010101100101011010101100100110111110011111100001110010010000100010100000000110111000100110011111100010101111101100000101010101010100011;
#1 $display("%b", po);
# 1  pi=207'b101000010011111101101010011101001010100011000010000111111001110000100001000001101111010100101011000110111100000111000101101111000111111010110110000100001010001001101100011110100000011001010100101001000110010;
#1 $display("%b", po);
# 1  pi=207'b000010001101101110011010110011100010001111110111100011001011110000111100001011000101011001001101110000000101010100011101000010100101100010010110110101011010111001100111010110110000101011000111101011000101011;
#1 $display("%b", po);
# 1  pi=207'b111101101001101001101000100100111000011101001111011101111010110011001001100000101101010010000110000010101101101000010000100110011100110100110110100110100100110011110100101010001111100100001111001011011100111;
#1 $display("%b", po);
# 1  pi=207'b100100001011000100101111111101101010110110101101111110010010100011100001111111100101010110011100000100010111100100001110111100110011101100100110100000000011011010111100001011100010110010101000011010101011010;
#1 $display("%b", po);
# 1  pi=207'b000110101001011010011100110111011111000000011100100010000101110101111011000000100110011110011110000010001010001011000100000000101001100000001100000010011101001101100011001111000101001101101101111010110010111;
#1 $display("%b", po);
# 1  pi=207'b111111101001110110000010010100000110111001010011111100000010000011001111111001001100110111000011111011001100100111101011100011100100011101001011011111001111000011000101101001100001100000011110001001100011011;
#1 $display("%b", po);
# 1  pi=207'b110111101101011000111101110101010100010000011100100101110001011110101011011001001101001110111010111111000011010100001010010110110110000110101001000000111000011001111110010110111100111111101000001110010100101;
#1 $display("%b", po);
# 1  pi=207'b001101110100110001111011000010101011101000111001100010010011010000011110001000011010001101100100111000111011101000001101001001111000011010111110010111110110111000110111110000010011010011011100101001100011100;
#1 $display("%b", po);
# 1  pi=207'b000000111000011101111100111110111011110110101011010110111000101010011101110101011100110111110110011101000011110111110110010110111110101011010001001001010011100001111101001001110000110010110100100010101010101;
#1 $display("%b", po);
# 1  pi=207'b011101011011001110111101011010101001000011001000011000001010100111100011010101101100011001100101111000111011110110110111011100100010010000011000000101011101011010111111100110000011001110010000011001101100010;
#1 $display("%b", po);
# 1  pi=207'b001110011111101110000100000000101001110001011101001100010010010111101110110111100111111111001100100010001100110100000000001010100101100000000011111011101100010110100100001011111000010111101000010001110110010;
#1 $display("%b", po);
# 1  pi=207'b110110111111011000111100100011110000101111111101011010101100110011100011101100001010011001110001010001100001010010101011101111110110010111001000011101101000100011111110001101100101111111011011100100101110001;
#1 $display("%b", po);
# 1  pi=207'b011101110101010100111101000100101101101101010000111101010100001010010110111000111110011011010011111010011101100111100110010011000011010011001001000000001011111000000000111110110110100001000110010110001001110;
#1 $display("%b", po);
# 1  pi=207'b101010101110100110001001010000010000101101000001001100010101001101010001101000101100010110111110001110011100001000001100110100101001000101000110011100111101001001111000010011000111000000010100110001111101101;
#1 $display("%b", po);
# 1  pi=207'b110011101011110011010000001110011111001101101101110010110011101101011101010101110110110111000011110001101000100011011011100110110100100011000000001011110000001101110110011000111000100100111100110100011110110;
#1 $display("%b", po);
# 1  pi=207'b011100000011001101000010110100000010001100001110011111000010101011110011111011111110100001010101100111001110100110010101101101101101010010011011101011100010011110111101001100001110101101010100001110010000010;
#1 $display("%b", po);
# 1  pi=207'b111101011001010010010010101110011111101110000000001001100101110010110000110100110110101001000101100000100100010110100001001000101000111011010101100001111010010101011000110101011010010101101001010111111000010;
#1 $display("%b", po);
# 1  pi=207'b001101100001100100011100101111100000010100011100001010010101101000001011100101100000011010101001010110101001001110110000111011100010101101101111101111001111111101011110001011101111001000011100101010110110101;
#1 $display("%b", po);
# 1  pi=207'b010101110111111100100111000111001000010100101000110000101111100010100000110110111010000101101111111001011100011101100011101011010100000110101000100011011011101101001001000001001010010100010110010110111100101;
#1 $display("%b", po);
# 1  pi=207'b111101011100110100111110001010010100100010001000110101010111000001000110111011101100110010101011000000100001001010000101001100001001111101011010000101111001011100011111100001110111110010101100000111110111010;
#1 $display("%b", po);
# 1  pi=207'b001110111110011001110000000010101110110000100011111010101101101001101111011101101111010111000010000100110010111111110111010110000000111111010100101110010111101011101010011010010000000101011110101000111101101;
#1 $display("%b", po);
# 1  pi=207'b111111110111011000111001000001011111100100000111100110010010101110110110011011101000111001110011011000111110000100100111010100110101101100101100011011011010110101001111011000100101001010100110111011111111010;
#1 $display("%b", po);
# 1  pi=207'b111101100000110010110001001000111001011101111100000001010011001010000001000010000000110101110111010010100101100000111111000101010010000000110011001101101111001110110100110000010000000011101111001000101011000;
#1 $display("%b", po);
# 1  pi=207'b100110001110011000110001101101011101100110010101010110101010111110010110000111011011101110110100011110011001000001001101101101100111101010010101010111101111011101001011010001010101001101101100111000000100111;
#1 $display("%b", po);
# 1  pi=207'b000011001111010001010011010000101001100010110001010010110101110101010011101011001101011010001101100110110000010001000011110001111001011010100011001011001001011011110010101110100111010101011011101101110001110;
#1 $display("%b", po);
# 1  pi=207'b101100011101101000000001100001111001011000111101101000111101010100001011100111001100100110010010110001010010011100000101110000110000000001100000100101000101001110001011110000001110100010011010010001011000110;
#1 $display("%b", po);
# 1  pi=207'b100001100010011100111100111110011110011111100011001110101101010000111110001011001111111000010110101001110011100001010110100101101011111001000111111100100101100011001001010000110101100100100100001001000000000;
#1 $display("%b", po);
# 1  pi=207'b000110001001110010111110101110100001101110011001010111111110011111001100111101001100010010110011011000110111011111010110011101010010000001101000101001110000111101011001101011001001010110001001001010101001110;
#1 $display("%b", po);
# 1  pi=207'b010000101110111000111010010001101100101010000110101001110110110101011010100011001001000100110011011110000101110000000110011010010000111011000111101100011010010100101011101111110110011101000110101101011100000;
#1 $display("%b", po);
# 1  pi=207'b010000010001111110111101110111110100000101011110100001100000101011011001011011101101101011101010000010001110111000110010111000100111001111100110101001111110110000011100011111001101000001100100000011011111000;
#1 $display("%b", po);
# 1  pi=207'b001110010101100111101101010010110110011110101010100000111110011100000011010010011000110001101100111000001111100100011111111110101010111011011111100101000110011110011000111001110110010001010101101001011100100;
#1 $display("%b", po);
# 1  pi=207'b001001100011101000011100000000011000000101001001111000000011100001000100000000011000010010010001111000101010101001111010111000000011100000001000010101001111110101011001000000001100010110110000100101000010000;
#1 $display("%b", po);
# 1  pi=207'b000000101001111111000010001100001001101011101100111101001111010000111011100001101000100111011101001000111100010000011111111001000011010011110111001011110000100110100010001001001111101010011101011000000101000;
#1 $display("%b", po);
# 1  pi=207'b100001001001000010000101000100001111000111101001010001000000000011000001010000101110001001101000111010111001111010101111100001001011010000101011011101101000100010011101100011110101100100011100101101111001100;
#1 $display("%b", po);
# 1  pi=207'b110001010011000000111110100100010010111001000110010111101100011110110000000100010111010010010110011100111101101111111000100110101110000110110101111110000111010011111101110111000101111110100100110011000110101;
#1 $display("%b", po);
# 1  pi=207'b110000111000011001111001110001000101010111111100010101110101001010001111100111111111111010110110101100010101101000001101101100101001011000001110110011101111010010011001100011010011100001101111101011110100011;
#1 $display("%b", po);
# 1  pi=207'b000000010000000001000110011011011110010000010000010000010111111110011100000010100001010000000010010011101001000110111111010101101110010100101010011110000110011010111011010000001110010010010011110101110001000;
#1 $display("%b", po);
# 1  pi=207'b101010011111100000111110111011100000101010010111010101101101110100011110010111001010101110011001100101011010000011111001101000111101011101010110110011010111101111010000110000100010111010111101101011100100000;
#1 $display("%b", po);
# 1  pi=207'b110100000011110000001000001011001010011011001010110001100011110101010000110110100101110000000011111010110110100011011111010101101010110011110110001010001010100101000011110011000110011010110011101001100111111;
#1 $display("%b", po);
# 1  pi=207'b011110111101000011001100111111011010011010110010011110111001001101001001010001100010001000001100000101011000110111101011110010010111000111011100010010001000000111100101010011010111010000110010000000101101111;
#1 $display("%b", po);
# 1  pi=207'b110000101010111101100101100011110100111000000000111101001000000001101110010100000110011111010100111011010101000111000000011011011010110010011101101101111110011111111110001101001100100100110011111000100110110;
#1 $display("%b", po);
# 1  pi=207'b110000011001001000000101101001101011001011101110110011111111111001011001100100001001011101110110010011010101101011100000100000000110101010010001010001110001000110010100001100011101110000000001000000010101001;
#1 $display("%b", po);
# 1  pi=207'b011010110001011111011011110100010100100100000101011100011101011001101111110000001000011011010010101110100011101010100101001111111110101110011010110111000001111010000010000101101100101110100110001111101111100;
#1 $display("%b", po);
# 1  pi=207'b111010000100011100011010001111111110100011101001101010111000100100110001100001011110011011100011111011011001100100000001100010110001111000011110110111101111010110101001010101101001011100011010011111110010011;
#1 $display("%b", po);
# 1  pi=207'b111010001011111010111100011111000000110000101111101011101110011101101001011100110011101111000110001110010010110101100101101110001001001101110100010011011110010011000001010110100110000011100010100000111010011;
#1 $display("%b", po);
# 1  pi=207'b001011010010100001100010010100000000110111110100010100111010101011111100111111101111111101001010011000100010111111010001001101011011010010101100101110010000001001000111100001111101110010001100100110010101111;
#1 $display("%b", po);
# 1  pi=207'b001100100011100010001010111001101010101111101100101110000100101011100100101100001100000101100010011100100010010001101100110010011000110001111110011100111110011001100000000011001110000100101000111010101010101;
#1 $display("%b", po);
# 1  pi=207'b000010110011101110010011001111010000100011001001011110000100001011000011011100110100010000011001010111010010101011010000111101000011000010011101101011110110111011001011001000010110001011011011001110011100000;
#1 $display("%b", po);
# 1  pi=207'b001010101011111010111100000111011111001010100001010101101100111101101111000010111101010101010010100001100000101011011001000000110000100001000001110101000101011110100001000000010101100011001110110111000100101;
#1 $display("%b", po);
# 1  pi=207'b100111100111010100101111101100000111100000111110001100010101010100011101111101101101111000100001110010110010101111101100111010000110100101100011100010010110110111100010110101011011100101000111110011100101110;
#1 $display("%b", po);
# 1  pi=207'b101110111110010101100111111011100110110011111101010101000101011010101011110000000011000001010111101010101100100011010001111010011011010010000011011101101000111110100111001010011100011011011001010110101001010;
#1 $display("%b", po);
# 1  pi=207'b110011101101011000011111110111010101111101010110110011100100110110100110101111111001100001000110001011111010011100111000111110100110001110000001001001001010011010100000001000101001111010011111100010111111101;
#1 $display("%b", po);
# 1  pi=207'b111010011000100110100101011010111000010100001001100110100011110101110110011111010011100111010111011110010010000001110100110101011110110011100111111000100000101100010110111010111010111001101001100111000100001;
#1 $display("%b", po);
# 1  pi=207'b111000100000000010110010100011101001011010010010000110110101101001011001001100000010110110111100011110111101011100011111110010111110110110111101010010010010101110111000010010011001011011001010010101001010000;
#1 $display("%b", po);
# 1  pi=207'b111110100111100000011101010101010000011010000101111100111101000100011101011001000010111110001111000100101010101100001100110010001100001101000000101110000101001001101110011110110011101110110111001101100000000;
#1 $display("%b", po);
# 1  pi=207'b111101110111101100010001000001001100011000010011000101110110110000000011100001111000011101101101010111111001101010111010110010100001000110101011011010000010101011000011010010011001011101010010110010000011110;
#1 $display("%b", po);
# 1  pi=207'b101000111100100001111100100111001001110110000010000010110111110101011101100000101110000001000011111010100010000110110011010000110111001001010100110000000100111010100111110101000000010010101100011110110111011;
#1 $display("%b", po);
# 1  pi=207'b111001000111101101000001111100001001101000100100011100010010100100111000000001111100000001001110010001101101010001001011011000010111000010111010111011001110111010101010101011001110101000000000100011000111010;
#1 $display("%b", po);
# 1  pi=207'b100101000101101101001001011011111001110100101100011101011110101001110101011001000101101101001111101111001011000111100111010101011110000100011100010111010111111101100000010111101011000100100010110010100110001;
#1 $display("%b", po);
# 1  pi=207'b111100101000101010000011000101110010111001000000100000110011010001111101000101100011110100110101101111011101010101001011000100100101010001011110111111101001011010110111111110011100101100110110011011010011100;
#1 $display("%b", po);
# 1  pi=207'b001011001011100110000001011001010011011011011000011011011111100000001000101111001010100010010010101101111110110100000000010011100111111111011011000011110000101010000101101110111000011000000101000000011010001;
#1 $display("%b", po);
# 1  pi=207'b001010010010111000111111110110011100011001000111101100110111110100001001001001100100101101000100111110000010011110111011010101110011101001000101100101110111000010110010110110000001001101100011100110000010110;
#1 $display("%b", po);
# 1  pi=207'b111001010010100100110100111001001110101011000100101110000000110011100100011100000101000001010010011101101001001011111100001100100000101000011100000111101111000001101100110000101001010101110111110011110011000;
#1 $display("%b", po);
# 1  pi=207'b101110010101011001101000000100101010001110011110001100011110010011011011100100111100010111011111110101001100101111001011010111001100100101100010110111010101011001001110001110100011000000011010001001110000101;
#1 $display("%b", po);
# 1  pi=207'b000000011110001101011001100001011000010011100000001010001101111101010011011110010001101011001110100111100110010010100101010010110001111111110100010101110001110010000100001100110100110110010000101110011110101;
#1 $display("%b", po);
# 1  pi=207'b000110010110011011110010100011101011111111001010111001111001100000011101110100000000001010000110111011001100100101111001110111100101111010011010111001100101110000101101000110111010000110010101110011110110010;
#1 $display("%b", po);
# 1  pi=207'b101011001011110101001001001001111111100001000010001001010000000010010000001010011110011001000000011011110011010111111100110000011101111100001101011101010100100010010100011000111100010011100000111110001010000;
#1 $display("%b", po);
# 1  pi=207'b100100111111001110001001110110111000101111100101110000100000100111000101110000000001111000011001001111111011100000110001101001001010010101110111010111111000001110010011110110100100000111111011001111000100001;
#1 $display("%b", po);
# 1  pi=207'b111001011100111010010010110011010010001010001011101001100001011101001000110001010111010100111000011010010001101000001011111101000111000010000000001100101011011010110110110011101011110000000000110100011001000;
#1 $display("%b", po);
# 1  pi=207'b011001011111001100011010000100100101000111010011110100101111111010010000011001100001101011010001100001100110001111000110110100010111001111010110000111101110001101000100110110011010110001011011110100100010011;
#1 $display("%b", po);
# 1  pi=207'b011000010111010111011010100001000100111111011100011100100011111011101110100101011010000001100001111001111110100101101101101111111101011101010111101111011101010011010010001010000110101110101000111000000101101;
#1 $display("%b", po);
# 1  pi=207'b110110011110100010000111111010111010100001110100101001011010111011000011110100001001111100010100101011001111100000100000110001110100111010110101101101011101100111000011010001100101011010110100101100111001111;
#1 $display("%b", po);
# 1  pi=207'b100100001111001110011000011101011001110010011101110000011111000010000010110001001001011111010111101000101110001001000010000011000000011110011011100111010001101010001101001110110100100100110000111100010101010;
#1 $display("%b", po);
# 1  pi=207'b011101110101111110011111101000100001100010000000001111010010100001000000011001011111111100100010011010111001100110111111010011000100010011001001001000011010111101010100001101000011000000111101000111110001001;
#1 $display("%b", po);
# 1  pi=207'b001100100100000001110100010011011010101011001000000111111100011001010101000101010011111110111110100100000111101100000101000000001111110110001000001101100101001111001000010001100001011101100100010011010010101;
#1 $display("%b", po);
# 1  pi=207'b101111011010110110100101000010111000001011110110010111000110011110100000101000001001110001011011111100011110001001100111110001110001010011010010001010111000011000100111010110110000000110101001010001101001000;
#1 $display("%b", po);
# 1  pi=207'b010001000001100100010010110000101110101111011011010111100000101000101111110010100010000000011000100101000001011100010110110010110011100111000011100000101110000000110001111101101110000111100000101110101101101;
#1 $display("%b", po);
# 1  pi=207'b000110000000100000110111010011101000011101000001110011011110001000101011000010011000111010001011000111111001011000010100011101100111000100010000010111110101111110110010011101101110111110000101001000011101010;
#1 $display("%b", po);
# 1  pi=207'b000111111010010101100010011101101010111110110101101100011011101111101000110100001011101101001010010100110100111000101000001010111010100100001101011101110100100110111000101101000100011101010000010111011010001;
#1 $display("%b", po);
# 1  pi=207'b000011110111010100011101011011101001110001111001101000010011111111100110011100000110010111000100011011100101111011011101101010101011110001000101011111110101000000110001010000001011100101110101011011100110110;
#1 $display("%b", po);
# 1  pi=207'b011111011011111110100010110101011010010101010101101001111101001101000100010001000000010010010000011010100011101011000110000001110101001100011000011010110101111001110101101000110001000011111110011011011100101;
#1 $display("%b", po);
# 1  pi=207'b111001010110100011101011011110010011001000101110100100110111011100101111110001000001011100011110000000010001001011010001000010111001100101110101001110000010011011011011001010111111110010000010001111100011000;
#1 $display("%b", po);
# 1  pi=207'b101000100100111101010110111101111111111010101100101001110000111101110000110000111001000010011011011011000010000100111010011110101010010110100010111000011110011000101001001100000110011010011000101111001010111;
#1 $display("%b", po);
# 1  pi=207'b011000111011100101011011100110001110111000001011011110101110010001101110000101100001111101100110100010111110010110100010101010101111111110111100010100111110101100111111110111101101100100111111111011000011101;
#1 $display("%b", po);
# 1  pi=207'b010100000111011010001110010011100100001000110101011011011000101010111110001001001101011101100110101010010000011010011111100001000110111000000011110101101000000010000010001000000010110010010000101100011110101;
#1 $display("%b", po);
# 1  pi=207'b111000010010111001100110100000000111000011001101110001010110101101101110001011001011100010000100010011111111010010111011100000001101001110010111000110010010101111111000100110101101000111001010100101110110101;
#1 $display("%b", po);
# 1  pi=207'b110110101000110010101111001010010111100101110001111001110010101110101100101001111000000011110000011110101111011111001111001111011001011111110111010100110111101110000001010000001000111111001110010101101001010;
#1 $display("%b", po);
# 1  pi=207'b110100010001110010111101000011011110110000010111000011000101011011111000110100110010001111111001011110100101110110100110001110001010100110101011110001100111001101010010001001110101111000010010001010110110101;
#1 $display("%b", po);
# 1  pi=207'b110100010000011010000010100101111100011000001111000000011100111111110000010110010011100010000010111110010100111101000101100100110110111010010101101101110000010011000001000111000110011001111111011011101101101;
#1 $display("%b", po);
# 1  pi=207'b001101000101111101111111011101110010010000101110001110101001010000110101100111111111011111000111110101111111111101110111110010010011001111110111001001001111010000001001000101010011101000011000000111000111100;
#1 $display("%b", po);
# 1  pi=207'b100110000010111001010000110011111010001001100100101111111101101010000001100110001100100101001011000111010010010011110100011101010110000101011011100000111011100101000000110101100011010111001101000100100001110;
#1 $display("%b", po);
# 1  pi=207'b100100000101011000010010101100111111101011010001010011000101001111101110100001110000101001010010011111111010001001101011110111000101001001100011110001100110110101100010011001011101011101011101110110010100110;
#1 $display("%b", po);
# 1  pi=207'b101110111110001111110110100101100000000110001001101111100000010011010011111111111001011001110011110101101000001111001011001101111111010001101001010011010100101011100100111111011100110101011100111100100110010;
#1 $display("%b", po);
# 1  pi=207'b111010001011100000011111111100000100001001011100011000010111011010001011101001010101111111111111111001100010010000110101111001011011011101111100100011101111111001000100110110001010001111111101100100010111111;
#1 $display("%b", po);
# 1  pi=207'b111100000100001000000111111011101110110101100110000011001111011001010110100011101100011010010010100100010110111001101101110010001100101111110000100111001111000111000010011000101100000010011100000010111111010;
#1 $display("%b", po);
# 1  pi=207'b010111110110011100111101011001000010010100111111010110011001101110101001110111111101011010100100111010110100100110001100001001111011000000000011011110100001100000010111100001101110110100101011000101001011110;
#1 $display("%b", po);
# 1  pi=207'b000011100111010000101001101110011110101001010110001011110100110100000110011000110011000101101111000010010101111000110110100000000001000010010010110111000101000000010101000001100111011010100110100011011011010;
#1 $display("%b", po);
# 1  pi=207'b010011010110111000100011001000010011000111101101000110000001011101000110110010001010010001011010110110100110110010000100010110000011010010110001010010001110100011100101100111000001001111010100111110000100010;
#1 $display("%b", po);
# 1  pi=207'b011001010010110111110111011110111111010111010100001000001001011011010001101111111101001101100011110000011000111011010001000010100110010101101110101111001101101110111100000101001011110110011100000100101000010;
#1 $display("%b", po);
# 1  pi=207'b011101010011011101011111110111001001100000101101101100111100111010010000000010110111100101011010111111001001001100010011010011011100011010100111011011001110010110000000010101110101011001100111110101000010001;
#1 $display("%b", po);
# 1  pi=207'b101001010010010110111000000010011100000110110001101110101110000111010101001101111101011000010010110110010011100111111111011100000110001100000110011010101010110111011100101011000100101000110011000010001110011;
#1 $display("%b", po);
# 1  pi=207'b100100011100111111110111000010011011110100110000110001110011000100111101100111101001000000000001101101000110110011000011100000000100111110111101111111111100111001010000111111001001101001110110101000101110100;
#1 $display("%b", po);
# 1  pi=207'b111100111100000101000110100101011101101000111010100001000100011111011100110111010110110011110100110111100110001101001000111010010001100111100111101111100110100111101110001011000010111110101000101101001000101;
#1 $display("%b", po);
# 1  pi=207'b010011001010100011111001101011110111001001111100100111001101011001001010101011110011011101001101111101111111000110011101001000101100110100010001110011000011111110011111001001011100010000011001010111011010000;
#1 $display("%b", po);
# 1  pi=207'b011001000011110010111111001110011010100110001000000110011011001101000100110000100000010111011111011100011100101001101111111011100101110110111111110010100110001011010100010101101001100111000111101000101000111;
#1 $display("%b", po);
# 1  pi=207'b000000101101000010001100010011001101100101111000101100100100101000010111111101110011001110101001011110100111001110010011100010011000101000000000010111110101001010111110101110100111100100001111101010111100100;
#1 $display("%b", po);
# 1  pi=207'b111101111101101001001110000110001101010001001000010110101001011001000110010100101011110001000001010111001011111101101000000111011011110011010011101011000101010111001010101111010001100111111110000000101010110;
#1 $display("%b", po);
# 1  pi=207'b111111111111111001010001110110011011001000101010010010111100011010011101011010110001001101011110110001110011001101001101101001101001000101110010000010100111001110111000100111010000010000001101101000111011110;
#1 $display("%b", po);
# 1  pi=207'b110001101001101111111000100010101100110111010100101011101000100101100011010000010010000010111101000111111100011011010000100101010001111100100011010010010011010010110011011101000001011101011101111000101011011;
#1 $display("%b", po);
# 1  pi=207'b110101111000011000101110100100001111001011100000000000011111110101011100010000001100100111100101010010101100011011111010011000000011000011111101010110001001110011111100000101101000000110000100001011110000110;
#1 $display("%b", po);
# 1  pi=207'b100100011011101011001001100111011001010000001101001110010111111001101011011111001101001111000001111001010100011010101001111100000101100101100000101001011111000000001110010111100101000001001000000110001000001;
#1 $display("%b", po);
# 1  pi=207'b110001000111111111101101101011100011000110011001111110011100000010011101101001110001110111111110101110001101001000001001101001010000111000010111011000100110111011000100111111011000001000111111000000110110000;
#1 $display("%b", po);
# 1  pi=207'b111010000010000011101101110100011100010100111110010100001001001011010101001001110010011011111101010010111111101011110110010001011011001001010010100000110110011010100110101001010010110110001111000111100010011;
#1 $display("%b", po);
# 1  pi=207'b010100001111011010010011001110011110111010101011100111100101000101100001011000001010101101011011001010011010110001111001001011110000000010011101001100001110001010101100011111001000101101100001011001100111001;
#1 $display("%b", po);
# 1  pi=207'b111011100111110100100111000110001100001011001011111000101001100101001110001011101111111011110101000011010111010010000011111010100000011000100000000101000000100010010001110110011110101111011011110111110011101;
#1 $display("%b", po);
# 1  pi=207'b011011111010101010000010101111101110110110010001110000110110101001001101100000101000111011010111000100011100111000000101010111000110000100100000101110010001101011010101011001010111000111000101010000100110001;
#1 $display("%b", po);
# 1  pi=207'b000100100100001000101011111000011010010100010100101001110100110001011101111000111110111110011010111001100010101101010111110010001100110110011010110001111000111100110000001000100001001110111010010111111111101;
#1 $display("%b", po);
# 1  pi=207'b011110001101111110101111000000110100011000001111010110011100101111110110111101000111011101110000101000001001100011000111101001000110001001011001101110101110111110000010011110000001110101111101001001010100011;
#1 $display("%b", po);
# 1  pi=207'b001110001100011100011101011010110000010110111111110100101110110011000001101010000001011000111000011111011001010111110110111011110001011010000010101111011110110011000000111010011110111001110011011110100000101;
#1 $display("%b", po);
# 1  pi=207'b101111010111001100110100001111001100101000100110110010100000100011100010011100100010010010111011100011101101110111011111111010100011000111010110111111010001101010011011010101010110010100011101111111110000011;
#1 $display("%b", po);
# 1  pi=207'b110001101001101000100110111111010111001100100000100011010001101001010010111011101101011010100111010110011111110011111000000101101010101011001001101000010000001011100000011110110111000001110111111010101100101;
#1 $display("%b", po);
# 1  pi=207'b000101011100011000001101100011110101011100000011000101000111001101100100101100101011100011001010001011011100011001010010000101000111001101100001011001110100110111100111010101000000110000101111100001101100100;
#1 $display("%b", po);
# 1  pi=207'b011110111001110000111111011010100100110001101101110100001100100010110111001101101111010011100000100010011111101111111100001111101010011000101110101001000111111111001100000110111101111110011100011101110010010;
#1 $display("%b", po);
# 1  pi=207'b011100110111000010110101111000110001101010111100000100001010111101000110001001101110100000000011111100110100001100110000110110101010011111100111000000010010010010111011010000111111101101100001001101111101010;
#1 $display("%b", po);
# 1  pi=207'b011011011011101011110010101100000111001101111010111101111011001010111010111100001011110001100010000100010110001001100101000111101101010010000000111001101101110000111110010100001001010110101010110001010110101;
#1 $display("%b", po);
# 1  pi=207'b000101100000001110011101011010011111110111111010101001101110001111111001100010100100110000111011100010110000110110010001101110100111101011011101101010000110101010101101000010111110111110110011111101110110001;
#1 $display("%b", po);
# 1  pi=207'b000100001100100110100011000010010011001010100110001110100001100001101100011101010000010101011011000101100010001101001000110000000111010011110110000111111100111101111101001001110101111000000101000111011011011;
#1 $display("%b", po);
# 1  pi=207'b111000100110010101000011110010111001011100001100001111001100010100000000000111110111101001111100101101010110010111011101101111000001101101000001100011000001011011001110001011010111001001000110111001011111011;
#1 $display("%b", po);
# 1  pi=207'b000011011000111110100110000100000010100111000011001100001101110100101011000101000111101011100111100111000011101110000001000101011010011010001011001010111000111001111010100100100100111100101100000100110101111;
#1 $display("%b", po);
# 1  pi=207'b000010001110001011111011110100100100101010101100110111100010010000001010011001110010001110111101100001110001100110000000101101111100011111011010101010000000101010111100101101001010000011111100011111110000110;
#1 $display("%b", po);
# 1  pi=207'b101010001101010000000100001111110110011011010011100010110001101000100110110101111001010001101111010010101111101110111001101011010001000000110111011100111101001101101010010111000010100001011011110011010111111;
#1 $display("%b", po);
# 1  pi=207'b011010001111011010001101010101010111100001010101010110000111000001100100100100011100110110010110100001010111010000011100001111111101011010000001000110000101110111100010111101100111010000100001001100000011100;
#1 $display("%b", po);
# 1  pi=207'b000111010110111111100001000101011111110111000000110101100111101000010011011011101010011011100101001010001101011000011001101010011101010011100011100100001010011010101011101101101010110101011110010001000101001;
#1 $display("%b", po);
# 1  pi=207'b110100100001101111000000100001111001011010101110110001101101100101101100110001010111011000100100001110000000110111111110001100100000100111111100000110011000100101011010001110101010001101011101000001111011001;
#1 $display("%b", po);
# 1  pi=207'b110101001101000011001100011101110011011010011000011100001110000100110000101101101011000100101111010010001100010110000111111011001111100110100010011110000110111000010010000110110101101111111101011101000001111;
#1 $display("%b", po);
# 1  pi=207'b000011000101011011100011111101101111100001001000110100001101000101001110000101011100101100011001000010010111101111011100000010011100001101000110001001101011011010000110101110100010000101100111110110100011011;
#1 $display("%b", po);
# 1  pi=207'b010100011111101000000011100110110101110111011000110110011101001101000110111010111010111101101001010011110000011111001001001011011010111011010001110100011110100110000101000100100111100101000101110110010111110;
#1 $display("%b", po);
# 1  pi=207'b000001110110110101100001100111010001111010001100101100111101010000110101110000100110010111000000000101000111000100101010010100101111010010010001110111001011100010111111000001000010100011010111000100001101010;
#1 $display("%b", po);
# 1  pi=207'b011010111000001111011111111000010101101011000101011110001110111110010110000000111010110000010101100101011001100010011100111101101000100000010111000000100110100001011000000101100011000100111100010100100011100;
#1 $display("%b", po);
# 1  pi=207'b100001101100101111100000001001001101000001110001010100001101110010101011010101000111011000111010011100001100100011110101110000100111001100011111010011011111011110000100101110101001111010011011111011100011100;
#1 $display("%b", po);
# 1  pi=207'b011001101110011110101000111001100101100011111011011011001011011101000100011000100001110001100100010101011011111000001111011011001111110100000000111010001011110001010110011111100101001101111011010110000000111;
#1 $display("%b", po);
# 1  pi=207'b100101001101000000111010111011100100010110110001110001010100010000011111010110001010001011100010000011100110010010111100110101000010000101010000110110010101001111000011010011101011100010010101010110010011100;
#1 $display("%b", po);
# 1  pi=207'b011000010001100110111000100100101010000001001110000011101011101101101011000000111100001000011001011111010000111000011100010010011100101101101001110110101111001001010111101000011010110010011111011101110100011;
#1 $display("%b", po);
# 1  pi=207'b100101110000010001110011111000101110000101001011011001010111101100011010100010111100111101111111101100110100100001000100001100100101100011000111110010001110000011010101010100001001001101101110111101110110000;
#1 $display("%b", po);
# 1  pi=207'b100001000000111000010000010001111010010111111110100000110010101000011110011110001001101110001110000000110010010100111110101010000101111101011111110010010111110111001011110011111011101000011111110100001010110;
#1 $display("%b", po);
# 1  pi=207'b001011001000011011101100001110011011011001101000100001001011111001101010000001100000110000100100001111010110100010111010001110001101101110011011000111100100000110011011100010000100110100011000001010010001001;
#1 $display("%b", po);
# 1  pi=207'b111100000101110110010001010110110011001001100111100000111001101011010101011001111001111011110000000001001001110111000010111101101101101111111001011111111100010011111101110100100101000011100100111011100000011;
#1 $display("%b", po);
# 1  pi=207'b000111101101010011001101000110101011000110111010010100110011000111100000001001010000100000111001110011100001100011001111001110110001001101010011101111101010100111111010010101111001111100010000111110101110011;
#1 $display("%b", po);
# 1  pi=207'b010100001101101001110000000100001110011001010011100101110011001111111001110000010001010010011011101110101100011111110000011111110100101010000101111110111100101010001110000011001010000110001011011110000010111;
#1 $display("%b", po);
# 1  pi=207'b000010001011100011100110011001000101001011010101101011111010100010001011111111000101000111100000011111111101010101000011110101100000100000110100100001000101100101111000110110101111110001011010000111000010101;
#1 $display("%b", po);
# 1  pi=207'b010001101001100001100101100110101111011010000101011110100110001110111000100000011001101000110000010010010011010001101110100111100011101100000101111100000011101001100000111111000011011011110011011111010010011;
#1 $display("%b", po);
# 1  pi=207'b110110010001100011110001000010010100011111110110111011101101100001001011101011000001011000101100110111010101010011010101100100100001111000111100000010000010011000110110110001001001001001000010001111101100001;
#1 $display("%b", po);
# 1  pi=207'b110101000101100001001100000111111001010000110101000100100100001000111000100000100111111011000010010110100011101011101101100010010001001011101011111111011110000110011000000101110011000000100011001110100111111;
#1 $display("%b", po);
# 1  pi=207'b011110011010001110011110110001011011111101011010100001000111101111100010011001111100011100001000101011000110000001100111011000110000010100111111010000011000010100010111100011001001000101100000000000111100100;
#1 $display("%b", po);
# 1  pi=207'b000101110011111100010010111011001011011110110011010010000110110110001010010001001111110110000010101100010011011110110000011001101110111111000110111111100111111011011001010010111110000100110100001111010010001;
#1 $display("%b", po);
# 1  pi=207'b001001111001110010111001110111100000101011111101001011101001010001111000000100010110110001101001000101101000101011011110101110101110011000111000000001000001101000110010110110101010111111111101000111010000101;
#1 $display("%b", po);
# 1  pi=207'b010000001010011110101001110111010011010110111010000100101000100110111100001010001111001111010100001001111000001000011100101010001010011011010010000001110011001110101111010011001101101011111000000010010000100;
#1 $display("%b", po);
# 1  pi=207'b101001100000010011000101001101010111010001000001010110001000111100101110001111010000100001100000100011001101100010101110100100010010000010111000101010100000111101110101110011001000001111010110111111100110101;
#1 $display("%b", po);
# 1  pi=207'b001110111010110101011100111001001100111011111101111110000110100100111111001001000001101101010001001111101000001111001110011111010111011110001101101011001001100101001000101001011110110011010110010100010111101;
#1 $display("%b", po);
# 1  pi=207'b010010000110110101010111010000000110001000110110110010001101110011000001110000101000000101001000010011001110000011000000100001110100101011011011100111110011110010010001001100100111000101000101101000111111100;
#1 $display("%b", po);
# 1  pi=207'b010100101110101110100101001010010111100111100111001000010000110110000000000011101000110101001010010110000110001011101110101111001111000001011110001101110000100100110000110000110001111110001000000101010011100;
#1 $display("%b", po);
# 1  pi=207'b100101110101000010000000010010001000110000001000100001100101011111010101101110000100000110100011100111100111110001110010110111101011100111001100110100100000011101101000101110110100010111110100100000010110010;
#1 $display("%b", po);
# 1  pi=207'b011110100111001011111110101011100111000100100010010001010110110000000001101110110110101001001111001000100100000101011010110011010011111100000011110001011101010001110000010110110100000011110001000001101110001;
#1 $display("%b", po);
# 1  pi=207'b100000101110111110011101001100111110000100000110110110100000111101010000110110000011111110101111011100100011100100000000001000100111011001001010101111000000001011000100010010011101101010010100001101000100000;
#1 $display("%b", po);
# 1  pi=207'b001000110101101100111110001101111100011101001111010010001111000010011010011000010100101000110100001001010111001111110100010010110010010011001101010010011001000011101101011110111001111000010111010010001010000;
#1 $display("%b", po);
# 1  pi=207'b011100001110010100110110110010011010010001101001001110100010101001110001000001011010010100100001000010011010001110110000000101111111001110001000100001001100000110011111001011001011100101100110100110111111011;
#1 $display("%b", po);
# 1  pi=207'b100011101010001010000011001000110110001101010100110111001001010011100110001001111111011100110011100010000001011101101010100000000000011011010001010010100100001010110000000010001110010001010110111011001110111;
#1 $display("%b", po);
# 1  pi=207'b100100000100010110000010001010010100010101100001010101001000100001101000110001001001111010101111100110100001110110011010000101000001111000101101000110010100100110100010001100000001101001110111010010011010100;
#1 $display("%b", po);
# 1  pi=207'b010100011111100001001000101011101111100101100100001000110000100000111111011111010111100000100101001001000101001001110100001010100010110011111000110110101100010110100001000001100101111000001000001001111101000;
#1 $display("%b", po);
# 1  pi=207'b010011010010011110110100100100001000110000011011011001101000001011110111110100110000001001011000000010001000100110100101011010001111110000001111011001011100000101111111001111100100011011111010101101111011111;
#1 $display("%b", po);
# 1  pi=207'b011101110000100010010001100001111100111011010101100011110011111000100000010010100011001001011100000000101010010000011100110111110101011010011101011011010110011100000110101010010111110000010110100000110111111;
#1 $display("%b", po);
# 1  pi=207'b100101011011001100111100110000001110101101110111110011101001111000101010101110100111110011110010010100011011110100101101110110100101001001011001100011011000001011011000101001000000101101011000011100010010011;
#1 $display("%b", po);
# 1  pi=207'b110000000010100110100000010111100000000100011110110010111110110101100010010111100110010001110010001101010010100110100010001100101111011011101110100011000010001010010101011110000111110010100011110000011111000;
#1 $display("%b", po);
# 1  pi=207'b011001111011101101111111010010110101010110100011111000000000111100000111001110010011101010001001010011111011001100111010101101110010100101010001111000010101010110110001110111001011001011011000111101101000111;
#1 $display("%b", po);
# 1  pi=207'b011010110000100000001100101000001111001001100011111011110100011011000100100101001111011110101010111010101101000100010000001111100010010000100100100100011010001001010100001000011010001110101100101001010000101;
#1 $display("%b", po);
# 1  pi=207'b111011111111110001001001011010100111010011000110001100001101100011000111110000100011101010010101111010010001010000011101010010010100100010001000100010111011100101111011100100010010010111100101111111110111100;
#1 $display("%b", po);
# 1  pi=207'b011010001010101011011010101111110001011110010000010010110001111111100000010100010111000000100000110100011110100100100011011101011001011110101110011011010000110101011101000101100100111110010101000110100000110;
#1 $display("%b", po);
# 1  pi=207'b001010001110100100101101110010011100001011011001010101101101001110100101110100011000111101000100001000110000100001111111110111110011110011001000101001111000101010010110001111101010001110101010000001000101100;
#1 $display("%b", po);
# 1  pi=207'b110011010111000010110010001010001110101010011010010010001110000100101101101111010100010010100011001010101111001000111100010111010001011100100011011110001101000010100011011101011000110111101101001100100000111;
#1 $display("%b", po);
# 1  pi=207'b100111101110000001101100111100101111011011010100101011111111000000010011001010010000010011001101001001110001011011110011011110010000001000010010111111111010110011100011010001000111100101010111101011010111001;
#1 $display("%b", po);
# 1  pi=207'b011101110000111000010111100010010010011011011111110100010100100101010110101111010000111111110101010101000111110100011010001100011101010000100011010110000001001011111101010000100001001111010111001111110010111;
#1 $display("%b", po);
# 1  pi=207'b100001101010111110101101111110000001000100000000011100111011001100011000101111010111110111110011010000110000010110100010001001001001011110001101010011110111000101111010010111111101010000110111100100100011010;
#1 $display("%b", po);
# 1  pi=207'b011110110010000100100001110110010100000010111011101001100110100011010010010110101110000010100110110011010000111100101010100100110111000010111011010111001110000000000111110001111100111100100000011010010111110;
#1 $display("%b", po);
# 1  pi=207'b101001100011110100111011110101000101011100100011001111100000100100000011100100100100111101010111100111101011011010101000011000001100100101000000110101011001100110100010110100111100100101010111010000000101111;
#1 $display("%b", po);
# 1  pi=207'b100011101000001001101011011001110101101101111101001111100110011101001111011111001111101000000011000011010001100010010101110001000110110111111010111001010000100101000011110011010000010100011111000000011100100;
#1 $display("%b", po);
# 1  pi=207'b000001100101010010100001100011110011110101110011100010011010111000100100010001101111110100111001011010000010111000100110111100100110010000110001001100110000101000001100000000000110110010011010011110100011111;
#1 $display("%b", po);
# 1  pi=207'b000111101001000101011000000010110011000111001001110010001001000010100011101101010010100000001111000110001000011110111110111101001001010010111100111100010010000011011111010010000010010111100011000100001010111;
#1 $display("%b", po);
# 1  pi=207'b010100101001000110101111000010110010101110111111010100101101100101000011011000111101110011011010111010000101010011000011111100110011010101010110100000111101010101011110010110010111101100111101100011100101111;
#1 $display("%b", po);
# 1  pi=207'b100110011100011000011011110110110010100110101111111000010000000100100101011001001011111001001010101110010111111110001011001110100000101000001101101110110110101001101111011010010110001000111001110010011101100;
#1 $display("%b", po);
# 1  pi=207'b111000011110011011111001110000110001100010111111011010101110011110010110101100100100100111000001100000100100010011000010001010011011111111010011000010010000000100110001110111110101000010001101001011111111001;
#1 $display("%b", po);
# 1  pi=207'b000010110100011111111010100100001111001010001011100010000010001111101101011010011100110011111001110011110000001111111101101101101001111011101101011101010001110111001111111000010010100000111000011010001011101;
#1 $display("%b", po);
# 1  pi=207'b001000101111001000110001110101011101101011000101000101101101011001100011010000111110001010101010001110100101100100110000000010111100001011101000111101010011001011111001001100100100000110010010100101100010101;
#1 $display("%b", po);
# 1  pi=207'b000111011101000100000011101101110110001010010111110010101001001110101100101110000001010011001011001000101001000101101111100111001010011100101011000011101010111110101000100000011111101010000111000110001010011;
#1 $display("%b", po);
# 1  pi=207'b110011000000000001111100110000010110001110011011100110111100001011101010110100110100011111101101000111001011000000110011111000100111010010101010101011011110010111100110100010000101110101111011001100000001100;
#1 $display("%b", po);
# 1  pi=207'b110001110111001000101100010011110110010000101000110101101110010000001000001101100100000011011110010110110011000011010101010001100011110100100010000100011101011111011010100011010001101111010000001110011100110;
#1 $display("%b", po);
# 1  pi=207'b111010010100000011000100101001101001101111100111001001100000001010000000100101101101111000000100101000001011010110100110101001010000001001110011001100000100000100110000001011010100111011001001101111001100111;
#1 $display("%b", po);
# 1  pi=207'b001000011111100001010110111001110100010110001010000010110000100110001101110000100000000111000011011001100010011110001011110110101110001100111111010000110010000111000101100100110110100001001011011011110000110;
#1 $display("%b", po);
# 1  pi=207'b000010100110011011111100001010111011010100010100110100011110111010011010110001000011101111110111010010010000101110000001000110010001100000010001011101110010001011010010101110111010100100010100010111001100000;
#1 $display("%b", po);
# 1  pi=207'b110101110111110110001111100111111011000100100101010101011100010010101000101001000101011101100010101000110100011101011010101100110011101100011110110110010111010010000000010100010111010100110101100010110111101;
#1 $display("%b", po);
# 1  pi=207'b010100110111110001111010001010000101110111001001101001101111010001110111011101001000101000010000010001100111100100001010101110010111010100001001011111000111001100011011010110001000010101011001111101101100111;
#1 $display("%b", po);
# 1  pi=207'b101001011100010101000011101011000100011001110101010010111100010011001010010000011011011011101110111101000100001101111010011011001010010110001000001010110011000010011001010101100010011010110101010010011011011;
#1 $display("%b", po);
# 1  pi=207'b100100001101000011010101111011111101101111011001001011010000000111010110011000010000011001010100100001101110100100011000001110101111101111101101110101000000100000111000101000101101001000110001011100101100000;
#1 $display("%b", po);
# 1  pi=207'b110111000011110010010100000011101110100000111011111111000011110101010011100110100110110111010010110111110101100101000111011000011001111010001110010000110110101101001001011101111100111110111010010010110000101;
#1 $display("%b", po);
# 1  pi=207'b110000001000010101111011001011001110011011000010010011000010111000111111011100110110010001010100010101110101001111010110011001100001000011110001101111011011110101110001011110011000110101011100000001110111110;
#1 $display("%b", po);
# 1  pi=207'b010010001110000101010011110111110001111010101001001011110001100100110011111001101111110001101110001101101010010101100001111000100100010011011110011010011111100101001001011000100111010000000110000101101100001;
#1 $display("%b", po);
# 1  pi=207'b100101111101001011000011000110101110011001101000011110101001011000001111011011111101010100001100111001011000110111011110101111101100001110101101011011110100011111110001011000100000100011001001110111011000000;
#1 $display("%b", po);
# 1  pi=207'b001001100101001000100100001010100010101101101101001011100001000110001001001011100100110001001111101011111010100101100011101100000110010010000111010100101011111111100100000000100110011000101011010000100110010;
#1 $display("%b", po);
# 1  pi=207'b101001010010001101101101010101000011101101011110011000010010000101111001010110100010001100101011001100000110011111010101011000010010111000100000001010010011001001001010011010001111011010010100111111000110100;
#1 $display("%b", po);
# 1  pi=207'b010000000111001001000100100000110011111010110001000011100100100010111000001000101111010111110110000110100101101100010010000100011111001110100001011110100011010011001101010100000100000000110011111101110100110;
#1 $display("%b", po);
# 1  pi=207'b010110110010100111011110001111010101001101111000110001100010001101001001001100100110011100101010001100001111010011010000001011100100011101000000000100001010100011100100011111001111100011110000100111011111001;
#1 $display("%b", po);
# 1  pi=207'b111010101111100100010010001010110111110000010000111011110101111111101101010101000111010100111101001011001011100011110100011011110101010000111010001001100101010100100001110000101111101111111011001100101000100;
#1 $display("%b", po);
# 1  pi=207'b100110010000010000010101111100010111010001011001111001111100000011101110110101101110001000111001110111010100101110010001101000101010010001111000011100000100110110001000111010100110110000111100001111010000001;
#1 $display("%b", po);
# 1  pi=207'b100000110111000001110011101001101010111110111011001111010110100010111111111001111101100101110101111010100010011100011110100000000111001100000111001111011100010110000001001011100001011001001111101010100011000;
#1 $display("%b", po);
# 1  pi=207'b110000000011000110110000111101110101000110000001101100001101110010000101000011101100000010000100111111000000010111000101010010101010111001100011101011111101100001001111010010101100110110111000000100110111101;
#1 $display("%b", po);
# 1  pi=207'b100111111011001011000101001010101000100011011001001001010100111111011000000010010001001101001010000101001000000100110101100001011110000001100111101011111111111000110001000111001101000111001011111011110101010;
#1 $display("%b", po);
# 1  pi=207'b110001111000111001101110101111011101000000110010100110000000011000101010100111010100100011100010101000101111011111010010101110000000100010001100010101001100110111000011110000111100100000111000100011101100101;
#1 $display("%b", po);
# 1  pi=207'b111001111000101101000101001001101001111011000101000101100001000101110000001000001110101101100000000000011010111001110010101110011111010110111011011000001010101100011001100010001000000010011000111101000010111;
#1 $display("%b", po);
# 1  pi=207'b111100111110101111100110000010011001000100001101101101000010101101100101001010111001001010100101111010001111110010110101101100000000101111101101000001000110111011101001010111111100010010110110110000101000111;
#1 $display("%b", po);
# 1  pi=207'b000001111100101000100010110110001101011011100000011101100001101101010010010110101100101100011011011110101110011111110111000010101111101010100000111000100001110000010011000001110001101011101011000000111101000;
#1 $display("%b", po);
# 1  pi=207'b011001011100111110011111000101111111110100000110011010011100000011000010111111100100000001010000001111110011100011010101000100001100011001110110110111001110101011100000111001001001010001010000111010010101111;
#1 $display("%b", po);
# 1  pi=207'b001111111011110001100011100101111110000101111000110110101101011010011010101000110100111101010010010101111110100010100111010011001001010001100101011011110111000100110000110101011001101011101100001011011010111;
#1 $display("%b", po);
# 1  pi=207'b001011110101101110101001111000000101110100011111001100000001000110100010011010111101011111000100101000101001110011010010111000111001011011101010110111110111101000111101010110001010000001010010011001011100110;
#1 $display("%b", po);
# 1  pi=207'b010110100010100111111101100010111110000011110010010010000000111001101011011110111011000110110101011100110110000110000000111011110011000111110111000101110100011000111001011111110010101000001000000001110010000;
#1 $display("%b", po);
# 1  pi=207'b010110010101101000011101100011011000111001111101101010001111111000010110111000000101110101111111010000000101101111101000110000011000011111011100111001101000101010000100100111001001000111111001011111110111011;
#1 $display("%b", po);
# 1  pi=207'b100101011011110001110001110000011001001001001011101010010111100011010110110011001100000111101110011010110011100111110110101101001100110000110101000100111111111101000100000110101100100110011000110111000010100;
#1 $display("%b", po);
# 1  pi=207'b011100111010110110001111110110000001000101101001010011001110010000101111101000011101101011100001010110011011000010011111010000001010011111100100111110101001101001100100001001101011111000100100101100101001011;
#1 $display("%b", po);
# 1  pi=207'b001101010111101011000100100010101111111111111100010101000011000110101000000000111001110000111000010100101110111100110001010101101111000100010011111011011000010101111011010001100011001011100111101111100000011;
#1 $display("%b", po);
# 1  pi=207'b011000111000001011100111000011011001111101100001101100010101110111001010100011001111101010101101011101011000111100111010100001100001010011101001000110011011100010010100011010010110011011001100100101111000011;
#1 $display("%b", po);
# 1  pi=207'b011001101010100111110110000100010001100001111101000001011010110010110101101101101011110011011100111111101000010011011000110010100110010000111001110101101010100010110110001101100010001011111101001100011000100;
#1 $display("%b", po);
# 1  pi=207'b110011010001111110101000111000101101010001010111110111011000110101010001111011100001001100100100101001000110100111101010110111110010001101111011010111111010111011000100101111100110000001100110001100101011101;
#1 $display("%b", po);
# 1  pi=207'b110010011001001010110000010001111011010001000111101011111101100101010000011011011110001001000111110011011001110001111111110001100011011001011001110010110000011111110111001000011110101001001100111100010111000;
#1 $display("%b", po);
# 1  pi=207'b000110110000011111000110100111000100010110101001101100011011000010100110100010001111011011001001111100101000011000100011101001101011011010001111010101101011110001111110011110011110101110010100100100010101011;
#1 $display("%b", po);
# 1  pi=207'b111000000010000111000100011100101001101000000001011000001001101001000011110100010111110011000001010100010000101110100010011100111111110111001011100000001110001110110001010101011011001001110000110110111111101;
#1 $display("%b", po);
# 1  pi=207'b100000010101111000000111011111111010101111101101101000110101110000110000010011010101000110011101100101010100000010101111001011101110110011001101001000100001110001011101110101010111111010101101011110000010011;
#1 $display("%b", po);
# 1  pi=207'b000000110011010110100000010000000000101000101000000111101110101000010011110010001010010100001101110010100111010100100101100100010001001010001011010100010000011111101000010010010101110110011110001000100000111;
#1 $display("%b", po);
# 1  pi=207'b111010100101100100100111100100001001010110000110000001111100101011111100100100110000111001011110100111111001011011110000100111110110110110001101101100100101111011010011100111001101000100101110001100100011110;
#1 $display("%b", po);
# 1  pi=207'b001110010010111101000000101110111001100001000010010011100001100011100111111110011000110000010111011110011110000000001110111001110001110111100011101100001111011010001100001100000101110001011100110011011011111;
#1 $display("%b", po);
# 1  pi=207'b110011111100101011110011111100101010011010110101001100101001101100110000101010011001111101111101011010101000001001011001011101010100011001001111110111010010001001001001101111101111111100001001101010101100111;
#1 $display("%b", po);
# 1  pi=207'b110000111111101000110011000001100110011110011011110101001010001100010100000000110110001000101001000000011100100101010011001101100110010000000100101001010011010110011010011100100111101101011000010001001100001;
#1 $display("%b", po);
# 1  pi=207'b100110011110000010111110110101101110110011011110011110010100010111100100111011100010010010110011010010101010101000001111001101111001111110001011101100101100000001110101111011101111000110101110100111010100111;
#1 $display("%b", po);
# 1  pi=207'b101010100011001110011101000111100111001000110011010101001110011101101110001000110011100110001000111010000011110010101000111001100110000101100100110001011110011110110101110111110000010011101110101011100011110;
#1 $display("%b", po);
# 1  pi=207'b010011000001111100111001001110001010111000101101010011100101001000001101011110010110100101000110111100100111111001001110110111001010011010110001000011110110111000011100011100101000010001100101111101011010010;
#1 $display("%b", po);
# 1  pi=207'b011000000110011010110110000111010010101100000001000001010011000001011110011001011000000000011100100101110001101110101100000000001001101111001001111111010010100111011011100100011010010100101110100100111100010;
#1 $display("%b", po);
# 1  pi=207'b101011001111111110001100110011101100101101110011100101010000111011100011010010000000101101011101000000110001101100001000011001000110010010011000000111100101110001111001010110110101110011010111011100100111000;
#1 $display("%b", po);
# 1  pi=207'b110110110100101000010001101010001010110101000110011100111110010010000110001010100110010111100110001100101111111110011000001101001010111010111001100111010010001011011011101110011010001001000001100001011111001;
#1 $display("%b", po);
# 1  pi=207'b100111110100101110110000110100000111100010110000000011100100101000100000010001001110010011011100110110010010010111111010001100101101101101010100100100000000100010101011001100011011111111000110011011001000010;
#1 $display("%b", po);
# 1  pi=207'b010100111100000010000101000000011011010011100000010100001111011011111010011110011100000110101001100000100011101111011101001110010001000111111000111111111000000011100111100100000000100111010100111010000110001;
#1 $display("%b", po);
# 1  pi=207'b000001010011010000000110110111011010010010100101110001111000101100000111010011010101000011011100011011011011101011000110101111010100100010111111000001000011100011010110111001100001011101110110101111011100010;
#1 $display("%b", po);
# 1  pi=207'b001001101010100000001101000001111101111100110111010000111111001100001010001110101111000010010111011011001010001010011110101110100101110110110010010000000111010000001111110010011001101001010100011101101100001;
#1 $display("%b", po);
# 1  pi=207'b101010000001001101101110100111011010111011000000110010011001100000001010000101110000001010111101011010101111011011111100101110110000101111001110100101001010011010001010000100001010110111001110111111111100001;
#1 $display("%b", po);
# 1  pi=207'b010011101110000000001011101010011101011101111001001111100101111010111110101001000011001100100111101000100100100000111000111111101111001110000110110000011000011101111101001110111111100000011110001010011101110;
#1 $display("%b", po);
# 1  pi=207'b011111101010101110001111101111110101010100011110010011111110100110110000010000101010110001110011011010101100010100000110010000111011100001000111000101100101000000010110101110100111011110010111000101001111111;
#1 $display("%b", po);
# 1  pi=207'b001000001100111110000101000110111110100010000000010010001101110011001000100011100011100101001001101001010010100110010110111001011111001010010010101100010101110011111100001101100101101100000010100000000110111;
#1 $display("%b", po);
# 1  pi=207'b001110111001000111010001000100111101000101111100111011000000100011001101110101101000010011100001001011110110101111101011011100001100010111110001100100111001100001111010010011010100011010000001110000110101000;
#1 $display("%b", po);
# 1  pi=207'b010100110001110100010000100101111000001000100000100110101010010000111000111001101001101111001101111010010100111110011101000011100001000110110111111001000100101101010011001111110011011100101000101011100100010;
#1 $display("%b", po);
# 1  pi=207'b010000011111010001111100010110011110101000100000011110001000011011001100000011010001000001110101000010000000010011000101010110000111010001011101100001110010111100101100110110101011100111001110111100001101110;
#1 $display("%b", po);
# 1  pi=207'b100011101010100101010101111110100111000111000110100010001101100001010111010101100101100001110100101010010010111010000000111111011101101011110000000011111000110011011111111001010111110100000011010011011010011;
#1 $display("%b", po);
# 1  pi=207'b101011000110001001011110101110101111010011101111111101011111110011000000001010000001100001110110010010100001000100001011011101111011001100000101101000110001111000000100000101011010001011010011100101011001101;
#1 $display("%b", po);
# 1  pi=207'b001001001001111111000011000010000100011110100101100001110101100010001111101111111000001110100010111101000100100000110101010100001110101111010110011000001010101110001000100011110101011011001100100100000011111;
#1 $display("%b", po);
# 1  pi=207'b110011010010001001101101001011000001110001100101010100111001100011010100110101010010010001000111111101011111011101101101100110001001011010001111011011111011000001001000010010101011011101110101001100110011100;
#1 $display("%b", po);
# 1  pi=207'b110000000100000011001001010110011111111100100011111000000100101011110100011010011101001001010010010100000001111111000010100110011011011010110111000000100001110000101001010110001111000100110001001000010000101;
#1 $display("%b", po);
# 1  pi=207'b010001000110110000000011100100001100011111110000000110010100111000011101000001011000100001111001011000101100111101100011010100000010001111011001111011000010010010000000001011010010011001001100101011000101001;
#1 $display("%b", po);
# 1  pi=207'b001000000011110111111110110100001110010010001010001110101010001010110011101000010100001100100111110000101110110010111110111011010111000101100110000111111001111001110111000000111000011111001010101010010000000;
#1 $display("%b", po);
# 1  pi=207'b010101011010011100011011001110000010001111110010100110110110100101110001010011111011000010110000010000111111101000111110001000110011101100000101110011010110010100010010110011000001111111010100101011011001010;
#1 $display("%b", po);
# 1  pi=207'b011101010111010110010101101011000111010110001100000000010011000111111010011001110100010111001101010111011010010011100110110001110011101100111010101110100011111000001010101110010011001001111110001100110111001;
#1 $display("%b", po);
# 1  pi=207'b110100010001000110111110100011010000001111001010010110110010001100010100000111111000011110010101010110000000101000011101000010000000100001010111000110000000101000001001100100011110111011001000010110100001110;
#1 $display("%b", po);
# 1  pi=207'b011101010000100001011110001010011100110000011100110111111001000001010000101100010100010000110101110100001100000111000011100000100010011011011100011100001110100100111100110101010110010110101010101100011110111;
#1 $display("%b", po);
# 1  pi=207'b111001010011001000100101100000111011010111111010101001010011101110011001011100010101111100111111100000010110111010101111111000000010011110000010101101110111101111111110110111101101011111101010110100011001110;
#1 $display("%b", po);
# 1  pi=207'b111110000011100101001100001001111010011010000000100011001111000111011011010001001000111001110010010000000011010001101010100111001001110011110100100101110010001011011111100100101111011110100110101101010111111;
#1 $display("%b", po);
# 1  pi=207'b001010010011010110100001001101010100100111011111111000001101100100111011111000111001101110111100001111001100111110101100001010010110101101011011100100110000000101011010001101001011110100010010001101000100011;
#1 $display("%b", po);
# 1  pi=207'b000111010000100010110100010100000001011110111110000011111110001100101100100111010001001111000011110011000010010011111011100001011110010100001100110111110000000010110000001111110110101000000101111100000111001;
#1 $display("%b", po);
# 1  pi=207'b011111111010100011101101100000001101000111101011001111000110101000100111011101100101000110100000001111000011111110001110001011111011011001000110100000110010000110111110010110100000101010111100000010011011010;
#1 $display("%b", po);
# 1  pi=207'b001101100001101001101111000110100001100111011011110000100001100111101110110100000110100110001000100010010000011011001011000001100010001011100111000111100011011100100011101010110001111111101101111111100100001;
#1 $display("%b", po);
# 1  pi=207'b100101101100110110111000101000001000000000111100111111010011010001010011011101111111111011110010111011101010001101001011100011011010011111110011100100101000110010000001111011110001101110010000010100100011001;
#1 $display("%b", po);
# 1  pi=207'b011100111100111111000011010000001100011011011110001001010111101110000101110101101111110011100000000010000111100110110110001111000010011000001110110010000000101111101011000001011111000101000010000101000110000;
#1 $display("%b", po);
# 1  pi=207'b110000101011000001101111111110011001000110001110011100010001100011000000011100101100010110100010011000100110000110000010001100100110010111010010011101101011000111001010100110001000111001001101010110010111010;
#1 $display("%b", po);
# 1  pi=207'b111101010011011100110100011111010101000001111110101011111100010111111011001001101110001010011111100101000000111101100011111110111100011101000101000001110000111100011100101010110000001001011011101000101010000;
#1 $display("%b", po);
# 1  pi=207'b101010000010110011000000001010101000010010100101011111110100100100001110000000000110111010101111110101110011001010011101111010011010011000001001111010101100010011011110000011010100000011011000111111011110011;
#1 $display("%b", po);
# 1  pi=207'b111000100111010100010100110001100111000111110000000001011011101110010101010111101010011101011000100000000101000011110001100001001111101101000000111010110000011101110110111101001010000101010011010001100110000;
#1 $display("%b", po);
# 1  pi=207'b011100010010101111100001110000010101001101010110010101001011010110010000101001001000000100100110111001110100001110101000101101011010110111001100100100011101100110010111000011101011011111000010101000110000100;
#1 $display("%b", po);
# 1  pi=207'b010110110111100011111110110010000010111111000100010011010100010010101010001000101010111111000011100010100101000010111011010100011001010101111101011011000011000001101110111001110110100001001110001011001101010;
#1 $display("%b", po);
# 1  pi=207'b111011001111001011110100011011110000100101100010000001101010100000011011111100001001101101110111011010000010000010001000011110111010101111111111111011111111011100101110101000110100101000010100100110000011100;
#1 $display("%b", po);
# 1  pi=207'b111101111111001000011011010101101010001101100011010001100100101011001100101111001000001000100100001100111001100001100110001010000111111000111101100101010100111000011011100010011010000100101011010100000001110;
#1 $display("%b", po);
# 1  pi=207'b100011111110011100011100010000011111001010011100100101101100101001100110000101100000101010011011110110011001011011011111110110110011111110110001011010001101010001100110100110110100011000101000011101010000011;
#1 $display("%b", po);
# 1  pi=207'b101110111101100101101000000111001110010011000111000111101001110111000000011100110100011101001101000000100101110001111010101001011101010011111011100010111001001100011110100001011111111001110010100101011110001;
#1 $display("%b", po);
# 1  pi=207'b111110100101101100000000010011100100101011110001001010001011101010001111000001101011111001111010001100001101011000010100011001000001011000110011000001010010001011100110101110001101111001001110101101111010100;
#1 $display("%b", po);
# 1  pi=207'b001001010110011010010010001100010100101111100110010011110111100111101000011101110111101110110010110100100001000101101100001101001000000001101010100101011010001000111101111101000101101101010100111001110110110;
#1 $display("%b", po);
# 1  pi=207'b001101000010111110000100010001010100110111100010011001110011101001110001100111000001000011001110101010011010111101101000010000011011010001101011100101110101101111001110010101110010100011100011101010111110101;
#1 $display("%b", po);
# 1  pi=207'b100000110010001000010101010100100010110011111100111010101010100000011011001101100010111110000011100111111110000101001010101010110111010011001011110110000001010000011111001111000001111011100110100010111100101;
#1 $display("%b", po);
# 1  pi=207'b001101101110011111000101001001000001010111110110001100110100100101011011111011101101001011110110001111100110101110101100110011010111110111000100011000010011111110101101100111010011000010110101101100011111101;
#1 $display("%b", po);
# 1  pi=207'b101011110110010011101000001110010111011001001100001000001111001100100101110110010111110101011110100000011111010011101110000101100000100111100101001000110010101111010000111010101000111100010010011101110010010;
#1 $display("%b", po);
# 1  pi=207'b001111010111111001100000100000001110011010000110100001100111000000100101001000111110001010001100001000011001111100010001100111001010010111110101010100111110000111110101001111011100000110111100000110111010101;
#1 $display("%b", po);
# 1  pi=207'b111110110110011010110100100111000101110011000111101011110111011010000110010001100010101110101111101010111011101010001000111111100111001110101100111110101110001011000110101000000101010010100111101001001100111;
#1 $display("%b", po);
# 1  pi=207'b101100100110001000100001011110001111100101000000110110110010000000010110011001111111111001000101101100100011101101010000011101000000101011101000000011001100001100111100101000111010101001010000011001001010010;
#1 $display("%b", po);
# 1  pi=207'b110010010000111000001110000000101011100001111110010011000110001101011000100000010101110110100001110100001101000110101101110111000111110010001000000111011110001111011101011001110101100100111111000110111011001;
#1 $display("%b", po);
# 1  pi=207'b110110110010011000001110101111101110111100000111110111010011001110000111110011111011000010011111001001100000101110000110100110010110010101111000111111100110111111011010111000010100100100111100110111111001111;
#1 $display("%b", po);
# 1  pi=207'b001101011000000011111101001110000011010001110001111001100100011111011010011000001001001111100110011000010011100010110110100001100011111001100110011111010001010001111111010110100110101101101111111111011000001;
#1 $display("%b", po);
# 1  pi=207'b000110100001101101010011000101011111001010011010001110101100100001000010001110111110000101010010011110110010011100011111100110101011011001011010110100000011101101000110000011000111110111100011010011011011010;
#1 $display("%b", po);
# 1  pi=207'b000001001110110100000100111011111101011100011110011010111010000000011100000100001111011010110111101000101101101110011011000111100110001010011000001111001101010100111101100111000100010111010101001011011011010;
#1 $display("%b", po);
# 1  pi=207'b100101000100100000111000100010010100010100110101000010001100110001001100011101010010110110110011010110010010001110110110000001101010011110001011101011101010101111111101010101001111000000110011110010111010001;
#1 $display("%b", po);
# 1  pi=207'b001010100011011111111101011111110010101011010000011111010100011111110010010001010011000001110100100101000110101010011100010111110001010001111101011100001000100001010100011011001100011001111101000110111111000;
#1 $display("%b", po);
# 1  pi=207'b101100101110000101111110010110110110111100101011100001001110101100001101101010001100010010001000110111101101001110100111101101011110011000111011101110110011011011000111110011000101111111000010110111011010100;
#1 $display("%b", po);
# 1  pi=207'b000001011101001101111010011011111011101110000000000101001110001101111111110110011101101000110000110010010101001011001001111000100111001111110100101101111111001010011111101100011101110110101010110100011110010;
#1 $display("%b", po);
# 1  pi=207'b010011100111010001001110110101000010111111110110010101111111001110110000100101000110110100100011111111010110011010000001010110000001000001101110010101111100000011100101010101110110110010100011011011010001000;
#1 $display("%b", po);
# 1  pi=207'b011111101101111011110010001110100000110000110111100110000001001100100111100010000111110111010110001010011110010011000000101111010110111011110110101000100101001000111010011100111011111011000011101110000011111;
#1 $display("%b", po);
# 1  pi=207'b000011101010011011001000000011011000110101100010011110010110010101001100111100011100100011100011000011111100110011100001011101111001011111101011000110010000001010101011010011101000101101000110100100010000011;
#1 $display("%b", po);
# 1  pi=207'b000111001001110110010110011010001011110100101110110110110001001110110000111000011101000000101111110101001101010011100111010100010101110011101110110010010011100101110111011010001101011110011101101110010111000;
#1 $display("%b", po);
# 1  pi=207'b001101001011011101010001011001001111110010010100110111001110100000111100001001111001101101101001100101011101000011001100110010001100101100111011011011000101101000100100101000010111000111101100110000111010011;
#1 $display("%b", po);
# 1  pi=207'b011100111011000011101110000001100111101101000001110010011011110101001001011001101000100010110010001111100100001110110011010110001110001000010001100100000010010110010000001101101001111100111001010110001001111;
#1 $display("%b", po);
# 1  pi=207'b010101000010110100101000000000100110011011111011110011011100000011010000101111111100101010000110001000000110100000101101110101011101111111011010001111011110100110100001000001111111110011111010101111111011100;
#1 $display("%b", po);
# 1  pi=207'b010101001111000011011000010101101110010101101001001101110110011101000110011100010010111110000110011111010011111000101100111110110111000011100001100110001110111101111111101010101100000100101110110110011001001;
#1 $display("%b", po);
# 1  pi=207'b110111000110001100010110010110100111001111010101000110101000100111011000101001111011110011001100000101000001110100010110001111110100100010010111010100000001110000111100101110101001111011100101011111111110110;
#1 $display("%b", po);
# 1  pi=207'b011010011010101100111100101001010110100011011101110101101101100111101001100001010101101101000010001101101011000111111101100011000001101010011110001011111001001010101100100000111000101111100101010000101000100;
#1 $display("%b", po);
# 1  pi=207'b110011111011000100010101010001110110110100100101100010111100011010100011001101101101100111000101001010101111100010101011001011111010110110011010010000000110100101110010000100010001101111010001101100101110101;
#1 $display("%b", po);
# 1  pi=207'b011010011100111111101001010101011001101111000011000011010000011100011001100010001111110010101110011100000011001010110000110101101010100010011100000100011011011110100000011111011000010100001011001000110101100;
#1 $display("%b", po);
# 1  pi=207'b101001100111001000101010110010010010000010100111011000000110000011000011010000110000100001111111110110111000111000100101100110011101001010100110101010011110111100001000110101011100011010101111111010001011001;
#1 $display("%b", po);
# 1  pi=207'b001101000010011011111010000011011010101111010011110100010000101110011111111011011100001110111010101001010101011001000001111000100110101110110101100111100101100101001000110101101010000011010010111110011100011;
#1 $display("%b", po);
# 1  pi=207'b010011010000100010001010100111111010010010011110111111110000010110000001101011101011110000011101100110000101001010000000000101011010101011010100001011001010100010001100010111010101110110011100110011011110011;
#1 $display("%b", po);
# 1  pi=207'b000001001100011010111010011110100010101010110010100101010000111110010001100111101100011101001010000100111100001001000000000011100111110101011010100101101010001100000100110101001110001101110010001111011010110;
#1 $display("%b", po);
# 1  pi=207'b010110110111110000000001110101111100001000110110011110010011101111100001001110011101011100110100101001101101101110010101111001010110011101000101111011110000101000101011000011011001111110111001111110010010010;
#1 $display("%b", po);
# 1  pi=207'b001100011000011010000001101010010110000011101011100011110000000101010101011001100111010101100010011010010010100001011111011110111001011000100110011100101111000111001111000010100111101101010110000101110100111;
#1 $display("%b", po);
# 1  pi=207'b000111101010011111011010100111001110001010001000101101111000011100001110010111000111001110111101010111001100011111100100111110011001001101110110010000000010100101110001101011101000011100010001101011000010110;
#1 $display("%b", po);
# 1  pi=207'b010101011010110111101011111110011001101111000110001011001101111011111001110110111111001101010111011111101111111101110001101011101000100110100101001110000101011100010100010101101101010101111110110011110001110;
#1 $display("%b", po);
# 1  pi=207'b100101001001000011110011111010101110101001110110011000011000010110010110111011100111110000010101011001110101010101010110101100111011111010011011101011101111110101010111010110101010100011110100001001101101011;
#1 $display("%b", po);
# 1  pi=207'b110111111100111000010000010100101010001111111111000100000111111101110000011011110100111010100111001001011100111011000101110000001000110110000100101100111001110110011100011001000010001001001001110001001000101;
#1 $display("%b", po);
# 1  pi=207'b000011111010100111110010101111011011001001000001100111111001110100010000100010101011001001001011100101001110000111010111110111110101101110110011010110100111101001110101110111011111100111100101010011011001011;
#1 $display("%b", po);
# 1  pi=207'b100000000001011100011011111110001001100101101011010010011110100000101100100011101010111011011100101111110011111011001100110001010101100011110000101111100011000111101110000100100011011000110100010100110101100;
#1 $display("%b", po);
# 1  pi=207'b110010000001001100010001001001110010000010111010111000000110010011100000000011010010001101011010010010010000001110011011111011111110110011011010101110100011001101100100111011001010110001110101000010111101100;
#1 $display("%b", po);
# 1  pi=207'b010101110001100111100111110111001100001000110011000001101110011101100101001001000101001100001101010110101010111110111001011001110111001111011110111000001101001011011000100111101100101001110000011001111010111;
#1 $display("%b", po);
# 1  pi=207'b010101110000010010111110001000000100110000000011110101001100000111110110001001011100100001110010011011110000110111110110011101110011010011111001101001010010111100111110101110010001000010000011101010000011101;
#1 $display("%b", po);
# 1  pi=207'b100111010000011100001011110110111101110000100011000011001101111001010110011110000101011101011010110100001010011001100110000010010101000010100011101111010111001010000101001000000011001011001110101110010011111;
#1 $display("%b", po);
# 1  pi=207'b000001110110111010101000000111010111000011101001100000011000110000011000011001100100001111111000110010100011110101011010001010011011110011011111001100011001010001010011011001110001001010100101000110100101101;
#1 $display("%b", po);
# 1  pi=207'b010000001010000011110100111110110011101010110100001010011110111011001101010110011110100011001101001111111011000110111110101010011100000110100001101010110001100001000101010101111110110010110000010110000000011;
#1 $display("%b", po);
# 1  pi=207'b010110110011111001011001111011100011100100100000111100011010101111010110001011101001001010110111010111000101101110000000101110100001010000100101010111011110111000100000111101110001101011010101111010110100001;
#1 $display("%b", po);
# 1  pi=207'b111010000001110111010100111001100000110100000100111011110001010111001001110111101111011000100000111100110000100111010010011101111111010110111010000110111101101100010111001000101001110000100100011000000010110;
#1 $display("%b", po);
# 1  pi=207'b111011000110100010010100111000011110111101110110100010011110110000010010000101100110111010000100010101101000101001110001000100001100010000011111000111101101111001000010111010100000111101001101011010111001100;
#1 $display("%b", po);
# 1  pi=207'b000111111101011101111101100110011110101111111011000110101110011001110000011000000001000010110100001011101000110111000011011011101100010011100100011001100101011100101010111101100110101101001100010011100101111;
#1 $display("%b", po);
# 1  pi=207'b100111010000111010001011111101110010111001110011001011011001011110010111110011111101110101100101100110001110010000010010001111111110010100110000001100100001100110001000110100011110110100010111001111011100110;
#1 $display("%b", po);
# 1  pi=207'b011010111010011110001101001101001100111001101101110110111000111001111101011110101100011101101000100001011001010000000011011100111101100000100010101101000101111010001101010001011001111111100011000000001111010;
#1 $display("%b", po);
# 1  pi=207'b111000000001100111111000101111000101111101011011000110010010011010111001001001000101000101010010100011000100001000011000101101010001011100111100011111110101010000111001010111000110110101100010010001010011001;
#1 $display("%b", po);
# 1  pi=207'b010001110010111000010111100011100011101010000011110111101111101111001011110110111010100100001010110001011010001011110001001000110001000101101001101001110101111000010001111110110101111011011110000110101101100;
#1 $display("%b", po);
# 1  pi=207'b100000111001000011111100111001101100010001001110101001111010001111000111111110001100010111011101000111110001010111010000010010110110001001101001011101111001101101011111000010001000101111001110110011110101011;
#1 $display("%b", po);
# 1  pi=207'b110101010101110000010111101001111000110100101100011010011101110101100001100110010010111001001100011111111011111100001001001111101000001000101110011111110001000101000001100001101111000110001110101010110100011;
#1 $display("%b", po);
# 1  pi=207'b010100111100001110011000000000111011100100010011100100011100010110010010000010000010110000101001000010100111110010011011011001011100110100011010110001110000111111010101000101111001100011110000110000110101111;
#1 $display("%b", po);
# 1  pi=207'b001001100101100101100011011111000010010101111010000001101001111010011110111100111111101110110000001101000110101101011111100000110110100101100001011110000010100101101100011000011100011010110000111111110000110;
#1 $display("%b", po);
# 1  pi=207'b010011100001000101110001010101000000100011110101011101111010100010110100001101011101000000011100111111111100010011100101011001111011110111001110111111010101101100110111000011101001110011110010001001110010011;
#1 $display("%b", po);
# 1  pi=207'b111010001100001110110111111110010011011001000001101110000111011101010110010100001100101010100100000000001111100000100101110110100010000110000001111011001111111111111010001011000011101110101101110001110000101;
#1 $display("%b", po);
# 1  pi=207'b111110000101001001111000100100100100110110001010101000000100001000000001011100001111101001001011010100110010001111101101100110100110001010101011100100001100010000001010000111001011011110001011101010010010110;
#1 $display("%b", po);
# 1  pi=207'b101101010110000000000001110010101110101000001001001111111001110110110101001000100001010011110101000011000100000000100110001010110010111101100000011110101000011001010100100101001000011111000000100000010011100;
#1 $display("%b", po);
# 1  pi=207'b000111001111111100110000110101001000101110111100001110100001100100001100111000100100110101001110111001010011100111010011111001100101111101000111100011111111000100011011101001011100110100101110101011110101011;
#1 $display("%b", po);
# 1  pi=207'b111000000010101011101010101110101101011111101010100111000111010001000100010110110000110100011111111111100001101110101000011001000001101000001101111110111000001110111001000000111000101111011011101000000000100;
#1 $display("%b", po);
# 1  pi=207'b100101000000101000101010010101010101110001101010000011110111100010010101000110100011101111000010010000111100111000010111011110100100110000101101111011010110110111100010111000010010110110101111111001011101000;
#1 $display("%b", po);
# 1  pi=207'b100011000110000100101001111010101101100100001011101111111010011100100101101001101100111011100000101001101001010000110110111010011011110000110110011000001010111000111010011111100011111010110101110011001011010;
#1 $display("%b", po);
# 1  pi=207'b011110000011010011101011010101011010010100010110111010110011100110110001100111111011001001111101001001001101000111000110000000100110100010011101111000111000010010011110011101011011011100001101001000110001001;
#1 $display("%b", po);
# 1  pi=207'b101011111010111011110100100100111000010111001101000010011011110110100010111110001001001101010000000111010001101100111010011000001100010000011010111100010101011000001100111011011111000101010100010011111010010;
#1 $display("%b", po);
# 1  pi=207'b111100111101001000111010111111111001011010011111110010000011101001110110111010100001110000011110011101011000001011100011000111111011000001100111011101100010011000000001111000111111111111110101011011010111000;
#1 $display("%b", po);
# 1  pi=207'b100100110100001000010100101010011010110001100111001111100010000100111001011101101100000010100111000001100010001010001010000000100101001011000110100101010101000111100001001101011110011010111001000111110010110;
#1 $display("%b", po);
# 1  pi=207'b100011100010100100111111011010010010101011101000111111001011111110011101101010110111010010011010011100001001100110101010011001100010101110011011000001011101110001100001011100001100011100011101001001101010010;
#1 $display("%b", po);
# 1  pi=207'b000000011011100001111010110010011000001000101001000010010110011100000011100001011110101011010100011010001011110110111110011111010101110100111010101000001111011100000010001101011001110101000001100010111010010;
#1 $display("%b", po);
# 1  pi=207'b010101110010110100100011001001010111001011001010010101111010110101011000110000001100011110000001110001011001011110000110111011011011001100010111111100011110111110000000110101010111000011001111010101110000010;
#1 $display("%b", po);
# 1  pi=207'b000111110101110110011001000010100001001111111000010100010011011000101001111010010001111111111111010000010110011100101101100111110110011110101000000011111110111010001110111000011000011010111110100100010111001;
#1 $display("%b", po);
# 1  pi=207'b111011000001000010100010101011100101110100100111100100011110111011000001110100011000101011110110011111000101011111010111010000100001001011101111010000010100111011001111000000111100100111011101111011000111111;
#1 $display("%b", po);
# 1  pi=207'b010011100010111101111011011100010011111100100111010100001000111000110000100000010011100011001000101000000111100100011011010100011101010001011001110110110111001001100111111000000100010010100100110011000010011;
#1 $display("%b", po);
# 1  pi=207'b111000000001100001000010010101011011110000101110000011010100010110000010000001100010001000101111110110010000000011101110100000100011101001011101001101000111011011000110011111110111000110011100011011001101000;
#1 $display("%b", po);
# 1  pi=207'b010110011000000110011110011010000001111111011010000111111100001111011100100100100101010101000001100001010111100101010000110010000001100001010101010111000100111110100111101110011101101000011011010000110000111;
#1 $display("%b", po);
# 1  pi=207'b100110001000011001111010010101000000101010010101000101011011101101110111110010110010101010010101100101001000110010101110001010100000010110101110100100010100111111100011100101010010001110010110100001001111010;
#1 $display("%b", po);
# 1  pi=207'b000001001111010110110010100111000110011010110010001000000111001011010101010011110011111011010111011110010101110000111100110111100101101111110001000010000000010100101001110111110111100110000110111100011100001;
#1 $display("%b", po);
# 1  pi=207'b101011010000001100010110100011100101100101001000110011101000011010100001011010110110100001010111010111000001110011100001011101100000011000000101100110111100001010111011010001110011100000011101001111100111111;
#1 $display("%b", po);
# 1  pi=207'b010110111001000100101111010100111111100111101000000101100101101000000010110011000101000110110000000010101010100000100100110001111010000011010011000001000000101010011100000000000001000001010011110011111001101;
#1 $display("%b", po);
# 1  pi=207'b010001110101110011101100010101010000011101110011011000000111101010100000001010110110100100000110010000000011110101001011000110011010111011101111011100010010100000111000111000100001010010000111001110001110111;
#1 $display("%b", po);
# 1  pi=207'b111111001110010101001011010110101010001111100100001001011101001110100011101101001000011101100001001001100100000110010111101001110101111010110010110000100000110110100010010010010001011110100101000101001000000;
#1 $display("%b", po);
# 1  pi=207'b000000010010110001001101000101001110011010110111001110111101100011101100100111000011110111100101001101000010000011111111000000100101000001101101011111110010101110000011101001010100001110111111110001101110000;
#1 $display("%b", po);
# 1  pi=207'b010111010100110001111010011110000010001001000110101101111010111010111101111110000100101101100010110011100111100011110100010001000000010100101010101010100011001111010011011001100011111000001110001100100000011;
#1 $display("%b", po);
# 1  pi=207'b110001011001001000110000101100100110100101101000000101011100010100011100101101111111010001111110100111000000100111111011001011100001001010101010110110111010001101111101101111000111101001111011010001000010111;
#1 $display("%b", po);
# 1  pi=207'b011010100100111111011111100011001101101011101010000000010101101001001111101001000011100110101011100110010111011100001110110101011011100111000100111011110111110110111010100000001000010101110111000000000110100;
#1 $display("%b", po);
# 1  pi=207'b000001000000101001010110010110001101110011001001000011110111110101011000011100101111111010111101111010110100011110100111111001010111001100110100011110110100111110010111000100010110101010000001000101011010100;
#1 $display("%b", po);
# 1  pi=207'b010000100011101111110110100101100111010000111011011111010001100001000011010110101010101000110010001101110010011101101100111110011010110011010100111100101100110110011111010111111111111100000100111001111110001;
#1 $display("%b", po);
# 1  pi=207'b101000000001101101110001101011111110111000011011000100111011011010001101110110101010111010011101101010000110010000001010000001110000000010011001011011101101001111011000101100100000000101101100101010101110101;
#1 $display("%b", po);
# 1  pi=207'b011101000001011000101101100100000100111001000111110010111101010100110011001101000010101001001000110101101001000110001100110000000011101010111111110100011011101110001110001110111010100100010010110110111100100;
#1 $display("%b", po);
# 1  pi=207'b010001001000010001000100011101101010001111001110011010111100101011000101010000110000000010100001011000100001111001010001111010011110011101100011011100000001000101101001100010011000000011000100100101110001011;
#1 $display("%b", po);
# 1  pi=207'b111101100111111110101110101010110000000110001100011110110000100101000001111101111010100011101100010010101110010100110111110101100101011001110010010101110000000010011000000100100101100011110000000100010100110;
#1 $display("%b", po);
# 1  pi=207'b100011110101111010100111100110110000001001111011110101100001001111101011000001000110001110100100111110111011100101101000000001101000011100111011001011110101001110111010111001110011010110001000011000100011001;
#1 $display("%b", po);
# 1  pi=207'b000000100010110101101101010011011000010110000010111010100100111101111000010010111001110110001000110001111111011111011000001001011001001010100110110111000100010011101110101011101011011001011001010001000101111;
#1 $display("%b", po);
# 1  pi=207'b011000100010000110110000101111100101000000001111100100000010101100100010100000010000000010101001000011110001101111110010001101101110011111000011000010110000001010010011000001101111111110100000100000011100010;
#1 $display("%b", po);
# 1  pi=207'b101101100101011001111100101000111001101110001011001010111110100001110000111010001110001101110010100111000001000001000100100100010100011011100010010010001001001010110000001101010001101011000010010110000000110;
#1 $display("%b", po);
# 1  pi=207'b100001111110001000101100111010010011000010100010011111101111001011000011011010000101111011010101011011110101001010101110011011000100101000110000001010100110111000110011000001001001000001100111011000010010010;
#1 $display("%b", po);
# 1  pi=207'b000111011000110110001101111000101100010000010001001010010011011111010010110010111011101100000010101001101100010000101110100011111100010000111110010100011000011011001101101000110110011001001011110101101001010;
#1 $display("%b", po);
# 1  pi=207'b001100111010100010110010101011010010000101001110100101001111010010000100011010101110111010011010011011111110100111000101010100000001100010100101000011101111001111110000010101111010111101110100011100111010101;
#1 $display("%b", po);
# 1  pi=207'b101111001010100101111000000101000011100111101011111011101011011100100111100100011101110101000100001101000110111111111000011000100011011001000111000010110000111100101100011101111000001100111001100001110000101;
#1 $display("%b", po);
# 1  pi=207'b000110011001111100011010011010000001010000110011000110000010110010111111011001110000101000111110001111111101011001111010010011111001010000010011011100000111001001110001111001111011010111000110101001101100000;
#1 $display("%b", po);
# 1  pi=207'b000001011011111000010011110111000101110001110110000001001000101000000010111000010011110001001010100110101111011110010100101101110101011101010111001111011001011110010101111001001101010110011010111111101010110;
#1 $display("%b", po);
# 1  pi=207'b010011010011011010001001000101111100000100111101111010111110000010101110110101100000011111000101110110110010100100110110010010010011011110000011111011101011110100101110111111010000000111111001101101110110001;
#1 $display("%b", po);
# 1  pi=207'b010111001010000110001100010001010111101111110100110100110111100111111011000010101001111010101011111000100010011101111000001011001110111011010111000100101010110101011111011000100101011100001101010100101111000;
#1 $display("%b", po);
# 1  pi=207'b011101101000100101000111010110011000111111110000011110101001100101111100000100111000011110000111000000100101011010001111010010000011111101101001000111010000111101000010111101011101000010010111111110010001101;
#1 $display("%b", po);
# 1  pi=207'b011101101001100100001111101101101000000110001101010010110001100010001110011011110100000000101011111010100001110110001101011001010011110101100001010001100110000110100001011101001001010101011100111011010100100;
#1 $display("%b", po);
# 1  pi=207'b110110100101110011000001000101001010111101000000111010110101110000010000001110001011111101001001100010010001011011001011011100001011101101101101110000110111000101011100011111010010110001001111111001001100001;
#1 $display("%b", po);
# 1  pi=207'b111000001101110101000101010111111111101001000000001100000111001011011100000011111001111111001111101011100110010001110111110111000111110110001001000011010011000110111101110001010110010011110100000100100010001;
#1 $display("%b", po);
# 1  pi=207'b101101100000011001010100000000001101110000010111011110001111010001000001111100000110011101111001100010001010010100100001100010001100110010101001010010110111100000101000000101100100001101111010010101110010110;
#1 $display("%b", po);
# 1  pi=207'b001110000111101001111110101011010111000110010100001011101000000100101111110010110101101011101011001100110001010101000000101000011000111100010010001101011111001110000101100101000111010010011110100011001010111;
#1 $display("%b", po);
# 1  pi=207'b110011010011100100011001100111111010011110100111100110010001110000000100000011011011100000000111000000001110000010011010001011000110110011010110111111010111000001000111000111111001010111111001100110100110000;
#1 $display("%b", po);
# 1  pi=207'b011110111101110011010110011001110010000011100010011001011110100111010001010001110110110000001100111010000010111000011010100100100010010101001111110111111010100101001111000010001011110010111101011110110111101;
#1 $display("%b", po);
# 1  pi=207'b101000101010001001100010111110101110100000011001111110110001010110101110110010001100000001101101000000000001101011110110100100011111100001001001011001111111101110000100110100100101001101000110011011001110101;
#1 $display("%b", po);
# 1  pi=207'b101101110110010001101101000101101110000100010000000101100000011101000000010001100111100110000100101101011101110101000101010011101110010010011101001110001000011011101111100100100001011010110101110110010010110;
#1 $display("%b", po);
# 1  pi=207'b001001010001001011110001100000001001011001000010011111101101011111101100011110000111101000110110110111010010001001000111101111001110010111110000110000010000001101000100011110010010011101110100100011111011000;
#1 $display("%b", po);
# 1  pi=207'b001100000110110100000011000111110101000111001100100100110001111001011011100011101011111010100111111001110001011110010100011100000000000111011000010111001100010010011000110010000010011101001011001010110001001;
#1 $display("%b", po);
# 1  pi=207'b010011100011101111101101001010111110001001000000001101001100100000000101000010001101000111000100100001111010001000111001000001001001000001010111000010010011100101000010101000001100001011111110011110111011010;
#1 $display("%b", po);
# 1  pi=207'b100000001110100100111010001011110001110000000101000001011010100011100011011110111111101100001110011100001010010101111001001111110011101100111001101010010101101000110101100100100010001111100111001111010101111;
#1 $display("%b", po);
# 1  pi=207'b000001000100000100011001011000010011101010101100011110010010010010110011011111111001101111000111110000011100010000001000110100100100111001100010010111110110110001000011011000011100110000110100011000000111100;
#1 $display("%b", po);
# 1  pi=207'b001011011010010110010111111100011000011000110111100111100101101000101111101001010101100111001010010111001111110011110101010011000111011111011011000011100111100100110101110001100101000001110010110011101100000;
#1 $display("%b", po);
# 1  pi=207'b110000000010101100011011010100100001110000000111110111001000000000011010110011001011000010001000101101010000010001100011001000000110011000110101000001011101010010110110011100011110000100101010000010111101111;
#1 $display("%b", po);
# 1  pi=207'b001111010010101100110001011010000101000011110100111011101100100010101010001001101110010110001101000110000111010110111011100011110000001101110100111000101010101100111110001001110010001110111011010001100000000;
#1 $display("%b", po);
# 1  pi=207'b001011001001011111101111100011110000001011000101000000001111101001110011000001111101000000011010111001001000100001001000010111001011111000111011001011101000010101100010010111010111011001000011000001111000110;
#1 $display("%b", po);
# 1  pi=207'b100110001111011111001010101100000110110101010111000100101000011010011010101001001001010100010011000011000011011111010101011101001001001010001000100010011111111001100111111001000110010010011011100101101100011;
#1 $display("%b", po);
# 1  pi=207'b011101101001101010100111111000101111111110110100010010011011000001100011000001110101011111111101000000100111111011110011001000110110110011001100111110011111010010101011001101001010111100000000111000111011011;
#1 $display("%b", po);
# 1  pi=207'b101010001111111101010110100010101101000101001000110111000100010011001011111000000011011000010110010000011111101010100010011101010010111111001001001001001111101100010000100100100001000010111000111001000011100;
#1 $display("%b", po);
# 1  pi=207'b111001100010110101101101101011001100010101011111101000001000011011100010101010001011010111101100000111011101010000000000100100110001011011010101110101011100100101011100001001001101101011011110111110010100100;
#1 $display("%b", po);
# 1  pi=207'b101001111110001011100100100100110101010011101101000110101100111010111001000101001010001100010101100100111101010101010011101101100100101011110011011010100111110010100111010001011000100110110011001100000110011;
#1 $display("%b", po);
# 1  pi=207'b101010111000100101111010000001011001101000111111000001110000100110000011011011100010111000000101110110000111001001110101110000100001001100011101111111110000111100111010111011000101001101111001000010110011111;
#1 $display("%b", po);
# 1  pi=207'b111011010111001010110111111110000001101000101011011001111100110000100001000110101001100111110011011010110101100001010111100100101000001011100110111000110010111111010111001011100011101100000000011000011111111;
#1 $display("%b", po);
# 1  pi=207'b010100101100010010111000000010000101001011000010001011011010111100110110000011011000110111110010000001111000111101010111010110001101000001001010101111111000010101111001011011111100011101100100110100010111011;
#1 $display("%b", po);
# 1  pi=207'b111101010110001010101011111000011101000011101100011010001001010110011010101001011101010110011101010101110011111001001010110010101110001111100100001100010110010011010001000110110001100111110010001010000110101;
#1 $display("%b", po);
# 1  pi=207'b011000111001010100000011111110100111110001010100001100101110001010000111000011110011010000001010010011000011100110100110101000101110100011111101011010000110101011011010011101011001000010011100110100101100011;
#1 $display("%b", po);
# 1  pi=207'b011101100011010100100101101100111010100000000010011110101010111001110111011111111101001101110100011000100100010101100000010000010011011000100001100100100110000001011011011101111111001100010111010010001000111;
#1 $display("%b", po);
# 1  pi=207'b011100101110000000001000110000100001101100011000001111011011001110010001100000101110001100000101001011000010000101000101101100101000111100010010001110000111010000011011000111110010010010101100001101110100001;
#1 $display("%b", po);
# 1  pi=207'b000010011101111101110101100101010101010100110001110001000011001000001111011101101010100110001111100001000101010110100110000110010110010110010010010011010111110000111001000010011001100010111101111110011000111;
#1 $display("%b", po);
# 1  pi=207'b001110000110111001000100110111111110111111001110001101110011110111100100011110010111100100111001101001111001101101000110111101110100010001111110000011110101101000100111001001110101010001010101011110001011101;
#1 $display("%b", po);
# 1  pi=207'b000101101101001101101000100100111011011111111111100100101111101100001100111001000000011000110110001001111010100011110001111011100101010011011010100110011101101111001110011110111001010001111011001011010101110;
#1 $display("%b", po);
# 1  pi=207'b001010011010100100001100100110111101111111101100101101011100110100010011000101111011111001110111100000101101101000000101010110001101001111111111110010111011011100000000011010011100011010100100010110011000001;
#1 $display("%b", po);
# 1  pi=207'b000010101000001000011101101110001101011101011111100011000101111111100010111101101101101101001100101110011110111001011110111110010010000100110001001100001101101010010100101001001111110101001111000001000101110;
#1 $display("%b", po);
# 1  pi=207'b010100110000100111100101110001111111101101001010111000100000100011101011001110100001110101111000101100010100101101011111111111000100010111000001111111010010100011100101111100011101111011001101101111100110011;
#1 $display("%b", po);
# 1  pi=207'b011000000101101100100100010011110000111010001111001100010001101010111101011101001011001101000011001100101001110100111000010100100011011111000110110100011010101001110100001110011110011111110000111001011000001;
#1 $display("%b", po);
# 1  pi=207'b111010010000001001110011011011110111110100111100011010000101001101101000011111001110111001110011111000100101101101001100111100001110001011010001111110000100000000110001011000011101111111101101010110111001000;
#1 $display("%b", po);
# 1  pi=207'b000011000001100110011010001001011110000000101001111010100111000011111111110111110100000110011111010101111011100100110111000001001000011011000011000100110010100001110111100101100011100010000011011010111100010;
#1 $display("%b", po);
# 1  pi=207'b111101101001011011101011101000010001001001001010100011001110100010100111110110000101110000101000101011001100000110110011110000011101100101101001011011011001011101010010111001100110011010100101010101000110101;
#1 $display("%b", po);
# 1  pi=207'b100000101100000101101110001101100101110000110010111010000001001001111100011100111110110110101000111101111001101001001000110111101101101110010011011110001001111001000001110010111011100101000100000011010000011;
#1 $display("%b", po);
# 1  pi=207'b100111101110110000001011110011100100101011000010101110010101101010111010111000011000100111111010100100101000111010111110111110100110100101001010111110100101100011011111111000111001001100000001111111000000100;
#1 $display("%b", po);
# 1  pi=207'b101011110011001000110001010110101001111110011001011001001001101010100101010100100110111010100101100000001100100100111001101011111011010010111101111011011011110100100000101110000010111011000110011000110110001;
#1 $display("%b", po);
# 1  pi=207'b111000000010010111000100111101001110010101001011010000010000011010111100100011101100111011111100110111001000011101110011110110101001110110111110011100001101000111101110000010111010111110101000001000100000111;
#1 $display("%b", po);
# 1  pi=207'b001010101011110000010101100101100000011101010100110100111100011001001001011000010000101110101000010000011011110100011110001000001101000001110101110001001011001100011111100000101011010110100011000011100111001;
#1 $display("%b", po);
# 1  pi=207'b100101010001100010001111001010001000110100101101111000110001100001011110110100011001110010100101000011011100001000011110011110001011100000001001100100110100001010101000100010001010101000000000011000110100001;
#1 $display("%b", po);
# 1  pi=207'b001100011110010101100011010011011101000011110011100010000001000111111010011111101010111010101101101110101100001000010001011010011110100111110101010011010101010111101011111101010000100111110011000001000011111;
#1 $display("%b", po);
# 1  pi=207'b101001100001110101010001011000101010001100101011011111011100111001000011111010100101010011000111101111110001101000000000101111001010101100110011111000111011100000000101101100001111010100011101111010010111111;
#1 $display("%b", po);
# 1  pi=207'b011001101010010100100010001111100110010010100001100010010011110100111010111011001110001000101100001101000011101010000000100000110111110111000001000011001110011010111001000100111010000101000110110100010011101;
#1 $display("%b", po);
# 1  pi=207'b010010111001011000010010101100100110011110001100100101000010111011000010110111111101100111010110100100101011010111110100011111110010000100001101100100011000010100110000000111101111011000011011010000000100000;
#1 $display("%b", po);
# 1  pi=207'b101111100001010000110101111001110110110110111000101001010010101000011000100010110000110111110101100000110010000000110101101101101111100110011111011001100010111101010100001101000010011100111001110011000100111;
#1 $display("%b", po);
# 1  pi=207'b110110110100001111100100001111001101111111100111100010010000100110110001111010011110110101110100111001100011101000011001001100111001100010010010010101111100010000111011010100011010101011111101010110110110111;
#1 $display("%b", po);
# 1  pi=207'b100101011001101001011110100101110101111101110000111010000001101010101111001001011101010001010110111110010100011011100011010110100010110001101101110100000011001001101111110011110001110011011100111010011111010;
#1 $display("%b", po);
# 1  pi=207'b000100110010000100001010010101100011100101101101110001000111111010111100000101100011111001010111010010001111001010001101111001010000110011110011110010111001100001111001000110101000110011101001111011011111101;
#1 $display("%b", po);
# 1  pi=207'b101010100000100110101101001011100001000000101101011000010111000100111100101010110011011010010000001110000011001011111111100100001011101110010101110011001000001101110000010010111100111101101100001111010000011;
#1 $display("%b", po);
# 1  pi=207'b000111100110100100111110001100111000111010010101000111011001100001111111100000010010111110001101110110010010111101100000000010001100110110111011011010111010010111010010000101100100000101100110000100010011011;
#1 $display("%b", po);
# 1  pi=207'b001110110010011000010011001001110100100000110000110001011010001010000111000000010100001101011101010001011110101010000011100001100001000100010111110011001000010011001110111110111111001110011011000000111101110;
#1 $display("%b", po);
# 1  pi=207'b011110000111101011000011100100101001101110110010110111011000101000001110001000010101010000011000010100001001001101010000001111001100011100011100101010011000000111111110110011011100111101110111100100111100011;
#1 $display("%b", po);
# 1  pi=207'b100111110100011100000100001100000011011100110101110100000001111011100101000010010101001101001001100000011101111100100111010010111100011010100011001100101111000101001101001011011011100011011010111011101100011;
#1 $display("%b", po);
# 1  pi=207'b100100000100100110110101000011001111100000001111110101111011110000010011100110100010100101011101111001010111010111011111111010010011011010010100001011110100000001110100000111111100100001111010001011010000101;
#1 $display("%b", po);
# 1  pi=207'b111111111111100101000001010010011100000111100011110100100101110111011100110011010011001010101001001001101101010000101011001011010100111011011001110111111010001011111111011111100010010110001110010101001000011;
#1 $display("%b", po);
# 1  pi=207'b011001000001011101010100001010010101101110101001011001110011010111001001100000101001111001000101010010111111101010100000011010000011111101110010110100101010001010110111010011100011101001101100111001101001111;
#1 $display("%b", po);
# 1  pi=207'b110110000000100011101011111001101111100101110011100100110011000001010011010111101000110010010010101100101010000000110000001110100010100001101011011100010100101100101111000101110001100111110010011111011111111;
#1 $display("%b", po);
# 1  pi=207'b111110100100000110101001111011100011111101011001000011110101110101100100110000010100110101000011010110101010110001001000110010111111100010001010101000110101010000111110011101001111001110111001001010110001010;
#1 $display("%b", po);
# 1  pi=207'b001111111011110001110111101101010110001110110111001010111001111000010101001111001101111011110001110101110101001110110010100010001111100110100011101101011011100010011111111011011101001000111000110111010100010;
#1 $display("%b", po);
# 1  pi=207'b001100110101100010100100011000011001110100111101000111000000000010111010010010101110111100001110110100011100011000101110011000010100100100010110010000100101111001001010101010000010001001010111000000100011010;
#1 $display("%b", po);
# 1  pi=207'b010111000011100010101001001010101000010111001000001111011101101101000001010111001110110011101001011111111111110010000111100011011111010001000011010100011000001000001101011110001101011000101100000111000011011;
#1 $display("%b", po);
# 1  pi=207'b000010010000110101001010110101100111010011110111110111001101011001001110011100001000101011011010111010100101101011111100011010000111011001011111010100100011111111011000010010111010001000011000101011100010101;
#1 $display("%b", po);
# 1  pi=207'b011101000011111010101100100110011011111101011001011111110110001000001101011100010110101100101110100000010101011001110111000010000110000011111111000000011001110000000110111000101100001000101101010011001011000;
#1 $display("%b", po);
# 1  pi=207'b111001111111000110001101110010011100001001111011100111101010111111100010000001000000011001000011101111000000010101001101101010011110100010001010111100011010010001101110000110000010101001110000111000010011011;
#1 $display("%b", po);
# 1  pi=207'b101100011010000011111111001011101010010010110101100011100100111001011110000011011101100000000111100100110101101101100100010001010110100000101101010111100100011010000100101010110000110111011101000001110110111;
#1 $display("%b", po);
# 1  pi=207'b100100001011001010100111011100010010000100000110111101010101011110011101001010110010000111111000110000111101010101001011101000010010100001110011010100101111000101011000011111011011001010111110000100101110010;
#1 $display("%b", po);
# 1  pi=207'b010000001000010001100010111100110110111010010001001001010110110000011101110110000100000101011100101111110110110111000010011000011101111100110101001101111111001110001010100010111000110111011011000000000111100;
#1 $display("%b", po);
# 1  pi=207'b011101010110000010001111111000001100100011010010111110001010010100101101101001010110000110111011001111001110010111001101111110110001011100110011001111101100001110010111100000100000101011010000100100011110000;
#1 $display("%b", po);
# 1  pi=207'b001111010011101011001101111001001011001011011110010100011100100011000011110110011101011001111010001100010000110001100011111111000011111101101001010010101110000100100111011101110111110111111011111110001101111;
#1 $display("%b", po);
# 1  pi=207'b110010010100110110101100100011110001100101101010110100110011100001011100101110000111001001001000001011111000101000010011000010101010001011000111000001110000011001000101000010101000001001110110001011100010101;
#1 $display("%b", po);
# 1  pi=207'b101000001001100110011001111101110010001111001010000110000100000001001100011101111100111111011000100010101111101100011001111111010010111101000101000100000100001100001111011001000011111000111100000011101100100;
#1 $display("%b", po);
# 1  pi=207'b101010101000011011010011000101110111001100010001001001100001101001001100010110001010100110111111101001101100100100100110101010111011100111100111000111100000100000011110000011111101011110101111100000110101100;
#1 $display("%b", po);
# 1  pi=207'b000011100100011100001101100101000111010110100001011100011011011000010100011110010110100111111000000111101111111000010001111010100110110110011100011111111011001101110111011010010110110110100010011010100110000;
#1 $display("%b", po);
# 1  pi=207'b111001000011000110000010001101110001010011111100001110110000010110010001011100011010010011110000001011110001110101101111111100111001010000010010100000010101110011000110000110110110110110000111100111111100010;
#1 $display("%b", po);
# 1  pi=207'b011010001111001101000110011101011001110110011000010101011111111000001011100010101000001010110000011111110001100001110001011011100010101101001001000011010000110110000000001111010010110100100110010111100100110;
#1 $display("%b", po);
# 1  pi=207'b011010100001001010000111100011111001000001110001010100001010110011101101001000100011001101101111011000001110001110011101110001010101001000001010011101100111101010101101011111000110010101110001010001000111101;
#1 $display("%b", po);
# 1  pi=207'b111011111110101111011011000000101010101001011001100100111111010100101100010011101001010000000010101100101101010110101111111100011110101011000111101110110011000010101000110001101001011011011011111100101110000;
#1 $display("%b", po);
# 1  pi=207'b101011010111000101011001011011100010001110100100110110111110100101110000100110110111010000100010111100010000111111100111110010010011001011100101000000001011100100111010111001101001011000110101101001100011010;
#1 $display("%b", po);
# 1  pi=207'b010000110011110000010010000010000001000111010011101000100010000010001000001100101111011010111010111100110001100101000010001100100111111001010101000000011100000011100000010110010010101110101100100000010110010;
#1 $display("%b", po);
# 1  pi=207'b000010100101011011110001000001010111001010001111100110110011010011001101001100101001011001101111100001000110100001000001100110111101100100111000101011011011101000111101101001111100011001101110111111111110111;
#1 $display("%b", po);
# 1  pi=207'b100110011110000111110110111011010101111010100000100001111101000100000001101000111000101000011001110011001101101111101110111011010101110101011011011100001001101001101000100110100011000001001010011111011010100;
#1 $display("%b", po);
# 1  pi=207'b101000010111000001011111011100101000100011101011011110100111011100000111010010011111010000011001011110101011110001111001011000001101101010100011101111110100000010111110011111100001111100001101000011010010010;
#1 $display("%b", po);
# 1  pi=207'b110101001100111100001111100001101101011000111111101011101010010011110100110111111001111001000010010010111100011111011001011100100001001100111011010111111011100111000011100101110010011010111101100010110101101;
#1 $display("%b", po);
# 1  pi=207'b110001100011000010100110101000011011101111100101001001101001100100010010100111110100000101001000100011001001111111101111001100001111000101110010101011100111001000001111010001110110000000101101011111010001011;
#1 $display("%b", po);
# 1  pi=207'b111101000010011010000111010001011110001010010000100110100100010101111001101010111110111011111000000100110011110110111000111010001111011110111001000010001010000111111010111000110010111001010001111100001001100;
#1 $display("%b", po);
# 1  pi=207'b001100011011111101011101100111101111010110100100010101000111101010000100101001010011001100011011101111101111010101001010001010010110000011101101001100111001010100111010010000111001111111010111100110010001111;
#1 $display("%b", po);
# 1  pi=207'b010100011001001111111010111000110010010001001101000001100101011001100101100101001001111000101011011100000001111010000000001100100000011001110010000001001100100101001110111100100100001000110111111111011010000;
#1 $display("%b", po);
# 1  pi=207'b110010110101100000010001011011110111110000011001111100101001011011011111111001010100011000010001010011001101010101100101011101111111111010001000101011100010010011011111110101110001011010011111010110011000010;
#1 $display("%b", po);
# 1  pi=207'b110111110101100001110001000001000101100001111010000010100110010010101011110111101110011100001011101011100101000100010111001000001010101110001001010011010001110100001110010111111100000001101011100000110111110;
#1 $display("%b", po);
# 1  pi=207'b100101000110011010110010111111011101011001000101000000010100110100110111101010001100001010010010111010010110010101011100110101011010001000010000101101000111110110001000011001011010101000110001010000111000111;
#1 $display("%b", po);
# 1  pi=207'b101000001000001100010001001100110010111100101010010111100101101000001010011011111101001010101000010101110111011000100010111010110100011100111011101001001011111110011011101011110111110001101111111101101011011;
#1 $display("%b", po);
# 1  pi=207'b011110010101100000011001111000111111000101101001110110000000001101111100100111111100100100111111110001000111110101000001100101000101110001100101101111010000001100100101110101111011000011101101011111101101000;
#1 $display("%b", po);
# 1  pi=207'b111110001111100011101100101100110100100100001111011001000100111111000001110000100011011001011010101111011100000011011010111011000100111100010001010101111111110001110011011111110011110100010101010000111110011;
#1 $display("%b", po);
# 1  pi=207'b010010111101100000101011001111110000110001110011111111101111000100010110111001100111010101001111101110111111001001101111001011111001000101111001001010100110001101000011100101011100010101010011011001101100111;
#1 $display("%b", po);
# 1  pi=207'b101110111100010011110101010110011100100001100011010101100001101001000111000010100011100000111101111100101000011000110111011000010101111011100001011010010010110001100100010101101100000000111010011100101001011;
#1 $display("%b", po);
# 1  pi=207'b000111100010111111110100011100010100110101011111010000000011101000000010110100100000111110111100010001001101111011010011110010110111100001100010010110000110010000001001110110011001111111010010001011110000011;
#1 $display("%b", po);
# 1  pi=207'b101111001100000011100110001111011110101111100001010110100000010101010101110000000001011001001011011100101111010010101100011100010111010111100001100111011110111101001001001110000100101100001111011000111101010;
#1 $display("%b", po);
# 1  pi=207'b110011000011011110000000100101110111001000001101111111001011101111100000000010110101011100101101000100010011101000001100101100010101010100010010001010110110101111010001110101111111001011001101101001000101011;
#1 $display("%b", po);
# 1  pi=207'b001111010000100011010110110001101101111100010010000110100110001011111100011110001010001000000010100101011110100111011010110010100001111010010101011110001010110001000100010001111010111000011001100100010111101;
#1 $display("%b", po);
# 1  pi=207'b111010011001011001101111100001001000011011001101000000001011000010011100011010101001010011000001111001010001111111000000011101011011110010111010110111100001110011111001001010011101111100100010001111011110111;
#1 $display("%b", po);
# 1  pi=207'b011000011011110001101110111101110011011001000101110101110011110110001100011011000000010000100000111001011001001110001100001111000010010101110110101010111100100111110011101010001101111111101110101010011101111;
#1 $display("%b", po);
# 1  pi=207'b011011101011010000101101010010010001000111110001001011001001110110111001110010111001101101011111010010001111100001001000101001111111111101111101110000001100000100110100001111010000110110111010100110011101101;
#1 $display("%b", po);
# 1  pi=207'b000100001001011001001100011100111000010100111010101110011111101101001011110100111011010111111001000000110110010011011010001100101110011111111101110100011111001100111000001101111111010100101001010100110010001;
#1 $display("%b", po);
# 1  pi=207'b100001001011011000100111010011101010111000001000000000111101110001101011101111110100101011101101010110101001010110010110011001000111011100000000011011000111110000001111111111000000001001011100110110110110011;
#1 $display("%b", po);
# 1  pi=207'b101110011000111011000101100110011011000101101101100110100101010001001000001000010100110101100100010101010111000000011101010111000011011100101101011111100001110000001001000111010101011100001011001100101111000;
#1 $display("%b", po);
# 1  pi=207'b100000000010000100101011000101100001111101000011100001010111101010110001001110110100111111000100101011110011000001001110101111110000001001110010001110100110100010001010010100110010110110100101000010101000101;
#1 $display("%b", po);
# 1  pi=207'b101100110010100100011011101101011010100011000100100110001011111011100100011101010001110001010101110100010010100000001101001000001010010011001101110100001010101101100100101100001101110111101101011111111001001;
#1 $display("%b", po);
# 1  pi=207'b001001111011011010111010011100011000001011100101101110011100011101100011100000011100101110110000011110110000101011010011010100110010101000101011110000110000000100111100101100100011001111001100000001100100000;
#1 $display("%b", po);
# 1  pi=207'b100101011111011100000001010000110100001111000100111000101110000101110101110111101010011011010011110001101111001001000111001000101101010000001101110010011101011100100011101100101000011100011111010100111010000;
#1 $display("%b", po);
# 1  pi=207'b111111110001011001111011110011011001100001000010110100000011010101011010111001110010000100101101110001100101000011111010100011111101110000000101111011000111101001011101100011110101010101101000111000011000011;
#1 $display("%b", po);
# 1  pi=207'b010000010010011101011011001000100000101000100110110001011010001001011011110100100000010001100101000111101001110111101000101011001011111110000011111000110100101111011101010101010001100111000011001101110001110;
#1 $display("%b", po);
# 1  pi=207'b100011101010100011000100111111110000100011001110111111010100011101000111011101011010000111110001100101100110111011001001000100010010001011000011111110011110011010101100101100011001111110110011110010010010100;
#1 $display("%b", po);
# 1  pi=207'b010000011110010000101100101100111100110101011001101001001110111110011100000010111100110010000111101110100011110110011001100000000000101001000101100110111010111001000101100110000110111101111011001010000000011;
#1 $display("%b", po);
# 1  pi=207'b110101000011001011111011111110100011010010001011100111010011111011001111001010100000001000101110101010000110000101000110111000010111011001001010001010110011101110000110001111011100011111110011101111110010010;
#1 $display("%b", po);
# 1  pi=207'b101111010000001101110010101101110101010010001000011110111101001111001001100101110011101010011011010110100101110010111001000010000110101000001101100001111101111101010010111000111011001111111110001111010110101;
#1 $display("%b", po);
# 1  pi=207'b111100100110011011111010101011001011100001110001100000100001000001001001110101111111010101011110111000111011000000100100111000011000111101101011010110001010101101000101001001011100000100000000010111100110000;
#1 $display("%b", po);
# 1  pi=207'b011100000001010001010010101100011111100010001101001010100100001001101011111111011100010110100001101010011100001111000111000011111101101101110101110110011010010110011000011010001001100000010101110000011100000;
#1 $display("%b", po);
# 1  pi=207'b111101001100000100000100110010110110101010010000010000001011101101111000010011011001111100101011111100001100100001111101111001011111100010111110011010111101100101100110111001011010101101101001011111001110110;
#1 $display("%b", po);
# 1  pi=207'b010101010111011101110001001001101010000111100110010000111011010100111100011110100011010100000011011010100001011100101100000110000001010010110000001010110000001010101101001111110000101001111010111111001101101;
#1 $display("%b", po);
# 1  pi=207'b001011011101100001001100101000101000101101011110110110000010101110111001011000010101100000010010100111101110110001100101000100010101010100011100010011010000001101101111010111011110001101011100011111111111001;
#1 $display("%b", po);
# 1  pi=207'b010010010000010101100011000011101011101110000001000100000111110011010010001010010110011100010001100111011101001011100011011011110110010101100111110010110001101110000100010100010110000101101100011001010001011;
#1 $display("%b", po);
# 1  pi=207'b101001000111100100011010111000100011010100001010101011000001000010011100000011111111101000001101010110100001110011111001000011001000011100110001110111101111101010110101001001101000000101100111001110110111001;
#1 $display("%b", po);
# 1  pi=207'b100011100101110011001011101001000001010000100010011001011110110001010010011110101100011111010001000001100111010111000010001001111001101100110110101101111111110011110100110111010111001011110010000110010101111;
#1 $display("%b", po);
# 1  pi=207'b110111000101111110010001000011010011010001000000001010100011011101100110001000111010010001011110100000010001000000010111001101101011111010010000000000001100101011110011001110000011011110101111001010001110101;
#1 $display("%b", po);
# 1  pi=207'b001000100101100011011110101000010001010000110001100100110111010001110011010110111010010111011000101011000100001100010011001001100011101100011011111101100100000110000000011010011010110010100101011011011011100;
#1 $display("%b", po);
# 1  pi=207'b101000010001101010010110101110101001111001001111011111010011001000111010110111101000110000110010011010010001100010100111000101000100011101100011111011100000110111000000110110100011010101111010110111100000101;
#1 $display("%b", po);
# 1  pi=207'b100010010110111011110010010010000011100101101000000100010010011101000001100000011011001110011101011000011010101000011010001001110001011101101010110011100100100011110100000010000010110000010110001010001100111;
#1 $display("%b", po);
# 1  pi=207'b000110011110110011101110001111110101001111011110001011000010101011111010111101100101110100100011110001100111010111110110100000101111010110010100001101101011111000011101000101101101110011010000100101110100101;
#1 $display("%b", po);
# 1  pi=207'b011010010111111100010000101001011000100100101110111011011100101101000011110000110100011101000010101001001110111101010110101101011100101001010101011101110110011101000010110111000100100010110010010010101000110;
#1 $display("%b", po);
# 1  pi=207'b111000010110011011000110000100100101001110100100110101000110001101101101101000101001001111000010111011100001011000000011010101101100010110100110111001111111100110001000110100011100101111110011110110111011101;
#1 $display("%b", po);
# 1  pi=207'b111100101010010001000010001000111110111100010001010010001010001100000110110101000100011111110110111111110101111010111111101001010101000101001101010001110100101111100111100110111010011110110101110100100110101;
#1 $display("%b", po);
# 1  pi=207'b111000011001000000111011000100001001010101111100011100101010110111110101110101101111000001111011111100000111110001101101101101000101011110101010101010010000110000101000110011000101010000010000010110111100011;
#1 $display("%b", po);
# 1  pi=207'b110100001100010111001111011000111100101001001110101001110001000101101011101101100011100110111001000101001111101011110100100111100110100101110010111101011101111110110001100110011000010101101100111100001000101;
#1 $display("%b", po);
# 1  pi=207'b000111101001101010110011100010110111101100010100110011010011110100001000100011011011010010001110100010110100001000000101011110100101010011111100010010110110101101100100011111011000110101110000011101010110111;
#1 $display("%b", po);
# 1  pi=207'b011000001110110110101100111000010010001101101110100110001011001110110000001000110101111110011011101011010111010101101100010010100000010110011001001110111101011101111000100100110001110001000010011011101011101;
#1 $display("%b", po);
# 1  pi=207'b001101000000111001111011000100000110100111110110111000110001011010100010111110000010110001101000000101110001100000111010011101000011100111000010011100111110100111100101011001111000111100100101111011111011000;
#1 $display("%b", po);
# 1  pi=207'b100101011111010010101011111100001111101111101111010101000101010001111111110111011111100001110101100011001100011100101111000101110010001010110001111010101011001000101010100101011101000111110101101110101001011;
#1 $display("%b", po);
# 1  pi=207'b110000001111000001101000001100001001111100010100001101101101100100000001001000001000111101101000101010101010000000001001011101000010011000101010111011001100100000010011001011111100011100101111001000110000000;
#1 $display("%b", po);
# 1  pi=207'b010101011011001001001110111100101100000111110011100001010101011001111010001001011111111100010111010001100110000100100010011110111010010110010101101100010100011000001110011110000101000110010001101101110110010;
#1 $display("%b", po);
# 1  pi=207'b111010011101101010000011111110101000011001000000000111101010100011010111101011001001001110000111110111110100101100010100110101010010100101101000111111110100100110010001101111111010001011011101100110100001111;
#1 $display("%b", po);
# 1  pi=207'b101001011101101100011111101000011000101000010100101101011000000111101000100001111100101000110111111101111101001001110010100100111111110100000001110010011010010001111001110110011100110000010111001001100011001;
#1 $display("%b", po);
# 1  pi=207'b110100110000000010100010100010110011011111010101100100001001111000110000100000111100001000100101100110110101101000111010111111110000100101010011101000010111101110001001110011100100101001010010101010101010001;
#1 $display("%b", po);
# 1  pi=207'b100100100111000001000110111110000111101000011100010001110111100010111000111101000001010100110000100001011000110100010110000000110110111001100110000011010100100001010110100010011000100111110010110100111010010;
#1 $display("%b", po);
# 1  pi=207'b010001101110011001100001100010011111001010011110111100011101110001011001100010001010100010000000001100011001011011000111001000110010010000111010001010111001010111010111111001110001110101011110001000011100101;
#1 $display("%b", po);
# 1  pi=207'b001111100100011001000011110000111110111001100100100111000111100100110001101011101001000000010101111001011100101100110010110010001000111111011001110111100000011111100101100110000001001000101111001100111001010;
#1 $display("%b", po);
# 1  pi=207'b000010101110111010001111000101000100010010000111001000001110010000101011010011110001110101110001100101111010111101000111111011000100011110001101101111010110011000110000000101111110100000010000001111000000110;
#1 $display("%b", po);
# 1  pi=207'b001000011100011010111011101111110101101110111011101010000001000010001101100000100011000100000011111100110101001000001100111011010111110100111011110111011101111101001010001000111001010101001010010010001101100;
#1 $display("%b", po);
# 1  pi=207'b100110001001111100001011110000011100010000011110111100000100110101000000100110010100011101101100111011001100000111001000110001101111010111001110000110001010011111100011001001010010001111011000000010100011110;
#1 $display("%b", po);
# 1  pi=207'b001111000110100010001100000001111000001001001110010110101111111011001000110111001100011111100000000110111000000011010010111000101000110100110011110110000001010101010010000111110111101101010000100011001110011;
#1 $display("%b", po);
# 1  pi=207'b011000011010001101101110001000011110100111101010111000000000111011111000111111001111001100100101100111111100000101010010010100001000111001001000111001110010001010111001111001100011011101011110000011101100010;
#1 $display("%b", po);
# 1  pi=207'b111011110110011010111111111101000111111110100100110101010010110010111011101001101110011111100010011100001100101011010101110001010001100000110000110010010110011101010011010110000010111111111010010000011111011;
#1 $display("%b", po);
# 1  pi=207'b010011110011100010001101110001010010111101101111111111001010010111101111100001001010110110010010010001101111000110100001100111110011011111010010101101111100111000011001100010100110101000011100100001110111110;
#1 $display("%b", po);
# 1  pi=207'b110110101010010000111000100110101011011101111111101001001010001101110011101100101111000100000010001011001010001110000000001001110011100110011001010010110110101010010100101101110010011000100000111110111001011;
#1 $display("%b", po);
# 1  pi=207'b100110111101100101100001000010111101010011110100111011110101111011110101011010010001100000010111011111001111010010110110001010001001011001100010100011010001011101000110111011111110010110110101010111010011011;
#1 $display("%b", po);
# 1  pi=207'b010111100001101001101111100100101011000010110111101010100001111111101110011000110000000111000011001101111100110110100010011110110000100011001110000000111101011111000010010000100110011011111101011100101000000;
#1 $display("%b", po);
# 1  pi=207'b110111011001101000001111111101001111000111001111011000111001111001011011111111101100000111001001111110001010110111000111111110100010011010101111101001000101001101111100111000101111111001010011010010011010001;
#1 $display("%b", po);
# 1  pi=207'b000110100101111101111100001000001011111001101100100011100111100010011010110111100010011010011110010101101100110111100001010000010110010001110111011010100101111010100100010110111011100010000010010001111111101;
#1 $display("%b", po);
# 1  pi=207'b111010010010111111000001011010100111000010110110101110111110110110010001000110110101100110110001010011111101001001010011101111001010000010010010011000011000110001011001011000101101001001110100000000010100100;
#1 $display("%b", po);
# 1  pi=207'b000111001101111101101110110011101111010110000001001011111111000010101011011110100010010010010111001100100000000011100111011001001001101100011010101010010111010100011111001111101010101011101101110000110111101;
#1 $display("%b", po);
# 1  pi=207'b011111000110001110110010011110111000100010000101111000010111101100101100000101011110110010111111010110000110001001011110101101011111000010111000100111100000011011101010001101000101001010111100110011100011010;
#1 $display("%b", po);
# 1  pi=207'b010010011101101000010110100011000110100101010000111100010101001101100100010011010101111111001001010001000010101000000101100101100110010111111000000100000110111100010101011100110011011010100110111010100110110;
#1 $display("%b", po);
# 1  pi=207'b111101000000010100101100111111100101110101110110110000100011011010111111001101000011001000000010011000010110101100000010100101001111010110000110111010110001000101001010011001000001111001100110101010111001010;
#1 $display("%b", po);
# 1  pi=207'b001011010110000110010001011101001000110111101010110101010111000000100010000001010100100101100101010110101000010000010111110011100111010001100010100001111110011011101110110001110000100111010010100110101100111;
#1 $display("%b", po);
# 1  pi=207'b010011010010011110111010011110001011001110011001101101111000110010110111100101110111001010110001010100010011111100111010110111010101110001100010000100001000001111000100101111000111011000110010100100101010000;
#1 $display("%b", po);
# 1  pi=207'b111100100100010000001100110111000010010011000101111001011011000000111111001010110100100110100010000100000101000101010101110101100010110111100011110001001010110110100101001111001100101100100110001000111100110;
#1 $display("%b", po);
# 1  pi=207'b111011001100001010100111010000111110010011101011000101100111011011010111011010011010000001111011101110011011111000101011101010000000111000011000000011110001001111101110101010111001001101100001011001111101101;
#1 $display("%b", po);
# 1  pi=207'b001010100101000011110111010100100011100011001111101101110110100110011111011001100100111111011010011001000111001001101000001100010101100111000111110010101001000111000101101011001111000011101011110100110101100;
#1 $display("%b", po);
# 1  pi=207'b011011111111001000011011011111111010010111111100111001000000100010000110110100010100011111011110001010000100110110100000111001011101010011000001101110110100010100001101000111110101011010100010000100010111100;
#1 $display("%b", po);
# 1  pi=207'b000000111111100100110000111100000111111011101010000101001011000101010110100000001100101101011010001100010000010010100010110010110000100010101111111111111100110110010010001100010011100000111100000001110000000;
#1 $display("%b", po);
# 1  pi=207'b011000100000010010110000000110000110011000011110000011000011000100100101100101010010111010010101111110011010111010101000101000110001110101100011001010001011000011101111101110000111001110111000001011010001110;
#1 $display("%b", po);
# 1  pi=207'b000111000111110100101000101010101010001111000010100000101001111101010000000001001010110010101001111001110000110011101001101011011001110010000011110100111110000111100111110101011011000111001001111011001110001;
#1 $display("%b", po);
# 1  pi=207'b011111010100100011000100001011101100000111001011101010111101001111101111110001001000000000010110100111110000111010000110101101001100000101110011011001000111101111000001011001001011111011110011001100011001111;
#1 $display("%b", po);
# 1  pi=207'b010011010111010100110101010110010101100111010010100110011011100000111001010010011011011110001101101011011010111110000111011101100111100101110101100101110001000101100000100100111000111010000010101000001011010;
#1 $display("%b", po);
# 1  pi=207'b011011111000010011100001000110110110011101011101110001010101100100101010101001001000101001100001010100110001110001010111011110101000001001001101111000011010110011010101101111100000011011111001010101010011111;
#1 $display("%b", po);
# 1  pi=207'b001001001001101011110100001100001010110101000011111111011100001100011101010101011000011111011101001101111000110110010001110110110010111111100110010110111010101111011111011010001011110111010110010010010101010;
#1 $display("%b", po);
# 1  pi=207'b111000101001100101101110011110111011100111011001111100011100011000011000100001001110000011001001001000110011010001110101001001000001001101010101011001100100011100101011001110000110101100011111010001001000000;
#1 $display("%b", po);
# 1  pi=207'b011001011001000111101100010011011111001110010110010110111110110011000110111101010001011100101001010011001100110001000011110100110110110100011100101001100110101100001000100011101110101110100010110110100100001;
#1 $display("%b", po);
# 1  pi=207'b100110011000100110100011111100111000111100111001111111111101000111101010110001000111001011111111000110001101101011100001001111111110111101100001101101111011111101001111011000100110001000111001001011011100101;
#1 $display("%b", po);
# 1  pi=207'b111001110000111110011100010010010011110000111100111000110000101011101111001100001011111111101011110001000111100101000111111110011110001110001100000101110101011011010000010100001010010010110110001110000000010;
#1 $display("%b", po);
# 1  pi=207'b001010010010011000000111110000100101011000100000011010111010101010100111010100011010011110010000001100000001101010110101101000001000000000010101000101010010101001011001010101110100100110101011101010111000110;
#1 $display("%b", po);
# 1  pi=207'b100001101000011110111001000010101010011011111011010111101100000100101111011000100001110100100100101011110100100100111010001100000100110010011011110100110010110110101000000101111000100000101011001000011111000;
#1 $display("%b", po);
# 1  pi=207'b001011110000110100000100011010011101001001111110101000101101001010011001100010101010111111000000001111001000010111011100001001110011001110110001101001000111100110000111001110101101110000011011100011100111010;
#1 $display("%b", po);
# 1  pi=207'b100010100011101011001010101000011010100010001000110110010011001110011010110110011100110001110000110001101110011011111100011000101110100010001100001101011001111101001100001010100110100011110100011110111001110;
#1 $display("%b", po);
# 1  pi=207'b100010101001100101111000010101101100010101011001101101101111011110100100011111111110110000110001101101000011110111011011011101110101010101110101101001011100010110101010010100111011001010011101010010011001010;
#1 $display("%b", po);
# 1  pi=207'b001000001110111110000110011011011010001111000101001010100100111111101100001001010111100000101111111010010111001001011011000100000010100010001111000000110010010010110110110111110100011011010101100001101001111;
#1 $display("%b", po);
# 1  pi=207'b000001010110111111101101111010101110000110101001111001001101011001001101010010011100100000011111001001111001011001101100000111110001101011101110111011011000010001110110100111111111111000100001101101111000110;
#1 $display("%b", po);
# 1  pi=207'b111000010011000110100010011001011001010000011100100101100111101101001110101110001011000101111110010101011100000101100111000100001001000100010110101000011111001101010010010011000010010111100110010001001111100;
#1 $display("%b", po);
# 1  pi=207'b011110001111100001100100010100010110110001000100101001110001111101000101110101111101000100001111100011100000011110111011110000100001111110110110101001110100011111000110100111010001101110111110001101010010111;
#1 $display("%b", po);
# 1  pi=207'b010101110100110000111110011110011111010111010110010010000011101001000111101110001010100000111111011100010001010011001111101000101101101000011111010101100001110100111110101100111101100001100001011100110001000;
#1 $display("%b", po);
# 1  pi=207'b111110001100101111010100111001101111101111100011110101111001101100000011011000100011111110001111101100001110001100011011110111101001111000110110101100100110000010010000111101110001111100100101111101010111000;
#1 $display("%b", po);
# 1  pi=207'b011111011000011100001000101010110111110111110001110111101110010001000011000010010011010111100110001011010110111111111000001001000010011101100000111011100101001100000001001101101001110101010110101010110111001;
#1 $display("%b", po);
# 1  pi=207'b000100000100110011001010001001011010110100000011001011100100001010101001110110100110010110000110101010100100110111111010011100011110100010111101111101000000000001101111101110000110100011000001001101010001111;
#1 $display("%b", po);
# 1  pi=207'b011011110010100011101000111010101110111100000000010001011101011000011110001111101000110100110111111101101000010000111001011011100001100101101111110000001001100001100000011100101011010101101010011010001010011;
#1 $display("%b", po);
# 1  pi=207'b100111101111111011101110110001110101000001011101101000111011101101001011110101010111100101110101000100101110010101011001000100101010011001101111101111100001110010100001101010010101111111000010100000111111100;
#1 $display("%b", po);
# 1  pi=207'b001010010010100010110011010100100100101110010001100011100100000010011100101001110101111101000011101001101010110101101100111011011101011011110111000001111001010000111010000110011111010000101110111101100111011;
#1 $display("%b", po);
# 1  pi=207'b010110001010101000011111110101100111100100001100000110110101000011010100100011000100011000111101010100111100100000011111110010110010100001101101100111101000100011011111110100101101001110000010000100111101000;
#1 $display("%b", po);
# 1  pi=207'b000001100111010101010101011101101100010001110011010001101011000100110101001011001001011011001001011000111100000000100010101010111001100010000011111101000010001111001110100000011011100001011011100000101011001;
#1 $display("%b", po);
# 1  pi=207'b101111001100110100001000001010001101100100010110110110011000110101100100000010111101000010110110010100100010111111101110011000010011111000101010110011110111110101100110111000111011100111011101110101110010001;
#1 $display("%b", po);
# 1  pi=207'b001110110001101100111000100110111100101011111000011111000110111010111010111100010101001111001011101111000010100000010011100001111110100011001110100100111110000001000111100101101001010000010000011010111110011;
#1 $display("%b", po);
# 1  pi=207'b101111101100100001001100111001101000010110001011000000000111110011011101100011100100010010010001110001001001101100001011110010101100010100101110100100111011111010001110000100110011011001000001100100101001001;
#1 $display("%b", po);
# 1  pi=207'b111010011111001111100000010100110010110111111110111111100001111011000011110101000100011000101001101000110111011010110111110010010011001100110000000110000001011011101101111011011101100011011101001001010101101;
#1 $display("%b", po);
# 1  pi=207'b010000111001100011101100111101101001010000110011111000010000111010010111000011011111110001111110010111100010000011110011110111000100011010000010110011101100000001000001111010101011001111100110111010101100101;
#1 $display("%b", po);
# 1  pi=207'b001000010101110111011100000101110011011001111100111101101000101111100101011001001010011010101110110000010011100010010110101010010111010001000001100011000000100101000100101011011110101010100111100010010101011;
#1 $display("%b", po);
# 1  pi=207'b001000111111101100100110111100100000111000100010000001000101101010001111001010111000101101101001101001110110111011010101110111001100001001100100101101111011111101001100001000011000110001101100100110110111111;
#1 $display("%b", po);
# 1  pi=207'b101000000011100001111101011100001011111001011100100001111010100110000001010110001001010001011111001111110101011110001100010100000100110001111010101100100000111011000011110010001000001011100011100010111100011;
#1 $display("%b", po);
# 1  pi=207'b110111100011011011110111000001111011100100101000111011101000001001101000101101100000000110110011101011110100111111110011000001001001000100011110111001000001010100010000101111000101110110000011010100101000011;
#1 $display("%b", po);
# 1  pi=207'b110011101110000110010110101010100101001001111010110111101001001110100011100111010001000110000010001100010000011110000111100101001001110010010011100110100111110001111101010110001001011100111111011111011011011;
#1 $display("%b", po);
# 1  pi=207'b110010110001111100001100111101100101101011011100000101110000000101011110101111101000111101101001011010100010110000110011101001101110000000010100000101010000110000011010000001101110101101100100000111010110101;
#1 $display("%b", po);
# 1  pi=207'b010011000101001001010100010110000111100001101011110110111100001001010011010100101110100001011010101111000100100111001010101101101011010101010001001000000000010011100011111010011010011010000101111000000101100;
#1 $display("%b", po);
# 1  pi=207'b111111011000100110101111001000110111010011011111100010000001000110011001101010001100000100000101001110100010101110110111010000110000001000010011010000011000000100101100000101001000100011001010000011100110100;
#1 $display("%b", po);
# 1  pi=207'b010001101111101011100010100110000000101111011100101011001011000001000000110011100111100000100110101000011001001000000000001111000000000111100000001100001011001110010101110111011001110010110000010010001001010;
#1 $display("%b", po);
# 1  pi=207'b100010011111100000010010001111011001011101001101000111011111011011010110001101111001110001100100111001101011101010011000010100110011101100100101011111111010101100101011000111111101100101010010001100001000100;
#1 $display("%b", po);
# 1  pi=207'b111100111100010000110101001110010011001101111010001101110011100011111000011101100100111001011110000001110000100000010100101010111001111000100000000011011110001111001000101011000011100001010000100100100100110;
#1 $display("%b", po);
# 1  pi=207'b110011100001001010100011100000001000010101000010011101010101011110011011010101010111001100010100010001100011111011100010001000010110100000010111100100011010111000111001100011111111001100011001100100001111110;
#1 $display("%b", po);
# 1  pi=207'b101100001100000101101010001011111011110011111001010000010001111011110000000110111001000001011110000111101001000000001111000101011010000011011000111011001110110101101000101110000100101001010010011111110011011;
#1 $display("%b", po);
# 1  pi=207'b010100000000100111011100100101100011000001110100000101011010001000100111010110111111010000010111110011011011011011110101100011010100001010111110101100100111001001110001100110000101101011011101101011111110100;
#1 $display("%b", po);
# 1  pi=207'b000111101101110001010111111100001100110011000110011101011101000010100000100011011100100100101001000001101001000111001001101111101110101111101111100101000101110101011100111110111000010110100010011001111101111;
#1 $display("%b", po);
# 1  pi=207'b001111010110001101011001011100001001101110001111001111110011010001001100011101110101110110100110011100110010101110111110011001010001010110000100000111001001110110000110100111000111100100100110011111101011011;
#1 $display("%b", po);
# 1  pi=207'b110111101000100001000110010010011000000110011110011011100000111001100111101110000000000011000100010101011110010100111110100010101100010110000011010011100110111111000110110111010110000001011001000010001010011;
#1 $display("%b", po);
# 1  pi=207'b000100110000001101010001001110010100001100111110111101000010100110011010011111111111101110001101011100111001110011101001110100101010010101111000111110010000111111000011111000101001011000011110111010100010000;
#1 $display("%b", po);
# 1  pi=207'b010100000111010101010100011111010010110010011001101011011101110111101010011011001101000111000001011110011111010000101011101011011101001111110010001011011100110000001100010011111010011110001001011000110111000;
#1 $display("%b", po);
# 1  pi=207'b000011100100100111111111000010011000101111010011001100111001011011000000000111110111100100111100010111000100011101010110110100001010110110100111010011101100011101001000011100001001010101001110011101001101011;
#1 $display("%b", po);
# 1  pi=207'b001001100011010001001000110101010101100100100111100100001011010000010111101001100001110001010011010101000101010111011000010100111110010010101101011111101101001100001000111111111101100011010000101011100101101;
#1 $display("%b", po);
# 1  pi=207'b001101110110101110001011011100110010111100110101000111100000100101111011110011110110000110010011101000111100010101001010000110001001101111010110001100110000011110110000010111100110101001011011001110011001100;
#1 $display("%b", po);
# 1  pi=207'b001011110001011001111100000110001001110110001111110001101111101100010111111101101111001000110011100100010100111100100011110110110000011100111010101111100101110100011000000100101011100010001001101000111101010;
#1 $display("%b", po);
# 1  pi=207'b110101011001110001100010110111101101111011101100100000011000011001011001011110101101111101100011101011010110111010111111001001000001111110100010011110111000010010011001101110100011101101101100111110100111101;
#1 $display("%b", po);
# 1  pi=207'b111000001001000110101110000010101001001011110000011100010111010111110011010101011101101000010111111000001100000111011010001011010110001001111011100001001011011000000000010001000101011011111111110110100110111;
#1 $display("%b", po);
# 1  pi=207'b101100111000000001100110001110110100000101011010110110011010001000011111001101100000011101011011100011011101001100001010010010011100101001101110111100001000100001111110100000101101111111100101101101011100111;
#1 $display("%b", po);
# 1  pi=207'b110010101000101011000010100000100010110000001001000011100001101101111011101001111010001100101001001001110010010001001001101111010001011110001111100111100100011101110110010100100010110100101111001100001110110;
#1 $display("%b", po);
# 1  pi=207'b010100110010000101100000010000011010110101101100100110100010010101000110100001111011011000110100010101110110011001100011110100100110101010001001001110101010100001011011000111110010110101000001001000000010111;
#1 $display("%b", po);
# 1  pi=207'b011011111100110011001010110100011001001010010100001010010000111110111101111111111000111100010011111001011100010101110010011101111000101000101001010100001111011111100001101011000001010110010011010001010111000;
#1 $display("%b", po);
# 1  pi=207'b111001000000111010110000101111100100110001001010000011000010111101011000010111110000010110010100011111010100101000011001001000100111000110010011101100101001110100101000011111111111011111000110110001101101110;
#1 $display("%b", po);
# 1  pi=207'b100001110001100010100001000111111110100101101110001011011000011010000101010011100111101000100010011011111000101011111001110101100100010010110111001010100001111001011111000110100110000100011110000000111010001;
#1 $display("%b", po);
# 1  pi=207'b100010010100100110011100101111000101010000111011111011110010001010110000110110111101011011101101001101100011100101111101010010001011001011110111001010101101000001000010011010111000000000001011111000011010011;
#1 $display("%b", po);
# 1  pi=207'b001100101101010001000010010010111011000111000100100111010110010110001011000000111100011110100000100000011110111110100001001010110000101011111111100111000111100101110110001001000010100101110100011001010000010;
#1 $display("%b", po);
# 1  pi=207'b001000011110010101101010110011100011011100010100001000011101101011111101100000001111011110111001101000001110111000011001100011110111001100011101001011000000110010110101111010000000110011111111001010101010101;
#1 $display("%b", po);
# 1  pi=207'b110001010110001010000000101101110010011010110011110110111011001110101010101000111111001111111011010011001101110001010110101011110100110011011011000101100111110011100010010100001001000100110101001011000101011;
#1 $display("%b", po);
# 1  pi=207'b101100000011111001110010001101110110010101000100111011010000011101110101000111110000100000100101101111011110011011000101001010111000010001010001111101001101111101011100101000101011110100001100010010000011100;
#1 $display("%b", po);
# 1  pi=207'b100100011001001101011110100000101011000101011000101110101101001111100110000001011111100011110000010101010110000000001010100001011011011000100011011000011000000000011110100111101001011001110101100000101001010;
#1 $display("%b", po);
# 1  pi=207'b010101110110111100111110000000100101011101000101010111011101001000011000111000010001010000111001100011000011000011100100100011000101100001001001100010111010100000011111010001000000000011000000100110001111100;
#1 $display("%b", po);
# 1  pi=207'b010100101100101111001100001110101010010011100100101101110001010010101111110101101100000111011011100000011100011000011010111000110100100100000101110111011110101110001001000001010010100110010001111001010101101;
#1 $display("%b", po);
# 1  pi=207'b111001011001000011010101000000111011100000110010001001101010000000101110011000100110100001010010110000101000111110011010110011101011111010110001101000011000110011100001100011111101001000001111001000011101000;
#1 $display("%b", po);
# 1  pi=207'b010011001101111101100100111011100111101010000110011101101011010110111010100001011111110001010001101111001000001101001100110000010111001101010000000101011001111001110100011110100011110101011101111011000001111;
#1 $display("%b", po);
# 1  pi=207'b000010011101111101011100101110110001001010000101001001000000101000011100000110010010000000110011000100101111010010000100110001011011000100000100100001111001111001110100111000101111011000110010110010000101110;
#1 $display("%b", po);
# 1  pi=207'b110000001011101101101110010010010100100000100010010101101001001010100011100010011100011101001011110001110111111000110001110000110000001010101000111000110001110100001110011001000111001100100000101100101011000;
#1 $display("%b", po);
# 1  pi=207'b011100110011001000111110110011100000000011001100001110010110101111100010010011100011110001101100111001110101100101000011011101000011100011010110100011110000100000110110100001100100011000110011001110000101101;
#1 $display("%b", po);
# 1  pi=207'b011010001110110000010100010100101110000111111100110000111110101001110110001000001100101001111110010111001001011001100110000110011100100111011001101011010010010111000010110110100010100011111101011110000110101;
#1 $display("%b", po);
# 1  pi=207'b101100111101110101011000010101001000000111001010100110101011011101010010111000110110011110000101110001101010010000111011000110100111110000011110110110101000110000100000001001110011111000011101001000110011101;
#1 $display("%b", po);
# 1  pi=207'b011110000010011001101011001000110101111110011110110100101101101011000001000011001010101100111110111010111001000011100101111001010000111110110010111011000111011010111100011110101110101110110000110110111100101;
#1 $display("%b", po);
# 1  pi=207'b111010111100000110001010011010000101001100000100100000010101101110101111100110111110110110100010110110011000011100011100001111000000101101000111001101001101101101011011111000011010110011110011010011000110100;
#1 $display("%b", po);
# 1  pi=207'b110111101001010001011100001100111101111000110110101001010010010011001011100111100001000111100101011011010111011010010010011011010011101010010000111010010111010101101111011010011101110000010110100000001110100;
#1 $display("%b", po);
# 1  pi=207'b101110011010001010010011001101111100011000011101000100000001101110000111100000000000010101001000111000001101101001000100110001000011000011000001111101000111001111001000110000001000100100110110001000100101001;
#1 $display("%b", po);
# 1  pi=207'b001011101010110100101011011011110110010001010001111001111100110011111110100101100111001011101010010111000110110101010011011110111100010001010011101111101011000110111001100111011110000010100111101111110011011;
#1 $display("%b", po);
# 1  pi=207'b111101001100111011011001101111000101010000111000111011010010000111110010101101100001000000101001001100110011010111101100110111010000110100011011001000001000000101010111111100011010111100011111110100001011011;
#1 $display("%b", po);
# 1  pi=207'b000001111101011110000111100111010101001111010001110010000111000010111100111111001111001011011101111011000010110100000111001011010010111011011001100110100110100000101010100111111110011100110110000010001010000;
#1 $display("%b", po);
# 1  pi=207'b101110110110011100110111100000001111110110010011011111010010110001001111110100101100111110010001000010101010101111110001110001000001101101010011010111111100000111010101110010001100000011001100100010000110100;
#1 $display("%b", po);
# 1  pi=207'b110101011110010111110111101000101010101000110010111000100010100000000000111101000011010111101001000111100001010000100111110001010001000001100000101010111110111011110110101010000110100011100011010110111111001;
#1 $display("%b", po);
# 1  pi=207'b110000011111111011101001010011011011011110100011001111100010100100110011100110101101000001010100010011110011001001100001000010100011010111111111000001010101110101001011001011001101110000111000110100110100001;
#1 $display("%b", po);
# 1  pi=207'b001011101111101110100010111001011100101000111001001110111100101111111001011100101011011101110000111111100110000111011001100110100011101111111100000001110111001010110000010010100010000010011101000111001010101;
#1 $display("%b", po);
# 1  pi=207'b100111001000001110001111110100010101010101111011011101001010110000111000100100101001111010010010010011111101101000000100100100111111000100100000001011010010011010110110001010111011101111011000011001111111110;
#1 $display("%b", po);
# 1  pi=207'b110101100000001111000010101001111011100100001111110100110101000000011100110111000110110101000100110010011101011000010001011011111110100010100111110011101010001111010100111111101001011010111100101000110000101;
#1 $display("%b", po);
# 1  pi=207'b000010001100000100110111110011000000010111010010100000001001000010010001101111011010011000010101101100010101100100100111110100100111111100100111011110011000100100110000101000111001110011011101000111000101011;
#1 $display("%b", po);
# 1  pi=207'b011110010001101111001010011011010010011111101001010001101010110010111100001111001101001111000100000110010100110000111100110011101110000100010110010000011100110011010010101001100010100000100111100001100101010;
#1 $display("%b", po);
# 1  pi=207'b111111100110100101101110101110111011100101101001011000001011000100000011110011010101101100110011010010100110110011111111111011110110100010110001110101100101010100110101010111001010011101010011110000111100111;
#1 $display("%b", po);
# 1  pi=207'b000010101100000000011110101101111100000100011110101111111110100010111011100110011010111101110100110111001000110111000000000111000101000001100111101111011011111001011001010111110110001110000101001110110100101;
#1 $display("%b", po);
# 1  pi=207'b100110001010000111001100001111011110001101011101100101110011100101110110111000100101110011010100101110110101011100111101110001110000011011111100110101001010110111111011011011010011011010111001111001110110011;
#1 $display("%b", po);
# 1  pi=207'b010001100001011110101100011110011111011101110011011000010111010111111001101110011001100101100111010110101110101110010010011000101010100101001000100110010101101100001100011000000000000010011001001010010011110;
#1 $display("%b", po);
# 1  pi=207'b001111101101001110110110101000111111101001011111001101111010001001010110001000000111111111000011111111100000000010001011101010100101101110010111011100100101011101000010101010110011110100010100110110110000110;
#1 $display("%b", po);
# 1  pi=207'b111101110101010000010100101000011000000010101100110110100110010010000001011011011001100010111110100100011001000001000110001110011000010011100100010110011110000011010001110000011101000011001110001111111110011;
#1 $display("%b", po);
# 1  pi=207'b011001110000000110000011101110101011111010000000011010100100100101010100001001110101000101010100100000111011001100001101110101011111101100010001101000001011101111111000111110100101100010110001110111000010001;
#1 $display("%b", po);
# 1  pi=207'b011100000101101001101001110100011110100010011011110010111001001010011010001000110010010110111101111000011110100111111011010100101100011000001001110101110010010011011111000001011101000010001111111110000100111;
#1 $display("%b", po);
# 1  pi=207'b100010101000001100000011000010001000010110100000110110111111001000110010101110010010110001000010110010111000100111100011011000110001100111001110011001110101111101110011111101100011000011001011000001001000000;
#1 $display("%b", po);
# 1  pi=207'b000100000000011101000110000001100101111110100000011000001001010000000001101001010001001011011011001010011000010010101011010110000001001101100000011101111001101011111100101100000110110110100011110100001110011;
#1 $display("%b", po);
# 1  pi=207'b001000000010110010000101110011011010100111010101000001001001010010111100011001010001011101111001001010101101001010110011100100101101000111000011011101010111100010110010011001011010010110111010111000100001110;
#1 $display("%b", po);
# 1  pi=207'b110110011001110101011011111111000001001010010101100111010110001100001110000111100001100110000001010110110000100011000100110100111101010111111100111011110111011101000000101001111100101011011101110001001000110;
#1 $display("%b", po);
# 1  pi=207'b000110001101010111001011101111001011010001100001111011000100101000010001111010100100011110011101110010011001101101010110011010011010111010110111010000010111110111110101111110010010100011001100010101010000000;
#1 $display("%b", po);
# 1  pi=207'b100100011001000110110100100110010100111101011111100111111001000110010110000000100011000000010000110111000101011000110010101111010001001100110000101101100111110101010111000110001010011011011111000111101010100;
#1 $display("%b", po);
# 1  pi=207'b011111111101110001000111111101100010110001101100110001001101101100001100010100011011000100010111011101101001111001000100111100010001011010001101100110010100110001111011000110001001001011011010100100100101111;
#1 $display("%b", po);
# 1  pi=207'b110110100001001000111000101101000001100110000000111011010001000110011110110110100010011001011010000110111100010011000101011101111111001010100110101001110101011110111101000000111000100111100000001111100011011;
#1 $display("%b", po);
# 1  pi=207'b111111111110110011000110101101011000100010110110001010111000010001101010100101001100010000000000101001100001000111111111111110001100111111101000010001101100101011101100001010111100110010010101000111101011011;
#1 $display("%b", po);
# 1  pi=207'b111101011111000001000111000101010000111111010001110111110010010101101111100100010101010111001001001101111100011111111110000000011000001100001011000001100001101100011001010010101011000101000101110100010111110;
#1 $display("%b", po);
# 1  pi=207'b100101011101000001100010101111000011011110101011000001110111110011101100011010110111001101101011100101011011101111110001110000011000111011011010000010010110110011101011001010001101101100110111010110100011000;
#1 $display("%b", po);
# 1  pi=207'b111110100101000110111010101101000000110001101100101000100101001010111011111101011110000010110111110100111010011100001000111110101001101001101101111010101011110110101111001011100110000101111001101001010011100;
#1 $display("%b", po);
# 1  pi=207'b000110110000011101110011001000110100101010100110110010111110000100110010100110100001011100011111111111001001011010001001100111111101000101110110101000111100000001101111110100101110111001101100010011011011101;
#1 $display("%b", po);
# 1  pi=207'b111111101000011011110011011100001101010001011001000000110000111110110010011110110101010010010000000011011000011000110000001110001010010101011000100101001000111010011011100101111111111010101111100111111010111;
#1 $display("%b", po);
# 1  pi=207'b110100111110001100111111001000100100100001010100110001110110111010111110000011110110011101000100111111101001011001111101001100111001010001001000101101110010101101111011100100011110111001010010000110010110010;
#1 $display("%b", po);
# 1  pi=207'b101101110010000100010001100011000111100011000110110001000010001100101101001101001111110101000011110110101011001010101001110000101101000001011111001101010101101001110100010010111100001101100101000011001111011;
#1 $display("%b", po);
# 1  pi=207'b011011000100010001101001100010011110001101101100011001100010111000101111000101001000010001110100111111111110100101010010100100010101011001000010000110110101101001101101110000001111111100011011011110010000100;
#1 $display("%b", po);
# 1  pi=207'b111011000111011000100011100110001010001001010101010111111110100010111000000011011011100110110110100101110101001100101101010101111010010001110100011111010111011111110110011100001010111001001001011011110110100;
#1 $display("%b", po);
# 1  pi=207'b100110111111001100111001011000101010110110111010111001100000110001110101100110000101011101011001011011111001111011000111110000011001100001000011011100000011010111100010101101001100001000100111111111001001010;
#1 $display("%b", po);
# 1  pi=207'b110000111001000100111101111001001011011101011001011000101111000111101101001101011001100001001100011100101011101011101010100011111010010110100100101110011110010001100001101110101010100111011111111010001010100;
#1 $display("%b", po);
# 1  pi=207'b001010011111100100111001100010001001110101101111010001100101111000011111001111111110101101001100010001010111110010001100101011110001100011110110111011110100110111100011011111100100111101101110001110111101111;
#1 $display("%b", po);
# 1  pi=207'b100011101010111100100111001110010011110100101000110000101110111110011110111001000011101011011110111101111101010101110011001111111110101010110100110100110100111111001111010101111011000110001001010111000011101;
#1 $display("%b", po);
# 1  pi=207'b001110110111101010000110011111111011011001011100101000111001110100011101111110010010010110011001110100001000110101110010001111111101101011100010010100000111000110001101101011101010001101110010011111000111000;
#1 $display("%b", po);
# 1  pi=207'b100111100100110100010110100011001101100001111001010111000110100110010110101010011100001001001001000010000111000011111000011101101011001111101011111100100000001010011011001001011010011000000111110001001000011;
#1 $display("%b", po);
# 1  pi=207'b010011111001100100111011110001000001000110000100110100111001111010010010011100011111110110101111110111101101100011010101010000001100101000011100001101100011011000100011101001100010111100111101010001001000100;
#1 $display("%b", po);
# 1  pi=207'b110010001011110001010101101010100111100010011011110100111000010001110100100011010010100111110100110010111000100011100001010001110001100101001101010001001010001101100000011001110010100001101111111000011011011;
#1 $display("%b", po);
# 1  pi=207'b010100111001111101101110101000110111111000000111001000111001001111010000001000011010110110110000000111010110001111100011001000011011001000010001010001010100001011001000010100001111101101011101000010111011011;
#1 $display("%b", po);
# 1  pi=207'b001110111000010001011011011110000000010010100000001011010110010101110101111111001011110011000001010010110011111011010001101101110100010001111101101101101110010101110100010101100010100110010010101101010011000;
#1 $display("%b", po);
# 1  pi=207'b000000011101001010000101100000100001111111010100000011000110001110011101100011000000110001111110100000111001101010001101001010001111001100011011000010100101101101100011010010110111111101111001001100111010110;
#1 $display("%b", po);
# 1  pi=207'b111011010110000100001110000010101101000010001101001010010000001101110111010100010001000111111110011101111111011100111001000011110111101001001011011000010100100111110101101111010101010011111000011101111110111;
#1 $display("%b", po);
# 1  pi=207'b001101010010000000001101101011011001111110100111001010000101110011100100100111111000100000011111001110000011101000001001110001110100100100000000101110111011100101001110111011010010010011110000000101100100011;
#1 $display("%b", po);
# 1  pi=207'b101111000010000001111001000001100100000011111111000001011010111011000100101011100010111000100101100011100110011001101111110001111110011000011000011010001100110010001101101111011000111010111000100001110100111;
#1 $display("%b", po);
# 1  pi=207'b011000010111110101010100001000010011110110101000010010100100001111111001001110101011001100001101010001001010001011010011011011100110111100110000101110101100001111100001011110010000101010001010101000100110001;
#1 $display("%b", po);
# 1  pi=207'b111111110010001011101111011001000110111101001011111101111000000000001111100010011001001110001110101010001010010000000010101001100101000100100001011100110101010100001010000101110110000110101010011010111000100;
#1 $display("%b", po);
# 1  pi=207'b001111011000001010100000010110011011111000110111101011000111101111011111010101101001111110010111001110010111101100010111000000011100000111001011101100011011101011011010000000101100100000110110010011111111101;
#1 $display("%b", po);
# 1  pi=207'b001110010001001111010111001000000011001000100011111111100100111111001000010110111111000111110001101100001110000001110000000101011110100101101110100000010110010010000100001110111010101011011111010111010110011;
#1 $display("%b", po);
# 1  pi=207'b010101010101010000000000101010110110010011101011111001101001011010011001110001010010001001100101100001000111111011111111110101010010101101101011001000000001001010111000000010011101111010001011110101011100111;
#1 $display("%b", po);
# 1  pi=207'b110001101010001000001111111011101011101011110110101101100100011010110001100010000011011010000001001111111011100111011101111011011001101000110110100100000111110110011000010100001100001110001010110101011000100;
#1 $display("%b", po);
# 1  pi=207'b101000100001011101100001001001101000000000100000010100110101100011000100101111101101111000110001001111001101011001101100000001001010111010011101011101101011111101100110110000111110011000001111101110101010010;
#1 $display("%b", po);
# 1  pi=207'b111111100111000101011111111100011110101010111001100000100110010011111010111001101011010011110010100100011110110000011010010001000111000010011100110101101111110111000001000100110110010110001100100111110000001;
#1 $display("%b", po);
# 1  pi=207'b100011111001011101110010011011010101100010100011010011001000111011101101000001001100111000011001000111101101011011001001011010100010111101010110100010011101110110001101000111000011010000111111111011101110110;
#1 $display("%b", po);
# 1  pi=207'b011111111011010111111000100100100011111011101110000011011101001000011001100010100010011110010001101011000001010111001011010010011111111101110101100011100010011110011011001000110110011110001110101010011111000;
#1 $display("%b", po);
# 1  pi=207'b000111111010110000001010011100100111100000001110100000101001001001100110011110110111000101000111100111111111010000101000111110010000100100111001100000010010010011100101000010110001010100101011111011101100011;
#1 $display("%b", po);
# 1  pi=207'b100111111001111011100011110100001001000110101111000001110110000001110001110110000110011111110100100111000000101001110101100111111111101110011110000010101111111110000011110110010011100111100111100001111100000;
#1 $display("%b", po);
# 1  pi=207'b101000100100101101011100101011100011100001011011101000000110001100010101000101011100001000010110100001100110101101011000101111110111101110110010010001100111100010111011000100011100000001010100101010100110101;
#1 $display("%b", po);
# 1  pi=207'b111111110100010000100100110001111001001101010100001100101001100110110010111000111110110010100111110010101001100001101110010001110000101001011010111010010001111000010100000000001001100001110101000110001011100;
#1 $display("%b", po);
# 1  pi=207'b110001010010101101100011110110101011110000000110001101110000101110011110011011111110110110011010011111100001011001001110001010110000111010011011110110000001100110111111010001100100100010101000101101101011011;
#1 $display("%b", po);
# 1  pi=207'b101000100011101100111001010010001000110001000100010101000111110011100100101000011010111000111000000110011110111010111100100100111110101000101101010110000010110001100011101101111100101101000001000100011111010;
#1 $display("%b", po);
# 1  pi=207'b010100001011010111110000011010111000101010001110011000010111010011000011110101111001000110111101011111000101011110111101010000110001010101001010111100000101000010000101100001001011011011101110100110001111110;
#1 $display("%b", po);
# 1  pi=207'b000100101100111011110101110100110001011011010001001001100011011101110100100100100101111111000110110010010001100010101001110000010111000111110010000000000100101001101100011011111100001001110011100111011001110;
#1 $display("%b", po);
# 1  pi=207'b000110010100111001010101010000110001001010110101010011100100010011000000101010111010101001010010011101001110001010110000000110010110100001011011110111101000010110111101101110010010000110011101010100111110110;
#1 $display("%b", po);
# 1  pi=207'b001010101100111000001010001011010010001000001000000011000111101001011001011000101011001011110001110101100000000110011111111001011011000011110111010101111000100111011100101001010110100100010011000101100000100;
#1 $display("%b", po);
# 1  pi=207'b011101001101110010011110111010101110100100001010101100001010011100110110111001010001110010010000110111001110010001011111000100101100011000110011000010110101100101110000011011001001001010000001000011000000001;
#1 $display("%b", po);
# 1  pi=207'b101010111110101110001111010001111100011111010100010010110101111000101110000111100111100011011101110110100111011100011001100101010101000110111100011010100100100001001001111011101010111101011000011011001111010;
#1 $display("%b", po);
# 1  pi=207'b110101101110110010001000100011011100011110011110000111110001100010110011011000011101010000110011111011110000000101111100110000101000110100011001001100010010111011010101111010000101111100110101011100000000110;
#1 $display("%b", po);
# 1  pi=207'b110000010000010001110010110111010000110111111101000100110101101101000001010101000110011000000010010011110010110101100000110110111001001010011101111101101110100111100101000001010100001101110011101100010000000;
#1 $display("%b", po);
# 1  pi=207'b000100110100001000110000100000101111101000110010001011101000010010010110101110101001110010110111000001110100011010010111100010111001000000000011110100000001010100000010001011010010110010011010110000011111010;
#1 $display("%b", po);
# 1  pi=207'b010101000011101000111111100001000000010000010010101100100000100000010010100101001110110100000101100111100110101000101110011011100111111100001110111010111010101001101101100000101100111100111110000111110010100;
#1 $display("%b", po);
# 1  pi=207'b010100010111110001011110000001111010011011010000011001011000110001001011000011100000011010011100100010101011011100001001101101111111011010111011110011011101010010110100100111110010101110000001110001100100111;
#1 $display("%b", po);
# 1  pi=207'b100101111001100100010000110110010001011101001001101010011011110101011110000101000000011111011001010010001001000000110011001101000011010110100001110110010100001001111101010111110000011110100001001000000011101;
#1 $display("%b", po);
# 1  pi=207'b111011001011111100001100100101011011101011111110101011000101100000110100110000001101010100000111000001001000011011100101100000101010111011100010000001100010100100011000111001101000100100001100101001001010100;
#1 $display("%b", po);
# 1  pi=207'b110110111110111010111111100111000110000000110001000101101011110100001111010110011000010000111011011010100111000010110110110101100011111000111000011110111100001010110100000100000010110111010110000001001111011;
#1 $display("%b", po);
# 1  pi=207'b110111110110011010110110101000001010000111001101111010000000011000111001001111101010100010001001101101110001110101101100001000011111010100110110011010111101101010111000001100010101011001110110010111011010101;
#1 $display("%b", po);
# 1  pi=207'b101010010101101011100010110010111101100010011101000100000111101110110001101000001110110101110100011101011010010100110110001101011110000001010110010000010110101000111001110011110010011110000110010110001100001;
#1 $display("%b", po);
# 1  pi=207'b000111010101101001111111001111110100111001101011010011110001011011011111111001110101101100001010001010000101000001001000011011000100010111100000101100010011010011010101011100000001000110100100000001111100000;
#1 $display("%b", po);
# 1  pi=207'b100011000010010110100000110111101101101101001101000111001001000100100011100001111101011111001010011010010111110010110011111001100001110000100100000101111001000001101000111001011100010000111110101000001110100;
#1 $display("%b", po);
# 1  pi=207'b011001010010000001101010010001011000010011101111100101010101010001111100111101111010110010011000110000011011111000000111111001100100010010110001001011000001111001000001011011011010001100000001101100011101010;
#1 $display("%b", po);
# 1  pi=207'b001111100111011011000111110110000110101101011000011010001001000001001010011100010101101001010011100011010111001110110110010001111000000000100010100110000100000011101001001000100100001101000100011000001100011;
#1 $display("%b", po);
# 1  pi=207'b011011101101101111010011100001100111000110011010110100000110000011110011110101110011010010000000010000111001001001000101101000110110101110100001110100111110010001111101101001001001110100011000100110011000100;
#1 $display("%b", po);
# 1  pi=207'b010101010111110100111001111010000011010000101011111111001010100100101010001000110100111101110001001110011110111000011110111111101001001101000100100111111001101101100101011001011110101001001011110000000000010;
#1 $display("%b", po);
# 1  pi=207'b010110001111010011011110011111100101011110011010111100011100011011100010010101100100010111111011010110110101010001010010110011110001110011111011111000000000011111010100011111000001100011000000001000110101010;
#1 $display("%b", po);
# 1  pi=207'b001011110100000111000100000001100111011010011011011000111110000110101001011100000011100101011100011011101010011101101011101101100100011010010011111011101000000011111011011110101111100101001001001101111101010;
#1 $display("%b", po);
# 1  pi=207'b010100111001001100111111101110111011000111110100110001110000110011001100101101110100100101101000001010011011110001100011100100101001000001001110001000000110101111110100001101011101001000101101011000001001000;
#1 $display("%b", po);
# 1  pi=207'b000101010010100100110011010011110001111110110011100100111010000100011111011011011010001110100011100101100111110011000100101110011101000101110100010100001111111001110101010111110100100010011000101110000000111;
#1 $display("%b", po);
# 1  pi=207'b100001110100011010111100011100000110101000001110111110001100000010001111110110001001111110000111011111100100111001100011100000100100010111010111100000001010010100001101100011100010110101001000101110011001111;
#1 $display("%b", po);
# 1  pi=207'b101001000111000001011011100101010010110001001000101110010100111001010100110111010111001000000111010000110000100110011100101111000000001100101100101111111010011001001111101010010010111010000000101000000000100;
#1 $display("%b", po);
# 1  pi=207'b000110111110100111001101011101010001110001111101011101101110111010011100100101111001111001000110000011011001000110100010001011100110111110010110010001111011110101111110101110000000010010100010100010101001011;
#1 $display("%b", po);
# 1  pi=207'b000001111111000011011000100110000011001001101000100010010100100010100011000110000101011000000001101100101010101111101110100000101100010110010101000110011001100101001010010010001000111011111110011011110100010;
#1 $display("%b", po);
# 1  pi=207'b010101011010001111010101101011101101001000111001010010100111000010100111110111001000010000000111101000100100000100110011011100101110101111000011111110101110111010000010101001110011110111000111111100010010011;
#1 $display("%b", po);
# 1  pi=207'b001100100000101001010010000100001001111101011101101110110000111100011011010110110101001010100011111100000010000110101001111101000001011101010110100110000010110110001110010101000100111001110111000001111101100;
#1 $display("%b", po);
# 1  pi=207'b010010010000011111111101101000101010100110011110111011001000100011101101010011000111100000000111110100100110011011000101110110100100001111011111100100110000000101011111001100101100001110010111110011000111000;
#1 $display("%b", po);
# 1  pi=207'b001010100011110000111110000110010101010000010001011001001000001111010010000001011110000011001001001111110010010100001111011100000000110010101010011101101001011110011100101100110100110110011101110110001010011;
#1 $display("%b", po);
# 1  pi=207'b111000001010001000011000101011111100111111011001110111000100000110001111101000111000111110100111111100111100100101011010101001001100010110000101110010100000110100111010000011010011011000100001010001101111011;
#1 $display("%b", po);
# 1  pi=207'b100011100111101001001110000100000100000100101100001000001110010111011010100010010101111000000010110110100001001000010001000101110011010101110000010000110101110011010010100111111010101110001011101110010010011;
#1 $display("%b", po);
# 1  pi=207'b011000001100000101100111000100110110001011110010101111000001111011010011110000101000010100100000111111001100111101100101110011010011101011111011111110000001111101000000100010011100110111001011000101111110010;
#1 $display("%b", po);
# 1  pi=207'b100101010001110001101011001111110001110100100101101100001100011110000111111101000011111101100100000101111100010000111100111101010110100100011110010111010101001000001000100001010101110001100011110000010011101;
#1 $display("%b", po);
# 1  pi=207'b110100001100101100011101111100111000101001101001010101001111111101111001010011110001101010100101111010111101101010100101101001001100110011000111101110101010101001111001110110100000000110110110111110101010100;
#1 $display("%b", po);
# 1  pi=207'b111010010110001000111100110101101010100111110001011011101101100111101101011011010110111110101010100011111101111000110011101111011000100011110011001101110011110111111011110010101100011000010010010100000111101;
#1 $display("%b", po);
# 1  pi=207'b010100111100111001000010110110000000001001111011111100110101100110000100111000110011001101011000101000000111000001101101010001100111111000101101101001111111110011100101111100011110111110000011100000110001011;
#1 $display("%b", po);
# 1  pi=207'b001011001000101100010011101100110111011101100010011001100100010011001100101000100101001111101000011101110100110010111001110010000101110000100000000010100111100100101000000100110001101101100101010101001111011;
#1 $display("%b", po);
# 1  pi=207'b110000001101110011010111110000000010100000100101111010001011101001111111110000110101001101100010101011001110010010110101010110101011001010110001100011001011001100110001101010011101011011100110101100110000110;
#1 $display("%b", po);
# 1  pi=207'b011000100001101011101110011111110110000100010011111111101101111000010011011111101010010010101010110111100011111101000111110001111001100111100110111011011011100111010101010111100001011100110110010001010100101;
#1 $display("%b", po);
# 1  pi=207'b111101001000100110000010100101011001000110011010111010100100101111101111110111100001111000100111110010111110111001011010110010010100011000001101001100111010111011100110001011000000100110111101101101101100110;
#1 $display("%b", po);
# 1  pi=207'b001110001101111100111011000111010101110011011111111011001100010111000110100011011101010001011000100110001100110100101000110011111011010011011001011010011000010110110110111010110000101011001001010110001111010;
#1 $display("%b", po);
# 1  pi=207'b101011000000011001010111000101101001110110010011101110010011100010010101010110110111010011001111010101101010001100000111110111000010001111000000010001001001011001000100000000000001011010101001101100000100111;
#1 $display("%b", po);
# 1  pi=207'b101110111110010101110101100100011001011001000010100011010000011111011000100010001110011000110000111100001011001100001100010110010110101101110001011111010011111100101010101111101100010100011111111100011000001;
#1 $display("%b", po);
# 1  pi=207'b100010001100001100101001100100011011111001011110101011001111101100011001000001100100001111101110000000100101101010101011010010011101111001110101110001100000110110100001111001100000110101101101100111110110111;
#1 $display("%b", po);
# 1  pi=207'b011010001111100000100100100001110011001100001111111111001010010110000010011110000001010101001010011101010001000110110100011011000100000000111000101110000000110010110110001110000100111001011100101001110111011;
#1 $display("%b", po);
# 1  pi=207'b000011110111011100111110101000011101110101011010111010001011001011110110001110100110110100110101101101010100101000010000000001101000010111001001011000001011001101010010110011000001000110000110110111100100111;
#1 $display("%b", po);
# 1  pi=207'b110010111111100000011010101001110111101100110100101111110011010000101110101001001000111000101011001110010101000100010100000110010101000001000011011000110110011111101101100110011110101010000101111111111011110;
#1 $display("%b", po);
# 1  pi=207'b001000011011110010111100111000100011100010101010000100000010110010010000100100001100000001000111000111100110010001111110101111000110100001111000001011101011100011110101100111000010101110100100010011101000000;
#1 $display("%b", po);
# 1  pi=207'b001100011011100100011101010101000100101101011010110011101010110111010101000111101001000001111100110101110000111101000010001100001100010100100101100010010000110101101011010101101110100000010010010010011011100;
#1 $display("%b", po);
# 1  pi=207'b110000101000100100011111100000011000011001001101011000011011000110101101100000001000001110100010111111011100010011111111011110111011101001010110101100000001101101100100000011011011111011011001000100110000011;
#1 $display("%b", po);
# 1  pi=207'b110110111110010001011010011000100100100111001011000010101001110010001100001001000010011110111011100110101110100100010000000010000110110001110010110101011010000100000011101101001011001101101110001110100001000;
#1 $display("%b", po);
# 1  pi=207'b101010000100101111100011110111000000100011010100110001001111111011011011100010100010000100000011101001111111101000010101000100100101111011110100010111101101011110101011011110111111001111000111000001101101000;
#1 $display("%b", po);
# 1  pi=207'b010101011101010001001111100101001110010010110101010000010001101011001010010011000001110110100010100101010001001110001001001011000010011001011010110101110000010100101011111101010001001101011111000100010000100;
#1 $display("%b", po);
# 1  pi=207'b000101100110010001000100001111011010101100111110000000101100111100000011000111100100101010001100101010110011001110101011100111101111100100100011111100101110100110110001101011100111001001011100111100111011010;
#1 $display("%b", po);
# 1  pi=207'b110111101001010111001001111010100010110000001011001010010010000111000000100110000001110000100101011100101101100101011000101010001111101111101001001100010100001101011010110001000011011010011110101000100011001;
#1 $display("%b", po);
# 1  pi=207'b101010101000111011001111111111100001111111010101011101100000000000101000001001011000100111100110010110010101001000011111000010100111100001011111100010011001101111001011110001000011011100011110011101100000111;
#1 $display("%b", po);
# 1  pi=207'b100110110110111101011101011101110001011100000110001000011010010100110010000000111010110001011010110000010100001100001000011110101011111100110110100110000001001101111010010100001101001011111101000101100010000;
#1 $display("%b", po);
# 1  pi=207'b101001011111011110100001001110010000110000110011110000110011001110011010011101100111111011000010111100010010000100101010110110000111100111010010111010110000001111101000111100100110101011000011001000011011100;
#1 $display("%b", po);
# 1  pi=207'b110011010100001101110011111111101110110101000111101111100110111111000100100010100010011110101111001010010111110111010110010101010101011011111001110111010010111111001101000001010010100111011000101011000110101;
#1 $display("%b", po);
# 1  pi=207'b100011101010110000001111001011010111000001010001110101100101110110111011100011110000000010111110000110111111010011001011100010010111010011011100010100010011010010001111101111011101101011011111000110110000001;
#1 $display("%b", po);
# 1  pi=207'b111100011010111101100100110110110010001000011110100000000011110110000000111101000111000010000101100101101010001100110101101011111001000011000100110000000100101010100111010001100001001101101111001011011010110;
#1 $display("%b", po);
# 1  pi=207'b101001101100011000100000000000001001011001010100110010010010001111001011111001101001001010000101100111111101110100111011101011100011111111011100110110000010100110000110111000001100101011110010011100010111011;
#1 $display("%b", po);
# 1  pi=207'b100111000001001001001001111000110000100111001000010011101001010100011111101110100000110000111000011000001100111011010110001111011011101010100111111000110110001010110000100010101001001110111011011011111001111;
#1 $display("%b", po);
# 1  pi=207'b110011011010010011000001001011000100101110110000001110100110001000010101111111001001011010011001011001001100111000110001000010011110001100101111001010000111100111100111011000000010000001000010011010000110111;
#1 $display("%b", po);
# 1  pi=207'b100100110111010100000010001001111001100110110010101010001110000111001010001001101010000101100100110100000111010010000111100000101100000000110010000001010001110101001001100100001001001010011100000001000101010;
#1 $display("%b", po);
# 1  pi=207'b110100011011101101011010011100111100110110110100011011000110000001111101111100001010000000000101010111100101101001100011011101110110101000001011001001000010010111100110000101011001010110011011000110001010111;
#1 $display("%b", po);
# 1  pi=207'b001001111011110111100101001111111110110001000001111010000100001101101111001110110100110001010011110111110100101110101000010101100000100000011101010010000111011101000100010110100110001100110010010000110100110;
#1 $display("%b", po);
# 1  pi=207'b011000011111011000101000010100001111001010000110010101000010100111000000010110000001101110110000001010011110110001100110101001001101011011001101001110111010111011011000010001100000111010100110110010101001001;
#1 $display("%b", po);
# 1  pi=207'b011010110100010101101100001100011111111110111111100011111110110001100110001100111101001111000101110110011101011111110011100100011010010011100000101100111101011000110111000010111011100111000110110111000100111;
#1 $display("%b", po);
# 1  pi=207'b001110101010110101100100100110111010110011010111011011110111000111010111111000101000011101101101101110000001000000111100111110100101011001011001000010011011111000110001100001010011001000111000100111101101110;
#1 $display("%b", po);
# 1  pi=207'b010110010110001100100001111010011100010101011001100000111000001011011001100101001011000101101100010101100010000011100010101000110111011011101000100111000011110111010000000111011110100011010100001101100010110;
#1 $display("%b", po);
# 1  pi=207'b001101101011010101010000100100101010100111110011110000111010110001111111101000100011001101010000110000110110110010010001110111000111011001110000110010110110010001101101010001110111011001111011110110110000010;
#1 $display("%b", po);
# 1  pi=207'b100010010100000001001110110011000101011011010100100110110111000110101000011011011010100100100110001100000011111110100011011010010100101101000010110000011110100100011010000101010110100111011111011111111111001;
#1 $display("%b", po);
# 1  pi=207'b000011100110100001010011000001110110000101111010111011001000110111010000011101010101100010001000100100010010001001011010001111011001100101100110011111100100111000010000111110000111000011110111100110011001111;
#1 $display("%b", po);
# 1  pi=207'b111010011101101000101010000101001010110010011110111100011110000110011101000011001101010000100111111111011000111100100110101101110000000100000001110110010011101100010111110110101100110001001110111100010101010;
#1 $display("%b", po);
# 1  pi=207'b100101011110011001000110010001011110010100101001011001010100000011000010010111111011110010000001110001011101100101001011011001101000101110100101010111001010010011000000100001010110110011011111110101001111100;
#1 $display("%b", po);
# 1  pi=207'b101110000100100010000011000101111011000011001100111111001110000000001111000100101100000100111010010011011001111101000111001111111100100001010110011010110110010100100000110110001010100100010001001110110100100;
#1 $display("%b", po);
# 1  pi=207'b011000101011111111001011101101001011000010101101110010000000010101100001110010110101111100011010000111010011100001100100110011111101111000000010010000111111010111111011011101101100011010100100010001010111001;
#1 $display("%b", po);
# 1  pi=207'b011001000000010010010000010010000001011000110011001000111000011000000000010111010101100101101101101110100100000101101100101000101010110101000101001100111011101100000001000100010100000101111001010010110101101;
#1 $display("%b", po);
# 1  pi=207'b000111000010110000100100110101010100010001110011110000110011011110101011100000011001111100000000000111110010000000010000000000000001001111010101011001001010100010001011111010101010010110000111011001101000001;
#1 $display("%b", po);
# 1  pi=207'b100110001100001101101111001110101111011110110001001001111101101101011111000111100110101001000111000111111000000010110000110011101000110110110110110100001000111011111100111110100111001111101010101111010001010;
#1 $display("%b", po);
# 1  pi=207'b111110100001001100100000011111100011001110000000101101010110010110101010011000111000001111001100101111101001111101101111011101000100001100000001111000000110011010001101110000100011110100001100111111000011100;
#1 $display("%b", po);
# 1  pi=207'b001110110011001010110101110001110101000010001110011001101111001001000000000000000001101011001111011001101101110111110101001100100110100011001101111110011101000111100111011100011010011101110110100110001110100;
#1 $display("%b", po);
# 1  pi=207'b010101111010001000100100000101001111000010010010110110101011110011110011101011000100010101110011101010000001010000110011010011100000011001011111110111001110101100100011000100100010010100011010101010100100011;
#1 $display("%b", po);
# 1  pi=207'b010110110100100100001111001100010010011101100100000110001111110011001101011001101100110000111111000111000011110100001110100000000011111000100010011110011011001010111100101001001000010000111110011101001101100;
#1 $display("%b", po);
# 1  pi=207'b001000110010000101110111011111101011101110101010001001101000100011000110110010001100000010001111011111001001100101111111001110110100100000001101001000010000111001011101010000011101010101110010101100011000010;
#1 $display("%b", po);
# 1  pi=207'b000011000011111101011011010101001110001111100001000101000100000000101100011001000101000100011000101110000100001011100001011001101110101011011010101011001110111001010111100111010011111110110100001011110001101;
#1 $display("%b", po);
# 1  pi=207'b001000110000000000111010111001110101011001111110111110011101011100010011011011101110000001000000111010110011001011100000111000010111001011011111101110011000000100001100011010000001010000010010000100001101100;
#1 $display("%b", po);
# 1  pi=207'b010110100001111101111001010100100001010001111110000001000001100000000101111111010101100001100001001110100010010100011001111101110010001001010101100000011001101100100110100111101000101110000101110001100010010;
#1 $display("%b", po);
# 1  pi=207'b111011111011000010101100101010000110011011101111010000011110001000100101101110011010011000001100001010010100110011100000100100111110100100010011110000101110001100000011001010011011000101111010011001111010011;
#1 $display("%b", po);
# 1  pi=207'b001000011100000011110111000010011110101111100101100011010001001110000101011111111010101010110100011001001100101011110100000010000011111011011110100001110101101110100111010100101100001111010111110110010101111;
#1 $display("%b", po);
# 1  pi=207'b100011000001110100110001001101100000111000101111001111001110100001000001101101010100111101010010011001100110001011111000001010101000101010111100000000111100100001000111110000001100001111010001000111010100001;
#1 $display("%b", po);
# 1  pi=207'b111100110100000011100101001011010110001010110101010111010110111111101101011011001101011110110010010100101110011101000011111000110101010110001100001001110100100010011001100111100010000001110110101010101111010;
#1 $display("%b", po);
# 1  pi=207'b101010111000111011111111101010010100101100100010000111100010101111000010100010011001000000011011010010110101111110010101000100110111001110111010110111101101001111110111101101011001100001111011110011100000000;
#1 $display("%b", po);
# 1  pi=207'b100100010011110111000110101100000101011011101011010110100001110011001010011100100100100001001100110011111110111001010111111000101111100110111101110111111011000011011000000001010001001010110111011101000010011;
#1 $display("%b", po);
# 1  pi=207'b100000101010011001111100110101100011110011000000001111010100110110001010010101001110110101001100010110110111101110111111011100100001010000000010001000101101010111001101010111111111010110101111011111010010101;
#1 $display("%b", po);
# 1  pi=207'b011010001011110000011001000110000100101101101000111010000100000001010010111010010100111111111111010100100100111001100001001111111101101011010100111001101110010111110101111010100111100101110001100001100110110;
#1 $display("%b", po);
# 1  pi=207'b011011110111101101000001001100011111100110111001101100000111000000110001000101011110110011011001100100101001100100101110101100101010001000000110000110100100101010100011001101001100110011111001011100110110000;
#1 $display("%b", po);
# 1  pi=207'b000011000101011011011111011001100000000111010001011100000010111001011110000000101001010101000010100001001111111100100001111101000000000000110010110110011110101001001111110000100010100110110001100001110111110;
#1 $display("%b", po);
# 1  pi=207'b110000010011110001111010110100111000101000001001101011010101110000011010000100001000111111111100110010110101001001011100001110011110110110110010000001100000000000100110110110011100100000111110000100101011110;
#1 $display("%b", po);
# 1  pi=207'b100110001111111100110110110110111101111110011000111001001110110000011001011110111111011000010110010101000011011100100101010010001011100101100001110011011111110110011111100110111100110100011011110101011010000;
#1 $display("%b", po);
# 1  pi=207'b000100101101111110011010110101111000000001000100001010110000000010111110011010011101100101110101000001111100001000100010111101011000011101111100101011010001100101110001111001110000101101010001110101000110001;
#1 $display("%b", po);
# 1  pi=207'b010010110010101111101000100001010000001000010101011010001001111100111110000001001010101100111111010010101101101110100111111111000100011100011100111001011111010001100001111111110000011110011010001001100010110;
#1 $display("%b", po);
# 1  pi=207'b000001111100001111000001101000100000101011011100011110000101010001111100001111100011110001010101110011111100111010011011110111010110110011000000001111110110100100000100111000011010100110100100110101000101011;
#1 $display("%b", po);
# 1  pi=207'b000100111110001111000001101110011111010000111101011101100011011110110111110000001011010010101100101001101000011111010010110100010111000110101100110010000101001010110001011100100001110101110110111110001001001;
#1 $display("%b", po);
# 1  pi=207'b111100000100101111001101011001111001010100001101110101000011001010100110101110011111000100101011001001001010010111100010101011011001010010110000111110101101111000110100110000001001011000010111011000010010011;
#1 $display("%b", po);
# 1  pi=207'b001100110110100011100100111010101111000001110111101100111010010011000010001011111000110111110110111001110001110110100100001111100110011000001000101111110001000101011101010000010011010001101001010010111111011;
#1 $display("%b", po);
# 1  pi=207'b000010111000010111110101010000101010000001010001011111000011111100001100110000001001001011100010001001110011010010010111010110000110001101010011100000000010010111000100010100010101010101011000010111111010101;
#1 $display("%b", po);
# 1  pi=207'b101100010100000000011000111110101101101111010111100111001000010011101100100100100100001001010101000011010000001101010100011100010001110111110100011110111011011100101101110100100010101001101101001101101011100;
#1 $display("%b", po);
# 1  pi=207'b101101011111111101100001011110111000011010101100110100101000100011110110010100001110100001001010000001100101011111010011011101100100001110101100101100011010101111000101000001100101010001101000110110011001000;
#1 $display("%b", po);
# 1  pi=207'b010100110011011010001111000000111010010100001011001110011001011110000100011011100011010010111010111101011001000000001010111001000101110101000110000101011111110110101000111100011111011111011000001111101001011;
#1 $display("%b", po);
# 1  pi=207'b100011111001010000111001010110110111111010100001110000100111100000110000100000000011100001000100111101101101000011101101111111010000001111010100000001000111001111011011111110110110000110110110000001011111110;
#1 $display("%b", po);
# 1  pi=207'b001101110110111010001000011010111100100011001110110011010100011011110101001010110000100100001111001010101110101011011100000000110100011000001001111110100111010001110111001100000000000000100011010111100001111;
#1 $display("%b", po);
# 1  pi=207'b110010001011111000000110010001111011110101100101110010001111111111010111111101100000001100111101010010011010100100101010000011100011000110110010001001100011100000000110111110110110011110101001001110111001100;
#1 $display("%b", po);
# 1  pi=207'b000011000101110101010011111001100110100000111101001011000101110000100001011001101101010100101100111001110111010111111100110001100100101011110011000100110001110000100000110110110101100011111111111110111100001;
#1 $display("%b", po);
# 1  pi=207'b010111000010100011001011110111010010110100010101000010111111101101110010100110110110111001101000000001001100000110010101001000000001010110001010011110111000111010011100001100101011100001001101010010001011010;
#1 $display("%b", po);
# 1  pi=207'b101001011110101001010100010100101110001111000000111001001011111101111011100111010100001011010001101101100000110010001010101001111001001010001010000100101011000001010110011011100110110111101011000110000100010;
#1 $display("%b", po);
# 1  pi=207'b011110100011101101010001110101011100001110000110001010001101011101000001011010110100111100001110110001010011000000010001000100010111100000011100111110101000001110011110000001110010101100101101111111001010001;
#1 $display("%b", po);
# 1  pi=207'b110110001011110001000000010110001011111110101111100011110101001110101001110010110001111000000101100000101010110111110111110100111101100001001011011010010000011100010111110101111000111100100010010101001001011;
#1 $display("%b", po);
# 1  pi=207'b010111001111011011111101011010110101100010100001000000000001001101000001111000111011101111011111001010110010100101011000011111111110001011001001011100111000011011010111000001001001011011000100000110011110001;
#1 $display("%b", po);
# 1  pi=207'b011001010001011010001000010110110111101001011111001111101110100000101011011110110010001110101001111000100100011101111111000011000001111010101101001101111011000010011000011101000111110000001100001100110000001;
#1 $display("%b", po);
# 1  pi=207'b110100111001000111110010001100001000011101011001000011011101010011111011010001100110000011000110100000111101010000010001011101101011001011010100100011101011011111101100110101010100110010001110110000110110111;
#1 $display("%b", po);
# 1  pi=207'b110010101110101101101010100011111010001110000001000000111100111001010100101100111011101100010001100011001011001001110100010010010111001000100000110010001110101110000101010100011011110011110110100100111101101;
#1 $display("%b", po);
# 1  pi=207'b001110100010011011100010111110110110101100010001011010000011101000101100110101100001010111011110110100010111110110111110111100101001001011110111000110011010010001001111101111100110110001001000110010010110011;
#1 $display("%b", po);
# 1  pi=207'b001111110000001000010110100010010110000000000001000001000100100010001100001111100110101100011010111010101010101111100100110101111110001010111111100011011001111111111110111011101110101001001110000110100101010;
#1 $display("%b", po);
# 1  pi=207'b001111101111101001100001010001101010100100010110111111100010000010100011011110001111101110100111110101101001000100001011101100010111011001101010011100110111110000000101100101001001110011011111000110001110011;
#1 $display("%b", po);
# 1  pi=207'b001110111011101111011011010111111100010000010010100101000111110101010110001100001010001101011000010001110111100100011011110001101010101011111111000111100101100001100100101100100101011100110111110000111001001;
#1 $display("%b", po);
# 1  pi=207'b100000001000000010100010011010011100101001100110111111100010111101111001101011001100101101010001010011101111011001100001011110000001000101000011000000110011100001011000010001010101011101101100011000010111101;
#1 $display("%b", po);
# 1  pi=207'b001001111100100011110111101011001011101110111000111100010110110110100100111010011000101011011101110111011001010011010001101001111110101001010100011101010110000000111001110110100001000110011010011110101100111;
#1 $display("%b", po);
# 1  pi=207'b001101100111111101101101100110111100111010011100111101010011110100011101010011010101110100110101110111010010001001101011000010001100010000001100101110000100100000111000010001000110111111010010111010001100111;
#1 $display("%b", po);
# 1  pi=207'b100100000100011000000111011111010011110110110100010000111010011011001101110101110101110101101100101001010111001110111011010001111011001010011000111011010011011000011000000101011000001101111011001010111001001;
#1 $display("%b", po);
# 1  pi=207'b110101101000001001011011010011011010011101101010000011111100101011100010100001101011110101111100011010101110111111011010011111000111101101101110100000001101111010011010101111101111111011001001001101000110001;
#1 $display("%b", po);
# 1  pi=207'b100000011111101000101010001110101111111010111000110010100001000101111110001100101011000010111000101000011000101100110101111011000010011100101101001001000001000110010010000100000110100010011010110110111000110;
#1 $display("%b", po);
# 1  pi=207'b001001110000110110011011101001101011100111001111110111011011001110110010001101001011111010001101111100010010101110011011011010100011001010001101101100111100011111111001101000110001001000100000111010101011000;
#1 $display("%b", po);
# 1  pi=207'b001001110011010110011100011111100011110111111000110011000110000110100000111111010000100010000010100101001000010011000110000110111011001001111111101001111111011100100011110100101101011111111000110000101100011;
#1 $display("%b", po);
# 1  pi=207'b101110000110001011111110011000000111101000100100011000110110000110110110010110110101101000101100001000110001110100110001001000000101110011000110101111011000011001110101011001111110111000011100001010110111111;
#1 $display("%b", po);
# 1  pi=207'b100010011101100001011011011001101110001001101011100101100011001010110111011100100011100111001100101011010011100001000010011111011111010010000001110110000000010100011110101111001000111101111110110010110101001;
#1 $display("%b", po);
# 1  pi=207'b010100000101100100001000001100100000101111010011111010011000101000001101011111000000001010110100110011000110111100011100101011100100110111100111010101011000100010110010001011101001010101100011001010011001011;
#1 $display("%b", po);
# 1  pi=207'b010000000000110010101000101010000001000110110001001101011011100011111110111001010101100100111110101001101111110001101100100100011011000100001011000000001001111111111011000101000110000011101100111111001010010;
#1 $display("%b", po);
# 1  pi=207'b100100110101100111010100000001100011100111001101101111001000011111111110100111101010011110000111110010001111100011110101111101101011001101101000011011001000010101011011110111001100011101010000111101111011011;
#1 $display("%b", po);
# 1  pi=207'b000001101001000000100111100001110111111001001000100101000000011011010010111010000111011111111100111100101100111101100111111000010001011101110001000001101101111110111100000001100001110011011001111110101100011;
#1 $display("%b", po);
# 1  pi=207'b111100000000100000110011101000100000000001100110110010100011011111100110001000011010110011010110100100110101010010001010000010000001100101001101011100111100010101101001001111111111110110001001001010111011000;
#1 $display("%b", po);
# 1  pi=207'b010001100010110010010000001001011100001000010000110111011111100001001001011101101001001100111111101111110010100110001111000001011001000010011100000010011111000100101000011011010011110101101000011101110101001;
#1 $display("%b", po);
# 1  pi=207'b000111100000011010010100001001010001100010011011110110110000101110110001000011000100100001011011000010100001100011001011000000011110101001011110101100000100100110110101011101101010000000100101100000000010111;
#1 $display("%b", po);
# 1  pi=207'b010100010001001100011110011101111100011011110101100100100110001101000100111110010001110111111000011101010110110110111001011010101110110111111111111111101010101000100011101110101111101010001111111101110100011;
#1 $display("%b", po);
# 1  pi=207'b011100010000101010000001010110000011100000101010000111100010110010101111110101100000011001010011000000100100111001101100000100110110010111001011011011111000101001101011111011100101011111010111001111110010011;
#1 $display("%b", po);
# 1  pi=207'b011011110110011100110110010011111101001100101100101100101010010111001100001111001110001010100100110101110011001010100110000000100001011101111100010111111011011110011011101001010010110010111010100000111101001;
#1 $display("%b", po);
# 1  pi=207'b101101100001100101010001011101100011111010101000101110001000110100100100110001101110110011101110100101010010110001001110010100111011000100101000000010001101010101111101100010111111101110111100001000101110110;
#1 $display("%b", po);
# 1  pi=207'b100101001001101001010101110011000011111111101010010111111000101101000000111011010001110000101111110000101000100111000110111000010101101001011110110110110101011100101000110010010101100001100000101010101100010;
#1 $display("%b", po);
# 1  pi=207'b001001010011000111001110001111000100000000001111100101100111110110101111110110100000000010010100101010111011111010100110010001101001011111001100111111000111011011100001010101110111101010001001111110100100111;
#1 $display("%b", po);
# 1  pi=207'b100010111110011100011000001000010110110110110001110000001110110100100100001010000011100111101111101101111010000001011100000101110000011001001110101010001010111011111011100111110111111101100101100010010010011;
#1 $display("%b", po);
# 1  pi=207'b011001011011100100000000110000110110011101011101001011000000110101111010110101111111111100010111001001101100110110010001011010100101001010011000010101011010111000001001001101110100110111001000011010110100101;
#1 $display("%b", po);
# 1  pi=207'b001111010011001010011100011111110101101101110001001011100110101010110001100010100110010000110010110010010101101001111011000011101000001000110110100011000011011010010010101000110000101110000100101110110100000;
#1 $display("%b", po);
# 1  pi=207'b101011100010111111011000101110111000011100011110001100100011101010011110101011111100000111010100001001001100100001100100111011110111001000000010000101100010001001100011011101111001100100001001110101001110110;
#1 $display("%b", po);
# 1  pi=207'b100110011110010100101101001101110010101110001011110011001101000001011111000110001000110010100111000111000110001101111101100100000111001110000110011100011000010110000110001100100101110000001110110010011011010;
#1 $display("%b", po);
# 1  pi=207'b110100001110111100001101001001000001100101010101100011100000001111111010011110010111000100100001101010100011001111101000100100111000001111110100101110010001111000110101100101110011001100111011001001000011001;
#1 $display("%b", po);
# 1  pi=207'b000110011111111000111111110101101110000101001010101110100010110111000000011001010010110010111010010000000110000110000111011010111010100011110101011110011101100000001110110100010110111111000110010110010010100;
#1 $display("%b", po);
# 1  pi=207'b110011101011100011111111001010101000100001111100001100101001100010001000111100111001011011110000111111111110001100010000110011110111011001001001010011000101100111101100011110100001110000010100001100011110000;
#1 $display("%b", po);
# 1  pi=207'b001010100010101011011110100001001100111110101110011000001011011011101100111101101111100001100111101100001011011010010111110100011001101010110000100111111000111010101100110011111101101111101100000100101001111;
#1 $display("%b", po);
# 1  pi=207'b000110000110101100101111011000110000010111111100011010111010011111110101001001010101011001110100111001010101111101101000101001000000001100011100000001111110000010111010110010101010000011101000010100010110111;
#1 $display("%b", po);
# 1  pi=207'b000101100000001110111000110001100101100000010010001001100101111011011100101110111110110001001011100111000101110100001010010101110000101101111111000100011101010100010010000010001101010001100111110101101111001;
#1 $display("%b", po);
# 1  pi=207'b111001111100101001111101000010011010001100100101100110111100100100011000001000101101011101010000110110010100101111010111111110001000110000000000100001011011111100010110111011100010001110101011011101001010110;
#1 $display("%b", po);
# 1  pi=207'b110000011000011101100100100110100101001110110110101001110001001010010000001100110011011011101111010001110001101100000111001111010100011011000111110011000111100000000100100100110111010000001000010111111111100;
#1 $display("%b", po);
# 1  pi=207'b100001001010110010111110100010101010100011100100100111111000100100011001100011000010010101110001110010000100010111111101100110001001100010101101110010001100010100111110111001011101111010100011000010101111011;
#1 $display("%b", po);
# 1  pi=207'b010100011100110110100011111101010001100010111100110110100001111010110011100110001101011000000111110011000100010100001111000000001000111011110101110111000100011001000011101101100101101111100110110001011111100;
#1 $display("%b", po);
# 1  pi=207'b100001110011001010011110011001010101011101111111101100110000101001111111011110011111000000111000100101111101111101111110010100011101100000101010011001000100101110100101101011000111011000011110001100000010110;
#1 $display("%b", po);
# 1  pi=207'b011101011000001110010011111000111110100110110010011011001110100000111001011100111000111001001010001000111011011110100110101100000011000111111000010011100100110000100011111101111101101110111111111000000111110;
#1 $display("%b", po);
# 1  pi=207'b100101110110001011000011110010011110010101010001010011000100100000111101101000111011011010111110011010101010110110110011101101001110110111101010101101010001010001000111000101000111010110110000010010100001101;
#1 $display("%b", po);
# 1  pi=207'b101001110100101010111100110111011000111011101000010100101101111101001010001110011100111001111010110000010101100110000111101000100111000100001110111110100010110001101011001010100001000111100000100111011011010;
#1 $display("%b", po);
# 1  pi=207'b100010110010010101000110010110101101101111111101001101000101100011110101110010011010100001001011010110111111100010000111101011100110011000011111001000000101101101000111100101000000100100000101010111100000101;
#1 $display("%b", po);
# 1  pi=207'b011001010010001111100011110010000110010010000101001100000111100011110011111010011101010101001101000001010001111011011111100010100110100000011001110101001001100110100011001000000001111001010111011111010101110;
#1 $display("%b", po);
# 1  pi=207'b000001101100100011011001101100000000001100010100101111000000011000110111101011111010110010011000110001101111001101010100111101001001100100001011100011111101110000000010110010101011111010001011011111000001111;
#1 $display("%b", po);
# 1  pi=207'b100111101100011111110110111001001010111010000100011010011111111101111110111000100101001100101100000110001000111001111101011000100010010101010000010010001000110010010101110000110111000101011111111011001001110;
#1 $display("%b", po);
# 1  pi=207'b110111000001000011110010101011001101001111001010000101010001101010010001001110011010101100111000000000110111111010000010010010100101110111101100000010101010010100100101011101001111111001011110100001011011001;
#1 $display("%b", po);
# 1  pi=207'b111110101011001010110100010101000000101100010000100111000010011110011111001010011101001010010010100110110111101001010000100001011100101000100110011010010011100110111110110100011100101100011111111011100111110;
#1 $display("%b", po);
# 1  pi=207'b110000001101110011011111100000011000110110110000010000111110111000100100001110110111110110010000001101000100111000111000111111101111010000100101101001101001100110010000100000101011000011011000001111000101010;
#1 $display("%b", po);
# 1  pi=207'b110101000101001110001011010100100010001101100101100111100100001010011010010101001110100001000011001001100010011010101000101110110110111010111100011000010010001111111110001010011101110010111111101101101111001;
#1 $display("%b", po);
# 1  pi=207'b010110000111000111100111101010001100101110001010101001000010101111001110001110100010000110010000010111001000001011101001010011010111110100001111000111101111000110100001000001110000100110001111011000011100111;
#1 $display("%b", po);
# 1  pi=207'b111011011100001100111011110100110001100011000110011000010001001010001100011001111111100100101101110101110010010010010000001001001010110000110100001000011010101110101011011010110101111010010100010010011101110;
#1 $display("%b", po);
# 1  pi=207'b001001000000001011100101011110111100100001110001101100100001000101111110110111101000010110100011010010011010010110010011101110011110010000111110110100110001010010011100111111010111000110000000100110101100111;
#1 $display("%b", po);
# 1  pi=207'b101010111100000001001010001000101011100001101111000001010001100101010111000011011001000100110011000111110101101110110110100110001111001110001111011101101011001000001110000110101110100111000110001001101110101;
#1 $display("%b", po);
# 1  pi=207'b110111110010001000110100100111010101001110100111101100010101101111010110110000011111110101100001011100011001011101010101111010100010111000101010101000000111110001110100101101001001000110111110110101001000011;
#1 $display("%b", po);
# 1  pi=207'b011100001101111010010110101111100011010110110010010111001101010000001100110011101100000101110110000101000110101111110001000111101100100100110010101111001101010100011011001010111100110001111000001001001001110;
#1 $display("%b", po);
# 1  pi=207'b100111111101110111110101001101100100110111110110010101011000100101010010001010110101001111101001100011001111011001010100011100100010110100110010101010011111011010110010101000011100001110101110001000000110101;
#1 $display("%b", po);
# 1  pi=207'b001001010011000001010011110001000000100111001010101111111011100000100110111101101111010010011111011000100000011000001110011111001011101110001001111011101110110001110100100000101111111110010101000110011111110;
#1 $display("%b", po);
# 1  pi=207'b110010001111011111110010101110100000011100100100111110001001010011100001111000110101111011110110111100110001000001110011110111010010010000101100010001110111011000101110000111100010101000100010101101001011001;
#1 $display("%b", po);
# 1  pi=207'b001010111101111011000110001101011101100100011001000010101010100000001100010011100101011101110011100101101011100100111111000000000000100101111011110110010111000000011101101001110000110100111000100111011000000;
#1 $display("%b", po);
# 1  pi=207'b000111110110100111111101010001001101100100001001100011110011010110111000010010010110111001111011010000100011010110101110100101010010011101111001110011001110001100110101110001101010011001010011101000011111110;
#1 $display("%b", po);
# 1  pi=207'b000100001010110101100010110011001001110011010101110101111000000101010100001101100010101111000111110100111111110101110011000011010110000101001101110011100100110111101100111110110010111000010001111101101010001;
#1 $display("%b", po);
# 1  pi=207'b110011110000101010111111101001111101101000000110111010100111011100000010011011110010111011101011001011001000100111000101111111000111110011110001110100101111001001100111001011000100101010010010010010111011010;
#1 $display("%b", po);
# 1  pi=207'b011100110000001110101010011110010101001110110010101001001111000001001011011000101100001000010100001101101100001000111101110001111101001101101110101100101100000000101111001010101101101111101101010111001011100;
#1 $display("%b", po);
# 1  pi=207'b000101001111111001100101001011000001000100010111110010101011101000010101000010001000011001000011111100011010111111011001000010010011000011001011110001001111100110000111010100010001000000001010001010101101101;
#1 $display("%b", po);
# 1  pi=207'b001111101001001101110110111000110010101110111011101101101011111100101001000111101110011110110110001010000110111100100001010110001101011110110000111101001100100001001101101001101101000111111011101101001100101;
#1 $display("%b", po);
# 1  pi=207'b111100000011111011101111010111110101111011000101101111001010111000111101111000000111100111001111101011110001000010011101111111111010000100100010001100011011100010000110111011101010001111010010111100001110011;
#1 $display("%b", po);
# 1  pi=207'b011010010010100101001000101001100110110101011101110100110010011100101100011111101001011110111011001100010011010111010100100100101111101000000111000101011111110110000101111000001011111111110110000100110000101;
#1 $display("%b", po);
# 1  pi=207'b110100011100000010110111100010010110011100101111110101111110000010101010100101011111111000011000010110101111000011111001111100101110000001000101101010101110000000111010110110111010111001101100010001101110100;
#1 $display("%b", po);
# 1  pi=207'b110110011110001000010101010001010110111000110001011101010001111101010100100010100110010101011000010101010000000100011110111110000101100011000000100111111101111001000110110000010000100011100001010111111111110;
#1 $display("%b", po);
# 1  pi=207'b001100110010110000001001001101000011000001001001111110111010110001001101000000100110001001000000110001100101011011010101010010101101110100001000000011101000100011001000111010111110110101111100001100111110001;
#1 $display("%b", po);
# 1  pi=207'b010000101101110001000010011001101111010110101010010000011111001001000001010001010001101011110111011111110100010100000010010001001000111101011100000111111101111001101010011001100000000110010010001000110110011;
#1 $display("%b", po);
# 1  pi=207'b000101100111011000011111001000001110111100010001110100010110100001110100010001010101111101100101000001010111010001011011101100110110111100100110111100010111110111101010000111010110110001011111101000101100111;
#1 $display("%b", po);
# 1  pi=207'b111000011010100111110000111000010111110110001110100010101101000111100010010000011010111010000110100011101101001010001101100100111010110000111110001110110000100000010101000111101010100110001011000111111000101;
#1 $display("%b", po);
# 1  pi=207'b111001110001110110101101111111000010010000101101110110101000010000011010000010111100011101011010010110010001011000010011100010001010101001000000000101001100110001101101001111110101010110001111110001011101110;
#1 $display("%b", po);
# 1  pi=207'b100010010101010001110110100100011011000010001101001110111010101000001100111100100100000011100101001010110110001111111010111010000011011011100111001000000101001000110100011000100000101000011000111111010110001;
#1 $display("%b", po);
# 1  pi=207'b000001001011001000000101001110101100011110010100001100011110101101101010011001001000000001101100101111010101000011011001000101101000110111000001010000001101000101110111000111001001010011001110100111011010001;
#1 $display("%b", po);
# 1  pi=207'b010001011011000110001101001000100100001101101101001011101000000110001111101010101100110111010100111001010011101011111100010110111000100111100110001001001010110001010011100000011001101001100001100010010000010;
#1 $display("%b", po);
# 1  pi=207'b110100011111111111001110110010000111101001011010011100011001111011001011110000000001000110111101111100110101110111010010011110011010100001001101001110101001011011100010010110101001011000010010110000101100110;
#1 $display("%b", po);
# 1  pi=207'b101010000110101010100001110100100010001111111110100011111110011011000011000000001100110100110011010010100101011110101001110000100010011110111111001001110000000100011110010101100101001011110010010110010110110;
#1 $display("%b", po);
# 1  pi=207'b100001111101101000110111100111011001000111011000001001100110111001110010100010000001011111000110001011111011000011000001101000011001010000011011000111011111110010110100011101111011110010001100010000111001101;
#1 $display("%b", po);
# 1  pi=207'b100100111111000000000010001001101100110010000000101100001100011001100001110010111010110000101101010001000010110001010110101011100101101011111100110001101100111101111101000011111100100000000001111100100111011;
#1 $display("%b", po);
# 1  pi=207'b001100100011100010100011001011111111011100110101100101011000110110110000110100110000010100000101000011110110101110011010001100001011011010001100101100011011110110000100001010010111111000000011111000000100011;
#1 $display("%b", po);
# 1  pi=207'b100001011111111101110100110100110000111111110000001110100101010111010100011101010011101110011001000111111101110101111000100110100011011110100001010010111100101110110011110010000110000011001001011001011100111;
#1 $display("%b", po);
# 1  pi=207'b001000111110010100001100011101010010110011010100101010101110011011010011100101000001011000101101111110000010101011011110101110010000110011011101111011110101100110111111111111100001010101110110110110110101100;
#1 $display("%b", po);
# 1  pi=207'b011110011001100110010001110110011010111001111110101100001110110010111101100101100001000101010001010000000100100001000000011001001110000100100110100111100110001001100000100110001010110110101000101000001110001;
#1 $display("%b", po);
# 1  pi=207'b001001011110110000010100001101000010111111110001111011001000001001111110110101010010101110011101101011110011000111101001100010111010000110100110010110001111000111001001011000100101100111010000010110010000010;
#1 $display("%b", po);
# 1  pi=207'b101001010111000011011011101010111011010110101110100111010000010100010110101000110011011100111111111110011011011101111010100010110110111010001101100000011111100000010110110100001011101000001000011011001100001;
#1 $display("%b", po);
# 1  pi=207'b100010001010000000011101100111111111111101010110011001111100000101110000101101000101111110100101101110111011001101101001001000100100100011101100100101100010100001001100010011011100010001101011111001000111000;
#1 $display("%b", po);
# 1  pi=207'b001100111011100010110001011001011001110010101010100011000001101100100110110010101011100110111101010010011111110111000100111100001110111110000100000001100011110001111000010101000100001011111100001000100001100;
#1 $display("%b", po);
# 1  pi=207'b101011000011010010101111111001010111101101001001110000110000100110010100101101111001101010011000000011000111001000110111010110111111101001110111000110100010101100000001011000000000101001110100010111110000011;
#1 $display("%b", po);
# 1  pi=207'b010110000101110011101010010011110101101101110111100011101010001010111110000101110100100101101111001110001101001010111011101100110010010000000111010000000010101110110000100111110000100001111100001011010100101;
#1 $display("%b", po);
# 1  pi=207'b000000100001110001010011001011010001010001001100110101011000100010000001101100001110010010010101010010011101111011010000010000011100011101101010011011010010001001000011100110000110100101110111111011011100111;
#1 $display("%b", po);
# 1  pi=207'b011110110110110111000101010011001011110101100111110011000111011111010111010100010010010011011001100110101100101110011011111111110000100010010001011101010011100010110100110000010011111101001111101011000010001;
#1 $display("%b", po);
# 1  pi=207'b010001000111010011010100011011110100010110010100111100100110010000101010101101100000000110110011011101001010101001101001011010001101000010001011101101001110101010011110100001110101001011111010001000100101100;
#1 $display("%b", po);
# 1  pi=207'b010101101001111111010000001011100111110000001111100001101110100011111110001001000100000010111100000110100101111111111001000001011100100010100110001101001001101011110011011000111101001000111000110000110101101;
#1 $display("%b", po);
# 1  pi=207'b010100010001000011111110110111101101110010011010010010111111100110100001101001000111111001111001100100011100001101010001011000110101101010010110001010110111001110010000001010100011010101001110110110111111101;
#1 $display("%b", po);
# 1  pi=207'b011110111100110111101010000001000000101111000101001011111111111100111101011001100101001100101000111011100110010010001011110101110111000000011001010011000110100000100101100100111100001110101010111000001010011;
#1 $display("%b", po);
# 1  pi=207'b010101101110100000110000010010000011010101110001011000100111010111101010111000010000101000110001001110111000111111101111111010000011110101000110110011111110000110000001000010110111110001000010000010101100101;
#1 $display("%b", po);
# 1  pi=207'b100001110110110000011010111001010110011001100100110011011000110100001110011100000000100110110001001111000100011001110010010011010111101011010111101001001001111100001011111100010100111101001011100111110110011;
#1 $display("%b", po);
# 1  pi=207'b100010011001101101100010000010101001001010010001001000111011110010010001010111101000001000000100011010110101001110001010010000100111110011010001111000010010110111111100001100111000110101101011010110111101011;
#1 $display("%b", po);
# 1  pi=207'b011100011001011111011101111100001010001111000111010111011011001100111000011000100101010101000101100111000011011110111010010010000010111010101111100011000101010011101100110010001101011011110001010101000011011;
#1 $display("%b", po);
# 1  pi=207'b001100100011100100010000001000100101110101100111011111101101010100101010110011011100110110001101000010000101100110001100101110110100010101001010110100101010000110110101100101010111110101010011110110000001001;
#1 $display("%b", po);
# 1  pi=207'b001000000000101101010101111111011001111000100100111100011101110101110000110000111001110101101010100001110010011101100000111111100001100110111110111000001101110100101011001110001100001000110111000010101111001;
#1 $display("%b", po);
# 1  pi=207'b111101110100101000010011110101110110111000000110000110110011111001001111110000111000000000100011011111110010010100100000101100011111111100100110100110110010001100111100111010101110101110011011000000100111101;
#1 $display("%b", po);
# 1  pi=207'b100010001000011001100000011001000000010010010001111011010110001011110110010100111111010111100101110101110001101010011010100110000010010110110000000101011011110110100101101110100001010001000000000110101010011;
#1 $display("%b", po);
# 1  pi=207'b110101011000000110110111000001101100001010110000001100011011001110111101110011101000001100100010011111011110010010000111100010100101000010101011010011101100110111001000100111110011100011101110000101000010110;
#1 $display("%b", po);
# 1  pi=207'b001011000010110001011011110111001100110000101111011011101100011100101110011101011001001101101110100101110000101101001011010011011110001101001001110010011111101001101100111010111010000111000101100001101101000;
#1 $display("%b", po);
# 1  pi=207'b100111001100000001101001000110000100010111000010010001111010100110000100110111111001011010010111101111001010100001110000110001111001011011001110010000110010000101000110111011111011101000011101111010001110000;
#1 $display("%b", po);
# 1  pi=207'b011100110010001110110110111011111011001000000000011101100000111101001101101010001010010010011001010101111000110111110101011010100100111001011111001011100101011110011011010001010100111101011101000011100001001;
#1 $display("%b", po);
# 1  pi=207'b010110111111101010000000000100111101110111110100100110011110101100000110111100011000001011110111011101010100110010111110101111111001000111001100111101000101011010100110001011101110101101100011011111001000110;
#1 $display("%b", po);
# 1  pi=207'b010110111001011010100100001100011111111000010000100011000110111001010110111100110011110001101110111101001010000010000110110010011100000100011001011000001101001100001101001100111011001100110011101110011110001;
#1 $display("%b", po);
# 1  pi=207'b011011001000001011101110101110011110000111100111100100011001101001000110110010001111000011100000101101101100001010100110000011100000111000010000011110110001110110010011011001011100111011111111100111010010011;
#1 $display("%b", po);
# 1  pi=207'b111111101010000011000110110100111100000111110010011011100111000001011110001011100011101011000110111100101110111001001001010110100011111110000000011110100000111101000111000001010011010010010001011110010010100;
#1 $display("%b", po);
# 1  pi=207'b010110100111100111000100110011000101110111011000010100100001111000100001110100010110111000101101110111001110010010110000100001100101000100100100011000111100100111100111101011001100001011111100100010000000100;
#1 $display("%b", po);
# 1  pi=207'b110101101001000000110110000100110111100101011110010000000011011110000101010001101011101001001110001000000011100111010010010000001111101000001101110111111101110011101011001100100101010011011011111101110111100;
#1 $display("%b", po);
# 1  pi=207'b110110001010001100110101111101110011101100010000011101011000000111110111100111010001000100000100010100010001110010000110001100000110111101001011111111001010000001010100011000001111010011000001101110111100100;
#1 $display("%b", po);
# 1  pi=207'b100110001101100101111010011010111010011101111011111101010011001000010100000100011111111011011011100111011001111001011110001110110001100010101111110111001111010101000000001011001100010011011100001111010111010;
#1 $display("%b", po);
# 1  pi=207'b000110110100000100111101100111001001001010100010110010101010010101100111001011010100010011100010000101011000100001110000101100001111110100101011010001111010011111011010100101100001110110110101100101001011000;
#1 $display("%b", po);
# 1  pi=207'b100010001010100111101101111011011100111110011011000010101110001111110011101100010011011010100110011100010100000111110111010001110011010110110011010000011001000001000001111101011011101111111000110101100000001;
#1 $display("%b", po);
# 1  pi=207'b101110010000101010110111010100100001000100101000100110011000111000101000100101101011000100101111000100100011001101111111001000010000000011011010101101101011100110011111101011110010100100011011011000001111001;
#1 $display("%b", po);
# 1  pi=207'b110110000111110101000010101010001111110010001100010001100111101101111001110110011100000101101000101010000110011111000111100001111111101001100001100001000011010011000000010111010110000100000101100110010010010;
#1 $display("%b", po);
# 1  pi=207'b110011111010010110000110110000011001010000101110000101010100111110000000001010100111101011100011001110110101111101100111000000011011011110001010110110111010110011101100111001001100001100000100001011000101110;
#1 $display("%b", po);
# 1  pi=207'b101011100000010101000101100011101010011101111110110100111010101001010111010011101110101110110011010101000100000001010010001001001100001001000011100000010000001100110110110010010110001101001001100101001010011;
#1 $display("%b", po);
# 1  pi=207'b100001100000000110010010101000111000000011110001010110110111001111101011111001010011110010010101100100011100100011111111110001110100110101101010100011100000001010110010111100101111110110000101111111010010110;
#1 $display("%b", po);
# 1  pi=207'b001001110011011110100100011111010110011011110111000011111010110000100100100110100000000000010001100111101010101001001111110011100101010000001000001011000100111011110101000101100011100000111111101101111101110;
#1 $display("%b", po);
# 1  pi=207'b000000101110101010101010011111010110001001111001000011001000010001011111111111000101101011101011010111011001101100100110100101100011010001011101011110101100110100110000000100000111110100010110000101001100011;
#1 $display("%b", po);
# 1  pi=207'b110110101110111101100111001000010010011000000100110010110101010001110011100100110000000111010110101100110111011011011100111110110001000011001110100001000111101111010010011010111011110001000000001101110011111;
#1 $display("%b", po);
# 1  pi=207'b101110001010001101100010111011011001010001000000101101111000011000001101001110000101100110100010000000000110110100001001100111010110111010010000101100111110010011101010100010111001000111011010001110111010110;
#1 $display("%b", po);
# 1  pi=207'b110011000110101101100010110011110010001101001111000110110011000110101010110100101000111001100110111010001110001011101100010101010010001011011000001101011010010100011001001111000001100001010010011100110101111;
#1 $display("%b", po);
# 1  pi=207'b011010001011011110010000001100010001101100111111010011011100111001100000000011110111110001011100101011001011010011101010000011001011000000001110111111001110001100001111100111111000101110010100100000010011010;
#1 $display("%b", po);
# 1  pi=207'b010011110101110111011100011000100101111101110000111100100011110110111110111111010000000010011000000100011010000011010100001010111110001100100111100001010000110001001100101011011001111010100001111001111011101;
#1 $display("%b", po);
# 1  pi=207'b110010110011010111110110101000110101111001001010111000011010111110011101101011100000110100001011001010010111111011000101110101001001011000110010000100000001100101100001101100101110110101010111001000010001001;
#1 $display("%b", po);
# 1  pi=207'b011000010101110111111100000100011011000110100010100100111101111000011101011101110111011111110000011000111011111101110111001011110110001111101101101011001100011111000101100000110110111000010101001100100111010;
#1 $display("%b", po);
# 1  pi=207'b101100001011101110001111001101000111100111100100010101111010000001001101110110001010011101010110001101101000100110111000100110000101111101111100010011001010010110100111000110111101101101110011110000101000111;
#1 $display("%b", po);
# 1  pi=207'b100100010111110001101011001100001000010000011111101010110101111110110010001100100111001110000011011000111010101101101101001011001011000011000111101000010001111100101100111111011111010101101001001000011010101;
#1 $display("%b", po);
# 1  pi=207'b011110001000010010101001101001111001010110000111011010000110111101101110100011110110000011010000000110111101001100001101001000001100110101001101000010100010000011011100100100011010010000100001011001010101101;
#1 $display("%b", po);
# 1  pi=207'b110110100100011101110000101001010000010010001111010100101101011101111011000000110000110000110110010000110101101000000000000000111111110000111111101011001100000110100110110000011101010110001110011010110001101;
#1 $display("%b", po);
# 1  pi=207'b000111101110111111011001010010111010100111011000101011111011000001100100101100111111000110100010000100001011001010110110110111011011110010010000000101111010000000110110110001000100111010011000100110111010000;
#1 $display("%b", po);
# 1  pi=207'b001101001101000100111010101010001100011000101001110010101110111001110001111011010000111010111111000000011110000001100100101000011011011010101100111001001100100010110101110100010001101101100011000101000001100;
#1 $display("%b", po);
# 1  pi=207'b011000100100011011011000010001111011011110010010100011100011110101000100000111010000100000010100001001110010001010110000001000000111100000000100001001000011000110111010010010011010001110010011001100100011101;
#1 $display("%b", po);
# 1  pi=207'b011010010110111000101101001101101010111101111111000111110010001111111001101011100100101000101111110001101011010110000100101010100110011000011010110100111101100010011111010100001110100110111011000100001111000;
#1 $display("%b", po);
# 1  pi=207'b111001010011000110001000110001001100011100010100001110001001110100010000110010000101100100000001101111111111011111001110000010101110100001000101110100100100101110010011011010000010100001110101011100000111010;
#1 $display("%b", po);
# 1  pi=207'b100011101001001110010000010010111100000110010100001011001100111001100000001011101110100111110011001000101011000101110101101000001100111100011010010001010001010110111010000110001010000111010000110011011100000;
#1 $display("%b", po);
# 1  pi=207'b101000100100011001100010010000010110010100000110000000001101110101101100011110011111111101110001011110101011000101011010110100010001011100100110010100000100100000010000001010011111110111111001101111001100111;
#1 $display("%b", po);
# 1  pi=207'b011000111110111011110001111101010001100101011101000111000100010000101111000110100011101000001110011100011011011000100101110101010111111101011010101111010100111100000101111111100010010110101000001111000110011;
#1 $display("%b", po);
# 1  pi=207'b101010011010001001011000111000101001111110111000111011100110100010011111010101010100000000001011111111000010110111110001100001101100110101110011001101110111010111101001011000101111010101000110000011010101001;
#1 $display("%b", po);
# 1  pi=207'b101011000001011000010101011011101110111010000111010001010101101100011100101111001110111100100100000000101000011000000110010111000000010111110001000011000010111110110010100001001110001101101101110101001111100;
#1 $display("%b", po);
# 1  pi=207'b010010110110001010000111111011110110110001101010110011001001101110110100011110111101101011101001010111110001110011010000100110001111101110010010010010101101100111110101110101110000111101110101000010000001000;
#1 $display("%b", po);
# 1  pi=207'b011000100100000100110101000100101001101111001111011001110011010010000001110000000000001010100101101110100110110101010001001100010111011111101110011010010001110100000000110010100110111100111011001011100101001;
#1 $display("%b", po);
# 1  pi=207'b110000011110111010011001000010010110110001011101011001111110000111100110010100011010010111111001000011101010101000100011010001111010000000010111011101001111001001110110111000100111000001000111111001101111001;
#1 $display("%b", po);
# 1  pi=207'b111010110001000110001110101010111111101000000100110001100110110111001110100010110011000011000000110010101101110011001101000001101111010111110000100001001111011011100001001001111010101011011110011010101111000;
#1 $display("%b", po);
# 1  pi=207'b010010011110111111101101001100111111000001011111110101101001001101001000110111101110001101010011001010110110111100001000111110011100100010011001111001100100001001110100101000011001011110101101101011001010110;
#1 $display("%b", po);
# 1  pi=207'b101111000011101010110001001011000111000000101001011011010000110000001001100100101100111111111000011011001110101111110100110000111000100101110010100101001001110010110000100011100001001100010001011011101010101;
#1 $display("%b", po);
# 1  pi=207'b001000111001110011001010111001111101101111001011000000000100110111110011010101101100010010110100010010100111000010010100000101111010101010011001011110110111011110100100110011111111011110011010100010111000010;
#1 $display("%b", po);
# 1  pi=207'b011111000101100011010001001100010000100101101011100011111010010111011101011101111000111111110101100111110111000000100001010001100100100010011110010000010111100010101011101001111111110010110000100001001101010;
#1 $display("%b", po);
# 1  pi=207'b000101100110100110110111001000011000000000100101011110101000000110010110110110100000010101011100010101011010101010001100011110101100000110110111000001001000001110100001011100100011111101111001000110101011101;
#1 $display("%b", po);
# 1  pi=207'b100110001011111000010101000101110001110001110110100011100001000101111010000111010100010110000101011001000100011000011111101111000100000000010010100100111110000011000011011100111100100101010011011001010000110;
#1 $display("%b", po);
# 1  pi=207'b001110100110010101101001011100101110010101001000011011101010001101000100101110010111111111000111000100100010000111111001101000010110010100001100111110111001100101000010001000010010110001010101001011101010001;
#1 $display("%b", po);
# 1  pi=207'b000101100111010101101000111100100011110001001111100001110110010011100000000100010000101010000100110100101011110110110000000001010010101100101001000100001011100101101000011100110110101100111001010101100001001;
#1 $display("%b", po);
# 1  pi=207'b010110101110100110010011110111000111111101000000111110011000111100010000110101111110001010011001011101000000011110011011010111010110110010101000001010101001010000000111010100011100100010010110011000011111000;
#1 $display("%b", po);
# 1  pi=207'b101101101101100100111101000010000101110110111001000110001011000100100010011111000110001001101000011110001001111010001010001111111101101001110111101010101010111000111110110110110011100010000011111100101101001;
#1 $display("%b", po);
# 1  pi=207'b111000110010110111000111001010010010010001000010010111110101010101011100111100010010111011001101000101011110111110101100100100111101000010110010100111001010100110101111100000001111010011001101110101001110101;
#1 $display("%b", po);
# 1  pi=207'b110111011000101000110110001001101000010011110101111010011100111101100101100001011100111000100010011100010011000111010111100001010011010100110000011010101011000101110110001000001100010101011111100011101101111;
#1 $display("%b", po);
# 1  pi=207'b101110010111001010001001011110110101101010010111110111001101011000110101011011001111111000001001110100111010110101110010110111001010110110010011100010100110111111010011001010101100010011101010110010010000110;
#1 $display("%b", po);
# 1  pi=207'b111011011010000000101101111111000000010011100010001000101000010010110000000100100110011000110001010000100111100110111100100110100101001100010000111010000011000110010111000100111000111000010010010101011101101;
#1 $display("%b", po);
# 1  pi=207'b111110100010000110000010000010101001101101001010111001111110000010001100100110011011010111010001110101001110110111110101100010001111001000000010100110101101001001010011100111111110110010100100010011100110000;
#1 $display("%b", po);
# 1  pi=207'b001011010111001010001011010001011111010000000110100101001101100011111101010001000111100001101110011111001110110011100001100101101001001100110001010001101111010001000011001011000010011111000100100110110001010;
#1 $display("%b", po);
# 1  pi=207'b010110110100011000110111110000101111111010111011111001100001100110100101000110101100000010111010011101011011010101101011100101101011011001110111001100010010100111100111000110000010011001100100101100000001110;
#1 $display("%b", po);
# 1  pi=207'b011111001101111011110011110111110010010000101100010001011101101110010010110011111111110101010010100000011100101000110010101000110101011110000010010110001010100100110001101111001100001010100111010000010001110;
#1 $display("%b", po);
# 1  pi=207'b100001101000100110111101110111100000111101100101101110110110000001001101001110010011000010000000010111011111010100111101110110110100111000011100011110110111011000101101001001000000010101111011011011010110001;
#1 $display("%b", po);
# 1  pi=207'b111001001100010100001011011110110000101100010010100111101000101100011101010101010101010000100000010101010101111110010111100100110010011110000010100111010100011000111010110101101100101011011110001001110110110;
#1 $display("%b", po);
# 1  pi=207'b010100001100000111010100110110100000010100000001101011000001101000110101101011100101010101001001111001101100100000100000110010100101011000000110100010001100101001100010111000010101011001111111111111010110011;
#1 $display("%b", po);
# 1  pi=207'b011011100001100001011000011100110100010110011101100000100010001111100100101000011001001011111111011100000100000100000111010000110111110000000101001111111000111000011011011101100110111101010000101110110110000;
#1 $display("%b", po);
# 1  pi=207'b001111100110000000000010001011101110001100101010100011001011010000101110000001000111100110001101101100010101110010000110100101100000011010110111010110011110010011000001010010111011110111001011110101101000100;
#1 $display("%b", po);
# 1  pi=207'b101000100000110000100010111000110101110011000011010110011001111111000100111100010000100100000110010110000100001111110111100011110010001010101110111001010110011110110010000100001101010110100100000101001010000;
#1 $display("%b", po);
# 1  pi=207'b101001101111011101010010001001111001111011010011011101010101100100100100011011110100101110001111001011011000001011001110101101101010111010010001111110101101111111111101011100010101011111010001100111011001000;
#1 $display("%b", po);
# 1  pi=207'b000100111111111011001111000010010111000110000110001001101100101110001101111101000011110111110001110001001101011000001100110011101101000110000001111101001111100100010011101011000111001110000001001011010011101;
#1 $display("%b", po);
# 1  pi=207'b110110010111101000111010110001100100110111100001101010101100001101011010001100010011001000100101111001010111100101100011101111110110001111011100000001001011000111100010110001001110101101111010001011000110010;
#1 $display("%b", po);
# 1  pi=207'b100111110000001110100101010101010100100100011000101101111110110100000001001001100111101111000111101110000110000011110011010000101011100110000001111110000010011001000011001101001101001111101000011010101110011;
#1 $display("%b", po);
# 1  pi=207'b110011100100101011111000001110010001011110001111000000000001011101100110010110111001010011110101001001001001100101101100010101000010111011111000100110100101001110110011001101111000000001111110111011011101011;
#1 $display("%b", po);
# 1  pi=207'b000001000101101011111000011110011010001101101100100110000000010101101001111100000100101110111111100000001111000110010010110100110000100011000011011011011100000010100100010101011100000011111110110001010111111;
#1 $display("%b", po);
# 1  pi=207'b111010110000010011011010010100010010111110001101010000000011011100010101010110111000010111010010101111000110100010101111010111101001010110010011010111100000110110001111100100110010110101110101011101111000101;
#1 $display("%b", po);
# 1  pi=207'b001100100011111011000100010111011010101011010101111010111101111111001001100111110000101101110111001001111000001011110111001010110010001010110010101101011011010100111000111001100101101100101100101001011001001;
#1 $display("%b", po);
# 1  pi=207'b010001000100001011010001000100001101001010010011111001101111011110110011111101010111000100110001111101011001001100111101001100001011100000101010100100000010000110000100011100110101001101100001010010000110101;
#1 $display("%b", po);
# 1  pi=207'b011011010010101111000001110011100011010000110000110100010001100011100000001001010100010000101100001011000010101011111100111111111111110100101101000001110010001111101000101010011101111011010001101010010100010;
#1 $display("%b", po);
# 1  pi=207'b010101110011000000100000111110101100111011100001011111011000010000101110101100101001010101010111101011100111111011000000001100010101100101111110010101100010110001111100110101010000001100010010000000101101110;
#1 $display("%b", po);
# 1  pi=207'b110111011010000101101000110110101111100000011000101111101110110101011100011100010100110010000100111000101110100110100001001100100010110001101100111000101011100011101011110110111000010011101000100000111001011;
#1 $display("%b", po);
# 1  pi=207'b001010011110000000011110010011101011100110010010110100110010000110110100010010111100100010110001011001010001010011111101010011101011110011111000110110110010000011000000111010011111111100100001111011001100111;
#1 $display("%b", po);
# 1  pi=207'b110000001010100100000111000001000100010001111110001111101110000011111111111111011010111101101011000001111010001001101111100110010010100011110111100111100101000111011111100000100010101110001010000100101010101;
#1 $display("%b", po);
# 1  pi=207'b110011111110010000101001011011110000111111010111110101110000111000000111011000101111101101001001100000110001010110011110011001111010100111011011000011111000001000001000001011110010110111011011011011101101100;
#1 $display("%b", po);
# 1  pi=207'b001011111000001001000110101011001010111001000011000000101101001001111100100000100101010101100011111001111111101001001111110011010001100100010001000000110101111101110001100101100111100001001100101101100100100;
#1 $display("%b", po);
# 1  pi=207'b010001111110110010100011111110000001011001110100100000000010110001101011000011101010101101000110110010110110000111011100000011010000101100011011000100010000100010001100000100100010011010111111111110000110010;
#1 $display("%b", po);
# 1  pi=207'b000000011111100011011010000101001001011011000000000011011010010110100101000110000001011101100110000100001111000110010110101110011100100100111100111011101011100011100001100000111010101011010001100010110000001;
#1 $display("%b", po);
# 1  pi=207'b000100011111000011000101011110101001110100101100100111111100001010001010111101110000100001111001000110100001100010000100111110100111001111011110011110010100110001010011000011001011100010010010110101000001101;
#1 $display("%b", po);
# 1  pi=207'b010001000110001011101001000110101101110101000000011100111010011101010110101010110010110101110000111100011001100101000111111011000001111010000111000111010111011011110111000010010011001101011111100011110100011;
#1 $display("%b", po);
# 1  pi=207'b011111001000011110111100011001100111001111001010100111101001010110111001010101111001010100111000000101100100011011101111010110001000011111101101011001010000000010000011111110000000001000101000001110011100101;
#1 $display("%b", po);
# 1  pi=207'b111001010000101000110100111111111000001010001111010010100110010011100111010100101000111001001110110011101100000001110100011001110100110001001001000110111011000111101001000101101101101111111110011100011111100;
#1 $display("%b", po);
# 1  pi=207'b111111001001101100001110010011111000001000100001111110101101011001100001001111110011011000101000011011001101010001001000000101011011000111100010101011001110111111010100001100110100011010000110101111001101111;
#1 $display("%b", po);
# 1  pi=207'b001101001100100010111001011010011111111000011100100100001001110101001010000100011011110110011010110101010111010110000110100010100011001101101100101000110010100001011000001100111101111010000001000101110100100;
#1 $display("%b", po);
# 1  pi=207'b011000000011111100001110001001110100111100100111000100101110110011100111010101111001000100111000010100010101000101111100101100111000011000100100110100011001110010110100110101011011000000010011001001010010111;
#1 $display("%b", po);
# 1  pi=207'b011001010011111001100110100100001110010001011110110100110101000110110111101100000001011011011010101110010010110100100010000001100110101001011001101110001100010100010000000101100110100110101110001111011111011;
#1 $display("%b", po);
# 1  pi=207'b100110011100010000110100001010111110110010010101000001000111011011110001001010110111001100110011010001001000000011000001110100001111001100011101101001010111100101011101001101101100001101110100000010100010110;
#1 $display("%b", po);
# 1  pi=207'b111100010001000101011101100011000111100001100011110010100000010100110010010110110011000100101000001010000110001010011110111001010000110101010101100000011111111001100000001000101100010110110110000000011101101;
#1 $display("%b", po);
# 1  pi=207'b100111110001111000110110010010000100101011101111111111000101000010011101101111001111100101011011011011100100111100100100000100111011110101110010100001100111100110110010111111101101101000101010001101011010001;
#1 $display("%b", po);
# 1  pi=207'b111101011100101110101001000110001110000000110010001100010100111101111010011100111000000010101111100001101100010111011110011011001100010011000110001111010100001000111011111010111010111010101110001100110100010;
#1 $display("%b", po);
# 1  pi=207'b100011101100110010110110010100011111101010110010000001100111110101011111000001100110100011010000111010111101000010001111100000011100110100101000100101010100011101101100101001010000111111111001111000001111111;
#1 $display("%b", po);
# 1  pi=207'b001010101111111000000111111010110110101000101000110100001100101111100010010101100001111101100010101101011110110000001010101111010111111000001010010100001111010001101010001110100101000011010000001011011111100;
#1 $display("%b", po);
# 1  pi=207'b100101101101000100001011001010000000000011000011001100101000100100100110011100100101011101001111010111110110101000001101110110000010011100000000101011111101010100010000111101000101100111010010001001110011000;
#1 $display("%b", po);
# 1  pi=207'b101000101100011111010011011001001101000000100010010111110001100010101100001101010000100000000110000110010000000111101001100111110110101100000001101011100100010011001111011100110110001100110000110010110110010;
#1 $display("%b", po);
# 1  pi=207'b001100000010100111011001010100101011000111111110011100111000011100110000101110010000000111000010100111111011010011101011001000110110101100110110001000010110001111010110111011011100011011001010001111011110101;
#1 $display("%b", po);
# 1  pi=207'b110111000000000010110100000111011110111111111000110011111010001100101001110000010000111001100101000111111111100100101000011101100000010001011100100101100000010101000000101010100111111101010001110000111001000;
#1 $display("%b", po);
# 1  pi=207'b011010101000110100011010011001101011000111011110010000111000001011100000101111001011010011011010001101011110000110110110011111000011011011111101011110001010110010111111010100111000101010000001101101110000000;
#1 $display("%b", po);
# 1  pi=207'b000010100111001111110110000111001111110000110100111010001101000000011001111011001111111001010110001100001101111111110111001000011111111111100100111111111010111111101001110110000111010001001000001011100000001;
#1 $display("%b", po);
# 1  pi=207'b101001000100110011101110011011101011011001100011001011101110001001110110111010011000110101010100001110000000000100100000011011100010110010001000011010000100110011001111110110000000111000011011011011100100111;
#1 $display("%b", po);
# 1  pi=207'b011100100111001100110100011110111101010111110011110110011010010100111010101110110100111000010001011011001011010001101101010010101111110101111100110011101001001010110001010000111011110011101111100000110000011;
#1 $display("%b", po);
# 1  pi=207'b101010101100101101001010111001011110100111001010100110111110111001010101010100111000100011110001111110001000100011111101011100011011100010011011000110101011010111010011000100100001100100011110011111100010000;
#1 $display("%b", po);
# 1  pi=207'b111011000010001011011100001110011110110010010001011010010111100110100101101001110101010100000011111001001000110110101001010010101000110001011010010101011101100111011011000100100100101110110010000000111001000;
#1 $display("%b", po);
# 1  pi=207'b101001111000011000000011110100010001100011000110011110010000010100110000100110111000010000000000100100110011111011011011010011110000101101100100011011110100000110101001011100010000100011011010110011100111110;
#1 $display("%b", po);
# 1  pi=207'b110101100001101100101010111111100110101110101111010010110110001110001101000000110100100010101000000110110001000010111100011011111110000110000100111111110010011100010001110011101011110010111110111001101011101;
#1 $display("%b", po);
# 1  pi=207'b001000101100011101101101011000000110111010111100111100101010000100000001010110001101100010011001101100100011111001000010101011100100001001000010101011010000001101010011011000001001100111010010111010000000111;
#1 $display("%b", po);
# 1  pi=207'b000111101000101101001011100011100101101100001011111010110110110011100001110010001011111001001110101111101101101101111110110110001000110001000110000000001010101110011000100001101100010111101001010101001010101;
#1 $display("%b", po);
# 1  pi=207'b011010110001101010011001001101100011110101101000110100110110011000101100111100010010110011011010000101011001110010011001010011110001000100000010000000010000111000101001100111111011101111111010010101111000010;
#1 $display("%b", po);
# 1  pi=207'b000000010110011001111000110100110111100100110110000001010001111001100111000001111011001000000011110101010000000001010111100010110110101010011010001001001001001000110011110001101011110101110111011110011100100;
#1 $display("%b", po);
# 1  pi=207'b011110010000010011010001000100001011010010110000000001100101111101000101101110011101101001110010111001101111000010101001110111000010001101101100001100101111010111010001001010100100100110111001110101011110001;
#1 $display("%b", po);
# 1  pi=207'b000101000001101100110000001010100001101100011000000000100111010101010100101110111100110111000001111000110101001001000110100101111111010110000101010011100001110011010110010101111001101010101110010011000010011;
#1 $display("%b", po);
# 1  pi=207'b000011101011110011100100111011110001111001100011101010110000000011000100001010001011011010110000011110110000000011000001110011000011010000110010010100010100001101111111101011000100101101111101110110011111001;
#1 $display("%b", po);
# 1  pi=207'b111010110110101111111000111101110011011000011111101101011101111111111001100110110001111111000011010000100001001111100001111000111000101011000000101010111110000000101100101110011100000001011101001110110111000;
#1 $display("%b", po);
# 1  pi=207'b101010001000000101000110111011011111101111000100111010001000010110101100011100010111001010101001111111001100010110101011011010101111100110001001001101011000011000010011111000111000011010010110101101010101111;
#1 $display("%b", po);
# 1  pi=207'b011000000110111000100000110011011110001100011101011000001110011110111111111111010001001111011110001110111010111000110001101101110110011010010111010110111111001010001011010010101001111110101010010110011000101;
#1 $display("%b", po);
# 1  pi=207'b001111111100010101010101001110110111110001010010111011111110110001001011000100100111001011011001000011110110000011011111010100110111111000011001110101101100010000001100000001111111100110001101010000010100111;
#1 $display("%b", po);
# 1  pi=207'b101101011001100010111010111111010010111010001101000111001011001010000110100001100001000000000010010111000000000000100001100100111100110001000001001011111110000011101010001011101101000000001000101110010100010;
#1 $display("%b", po);
# 1  pi=207'b011100010001000110011101110001010010111011000001001001011101101100011100011101011101000110000110100100011101001101000111001000000010011010010010111000000010010011001101001100010011001101000111010101101011001;
#1 $display("%b", po);
# 1  pi=207'b001001000110101101000011010000100100111111011010011111110100110000011110011000111001100011011011100110101110111011011010010010100100101000010010110110111101110110000110000110111011001000010000001111011111110;
#1 $display("%b", po);
# 1  pi=207'b110010010110011101000010001000110000010111101111000101111101011000100010000010110000000110010001000000110110110100000111000010111101000001000011001000110010000111001010001001010101010011111101101101010001011;
#1 $display("%b", po);
# 1  pi=207'b010001010000111100111001010010101101011100010011010001011011110101000010010000001010000110100111100010011111010011010100110101101101001111001000110101110001100110100010110100010011111011011101010001010110100;
#1 $display("%b", po);
# 1  pi=207'b110110000011110111011101101101000001010001001011000001001011111010101010110100000000010011011000001001010110000010001001010011100100100010010101111110000011001010010001011001010100100111000011100010111001001;
#1 $display("%b", po);
# 1  pi=207'b110011011111000010000100110011110000100010000100111010101100101000010000000100011001101010000010001001100101111110110001000101001001001111001101101011100000000111000010111010100110101101000101110100000101001;
#1 $display("%b", po);
# 1  pi=207'b111010111111101101011101111111010011011101100011100110100100011111110100010000100011101011001011111100101101110101101101110100101010010011000111111100110011011000001110010001010010010011111000110111110011001;
#1 $display("%b", po);
# 1  pi=207'b001010000011101001111001101000100000000110011110100100001100110110111101101010010110111000111010010100000101110110011001000101010000011101110010111011100000110000100011001111101000011011000100000100101100001;
#1 $display("%b", po);
# 1  pi=207'b101001000100101110110011000011010000000111101011000111100101111011011001110100110001000111000101010110110011010101010000011001001001000010011011101101010111000111110101110000111100101110010010110111110000000;
#1 $display("%b", po);
# 1  pi=207'b100101111001111111111101000011000001110110000101111101111011010111000110010110011001000010101111100100101100110111011001101001000011100100110110110100010110110011100100011010010111101101011001010010010001110;
#1 $display("%b", po);
# 1  pi=207'b110110110000000000100100000100100110000000100011100110011110101110011100110101101011001000001011000111101010110011101010001101110110111000001100100110011001111110111010110001010001101101010110110101010011101;
#1 $display("%b", po);
# 1  pi=207'b001011000001010000100110110110010001011101010100100011101001010000001011100010010100000100111110000100110100100100000101111100001101110001101100010000110110111011101000111001110001110001011110011010111010011;
#1 $display("%b", po);
# 1  pi=207'b101011101010001001000001110011010111101011101001111010100010000110010111100101111001101000111011101100110000011011011111100111101101000100001111111100011100110111001001000011001000000110010011111111011100110;
#1 $display("%b", po);
# 1  pi=207'b101101111101111100010000010001100000010100111111110110101110111011110000111011010011010011011000000110010010110110001110100000001101000001001100011011000101010001000110001001111001011101111000101000000110101;
#1 $display("%b", po);
# 1  pi=207'b001100100100101110110111001100101111110100011101100111110110001100001100111011001010010000000011010110000110100101100101000101101010001100100110100101110110110000011100000011110011000000110111111000101111011;
#1 $display("%b", po);
# 1  pi=207'b001101010101000000111000011111101100110111110010001100110001011001101111000010110101001110011110010001011110000011011111110001001011111100100001011111101000111100011100100100100011010101011100000001111111010;
#1 $display("%b", po);
# 1  pi=207'b100101101010010111111010011011110110001101100010110100011101000100100101111001111010101100100011001100011010001000000010010101101101101111001011110111010110010010110111110000101110011101010011010111010110000;
#1 $display("%b", po);
# 1  pi=207'b101101111000100110111100101110001101111011111100111000000000001001010001010010001110010000100000101101010101011111011001010100011010001101110110110011110011010011010110011000000001101011111100000110110010100;
#1 $display("%b", po);
# 1  pi=207'b101000101010011000010101100110010110101111011110101101010111010100111100010111101011111101011010001011001111111011100000101100100101100101010001100000110011010100000010100010111011110101100011101010111101111;
#1 $display("%b", po);
# 1  pi=207'b001100111001110101011001100111100100001000011010111011100011010100100100110110100000111100000111111010001011000010010111111011010101000001100010110011011000101000101111110100000011111101011011010001100101111;
#1 $display("%b", po);
# 1  pi=207'b101011000111011101010111101100111001000111001100010010101001000110000101000010111110101110111100111000111101010001101010110110010001111011000110101001011111101010000010100100000001011000101100011000111000111;
#1 $display("%b", po);
# 1  pi=207'b000010111010000000000001100110011011000100100000011101100010001100000111100100010010010111000101100000101110111101110110101000111010001011001011001111011111000000000001010111010101100100100011101111111000011;
#1 $display("%b", po);
# 1  pi=207'b110001101101001100000001111100010101101100001010111110011100001000110000000111001010011011111000001000000010111111101001000100011001010011011101010000111100101111011100101100100110011000001101010111110011100;
#1 $display("%b", po);
# 1  pi=207'b000111001010011001101110001101011010000111100100110100001110000010100000010111101001101011110000000001101010111001100010111001000110101111110110100110001010110001110110111001000011011010001000010111001111111;
#1 $display("%b", po);
# 1  pi=207'b001101011101101001101111111110101000000010000010111000101111000110000110100110011101001100111100100100011110100011111100111100000001111001000100111110100111000001100110000010101100110111010110010010000001000;
#1 $display("%b", po);
# 1  pi=207'b101101000010001110010011110111010010011101101000100000001011011110111101011000011101000001101110101101010010110110101010010111110100101101011100010110011001110110110011101010110100001010010011001000101011110;
#1 $display("%b", po);
# 1  pi=207'b101010111010100011101100001010011010110100001001010101101000011111000000001100111101010100010001101001001101010011011111001011001001010001010111110111100110011001100100101100101110110111010100001011101111000;
#1 $display("%b", po);
# 1  pi=207'b111101111100010110000000111011000101111010110011110001000010001010001101011111010111000010101010011001011010101101111011101101101011111101011110110110011101000110100001110011001010000110100111111010000010011;
#1 $display("%b", po);
# 1  pi=207'b110110011001111001000101000011111111110111001000110110110001011001111100000111011101101111101000100000111000101010001101110101011111001010100110100110100100110100100110100011011100101010110111000110100110001;
#1 $display("%b", po);
# 1  pi=207'b000000101001011100000001010111011111001010110111011001101000110010100001010010100111100110001011100000011010100110010000101110100000110011011111111010110100100111011100111010001111001001111000001000001001010;
#1 $display("%b", po);
# 1  pi=207'b000000111011001001110110101011001111011011010111010101000110011111001010110110000100000111001000101010000001110101001001111000110000110110000001100110001000101100011010011111000100001001101000001001100101011;
#1 $display("%b", po);
# 1  pi=207'b001100010001000101000111011111111101101110000010000100011010101000001001011010100011001011001001100010111110011110101100010001011010100000100010100010001001111011000110101010110110000110011011011110100111011;
#1 $display("%b", po);
# 1  pi=207'b101101011100001111000001111001001000111101110000111100010001011011001000100111011111001001011010010000001111010011010000001010110111011010111001110101110011111111110000100001110011100000011001110111011100010;
#1 $display("%b", po);
# 1  pi=207'b000011100101110110101011010100100110001000011110011101110000111001100110111101001100100111100110010111101010110110110110011111101110011011111111001000010100100000011010011101000000010011101010010001011001000;
#1 $display("%b", po);
# 1  pi=207'b111100011110111010011010000101100011001010010010000111111000001110100111001001010001000000001101110101100110101001111010001000111111011010100011110011111010111011011011011111100000101010110001100111000100011;
#1 $display("%b", po);
# 1  pi=207'b010100101001010000001101100101011000011100011001110010111100000001110000111011010101110100100001101001111001100101100000001001001101101100101001100001001001000100011110101110101011101110010010000100101000000;
#1 $display("%b", po);
# 1  pi=207'b001010101101101110011001011001001011011010010101011011111111111011111000101001000001010101011000010100011000101110000110001111110001001000110101110011000011001101010101010110010110100111001010101010001110110;
#1 $display("%b", po);
# 1  pi=207'b101101110101110010101111111111011110011000001111000111000110110111111000110110111101011010000001001101010010111100111011010011011110011101111110001100010111011011110110000110101001111011100101001101000111100;
#1 $display("%b", po);
# 1  pi=207'b111111010101101100011110011110110001010011010011010100110100111011010001001111101110010100110011011110010011011000111110010100010000010111000001100110001110100111001111111101001100011000010100001101010110100;
#1 $display("%b", po);
# 1  pi=207'b110000110100010110101111110011001000001101000111100100110000111100001011100101010101110000101101100001111001101010011111111000000001111110010100001001011010011010010101100000011100101110011110000010011001000;
#1 $display("%b", po);
# 1  pi=207'b001110101101010110100011101001000100110010011010101101111011000111010110001010011001011011111001111101011110101000011111101000000011101111100101001100110110100011000011101011011101010110000100011100100101000;
#1 $display("%b", po);
# 1  pi=207'b011101000100111000111000111100001110111010011110110100011110111011010101100010000101110000101110111001111010101101011000010100110000111010001110101000000101001100110101101000100010011101010100110100100000100;
#1 $display("%b", po);
# 1  pi=207'b000101010111110011010001010111000101111010111010010010101001110011110101100101100111000001111000010110111111101001011110001100101000001011100011101111101001101001111011100110000000100100001100110010000101110;
#1 $display("%b", po);
# 1  pi=207'b000101111101110110101000001100000111101111110110001011101010100010000010011011111101111111010001000000011111000111101100010110010010010000011010111101111110011110000111001110001010000100001011010100111011011;
#1 $display("%b", po);
# 1  pi=207'b100100100110000011111001100100110101110110101001110110110110001010010000110001111111111111011100100001110011000000001011100110000011010100000010110000000000010011010110001010011100010000000100101000111101111;
#1 $display("%b", po);
# 1  pi=207'b100100010001101101001101010111010110110010111111001001010110001101011101110011010101101011001101110001001100010101000100101100010000101101101101010100101110010010011110100010100000100001000010110010000010101;
#1 $display("%b", po);
# 1  pi=207'b111010001000111010001011000000111111010010101000101111100001010011100010011100110011001101110100010001100110101100000000011001001010101101110000001100010110010111010100010001000111100010110111000011011010111;
#1 $display("%b", po);
# 1  pi=207'b000001110010010111011001000011111011001110111101111100011111000110100000000000010000101010010001001000011000011101011111011000001010011011000010010111011100000000100110011111110010000101000111110010000001011;
#1 $display("%b", po);
# 1  pi=207'b110111011010010011001000010010110100101101011001111011011110100000111000010000111101011010100010110110000101101111000001011100101111100001111000110100010100001110101000011000110111100110110101110110110111000;
#1 $display("%b", po);
# 1  pi=207'b000101000111000010110111111101000111010110111000111000111000001110000101111100111011001110001001110011011111100100001100000010011010100101000100101001110001010101111101111111011000011111100110111010100001111;
#1 $display("%b", po);
# 1  pi=207'b001100101110111110101100110101110111000100001000010001111110000000100101110010110101101110100111000000011101100101001100100000001000101000000111001001011011001001101101000010001000100111101011110111011010100;
#1 $display("%b", po);
# 1  pi=207'b000000011101110001001101100000101100000010010011101000110111100001110010001001000101011010111000111110110110010011100100000011110011111011100110100001001110011111011100010000011101101000000100110101101101101;
#1 $display("%b", po);
# 1  pi=207'b011000100111110010101000111110110010011010010110111010100011000110010111100001010111000000011101111100100001101000010011001111110010110101110011101010011110101001000000101100010111010100000100011111000001110;
#1 $display("%b", po);
# 1  pi=207'b111110010111110000100111001001111001010101010110111101101010110000101110001110000100001010100000001110001000011100111011100100001010110000110110010100100010101101100000110111010101100100001010011101001111010;
#1 $display("%b", po);
# 1  pi=207'b101111110111010001011110100010000100101000001111110001011011010001011111101000100100110011011111010011100101111011010010101100001111011100011010000001010001110001001000100101000111001011001111001111001110000;
#1 $display("%b", po);
# 1  pi=207'b100101101100000000010001100100100110100100101000111011011001001010100101110101111000100011100011010000000101000000111100001000000111110011100010100010100110001100010111001001000111100110001010011001111010001;
#1 $display("%b", po);
# 1  pi=207'b000100000000111100000011100011000111101110100010110100101001011010111011101101101011010111001001010000000101010110111100000000110010100101111110011111111011001000110101100011011010000111000010010010011110000;
#1 $display("%b", po);
# 1  pi=207'b100101101000110000010101010100110101110111110100111000000000110011011001000111110101111100101010001011000100000110111010101100101110111101010100000010110010110001110111110110001011010101101111100010101101001;
#1 $display("%b", po);
# 1  pi=207'b110011110001011010011110111000101110010110111000110101111111000111100100011010111111111101001011111101100000110101100011000100100001001000011111100110001011000100011010110101000001001100010011000001011011101;
#1 $display("%b", po);
# 1  pi=207'b000101001010010111011101001000011111110011101111001100010101000111110011011111101101110011101001001100011001101010100100000001101100000011010111010111100110010010011010100000110000010100011101001101111010111;
#1 $display("%b", po);
# 1  pi=207'b111010101001100000000000000110100110001011101000101111100000101110001101010000101001001001111110011110000110110011011011111100100111110100010001000001101100000111001101001101011110111111100001100001010110101;
#1 $display("%b", po);
# 1  pi=207'b000001110001100001111111110011111000101010010111010000100001100110110110101001111101100111000110000011101111000111101010011001011010111101010010001100100001101100111001110111110110010000101101100000110101001;
#1 $display("%b", po);
# 1  pi=207'b111010100110100101010100011011011011011011001000110000011100011011111100010100110101100111000011100101111110100111000010100001100100000110101101011011010101100000001010101010111001001100000111101010010000001;
#1 $display("%b", po);
# 1  pi=207'b110011101111110111111101101110001010101001001001110101000100100100000011110001010000100001011100000000001010101111001101111101101010111001010001110110111110000110001001000111011001000010001111010111111010100;
#1 $display("%b", po);
# 1  pi=207'b111001111100110010101110100100111000101101100100000111110100001111000011000111101010110100111001001111110000000001101101001100101010001010000111000001101110011110010001100010010011101100100101011110110101100;
#1 $display("%b", po);
# 1  pi=207'b101100111101101010000100100100100100100111011010110000000101011111011010011001000101001010110100000101010010010000110001010100010001100100001111111110110101100010000111101110100100010001000011110111001010010;
#1 $display("%b", po);
# 1  pi=207'b100110101000000111010110011100110001001101101111111111001010100000100110101000000000001001111111100001011000011000110101000001000010111011101110100000110111000000111101101000010000101011010001110110110101100;
#1 $display("%b", po);
# 1  pi=207'b110100100101000101001111111011110010110000000110010111100000100000110001110110110000010001100011110110001011101100111001001011001011010001101001011000110001010101011010000011110110100001111111110111111101000;
#1 $display("%b", po);
# 1  pi=207'b100100111100101100011010111011100001011000000010001011000100100111100010001000101101101111100100010111111001111111010000001011011000110001100011010101111100101101110000001011101110011011110011000110100100111;
#1 $display("%b", po);
# 1  pi=207'b001010111110110111011110101010100101000010100010111010110111101101000010000100111011010010000110100101100010001011001011001000011010101111100000010101010110111000100101111111010011111101001000000011100110110;
#1 $display("%b", po);
# 1  pi=207'b110010000010100001101000011100001010111011111100011000111100100100111011000000111101110100110000100100010000100110100000110001010100111110011000010111011001110110001111000000011010011110101001110001110000100;
#1 $display("%b", po);
# 1  pi=207'b110110110100000110100011111001001110110000010010111000001100111011011000011010011010010111101001001111100111011101111100101111010010000001000001001010111000000100010111001011011111101110011010110010101010110;
#1 $display("%b", po);
# 1  pi=207'b001000101100001010100000000000000001000000011111010110000001000010110101111100010101100101111100001111010000001110111111100100000111110111011110010011110110011011001001110101111000000000110110111101001010111;
#1 $display("%b", po);
# 1  pi=207'b111011111010011010001000101110000010011011000001000000010000110001100011000000101010000100111101101011010000010000000100101110011000111001010001000010111111000000111000001000011000000000110101110100111001110;
#1 $display("%b", po);
# 1  pi=207'b011110110100010000001001001110100001100001010100101110110000001000101101000011101100110111110000000010100111101000111000000111000111111110110110001100110000110011111100000011011010001111000000101111000011010;
#1 $display("%b", po);
# 1  pi=207'b101100000010101101011000110000011110010001100110010101111111001111010100010110001110100100010100101110010000101101011101000011001010001001000110110101101010011011101001100100110101111001000110011001011110110;
#1 $display("%b", po);
# 1  pi=207'b010000110101011001101011010000001001100110011000001110110001001010100001110111101110111010001011011010101100001000010101001000111110101110110100000110111010001101011011101110110110001010100010100100010100000;
#1 $display("%b", po);
# 1  pi=207'b100111100010110011100010000001101110111000110011011101011100000110110101000000011111100010110100001010110100010000100110101010111000010000000010000111010010100111101100111100100101001101101100101000101100111;
#1 $display("%b", po);
# 1  pi=207'b111010010111111000011010111001101110010010110010110000110000000000100011000000101100001110100110101110000110101010111001101000110000101010010001011000011101110110110100110101001111001100111111100110110101101;
#1 $display("%b", po);
# 1  pi=207'b010101110010111101010001010011010011111111011000110010001100110101111001101011011110000101010110100111100101001101101111011100110010011111000111101010111001111101010000001111111111001100100000110101001111000;
#1 $display("%b", po);
# 1  pi=207'b011011011011101001011001111111110011011111101001011101001000110001011111011011100101110000110111001110101010000101100111010101011111100100010111100110111011010011101100101111001110011011001000000001110011011;
#1 $display("%b", po);
# 1  pi=207'b110001001101011010001101011100100111110011011010111110010001011011000010000111111101010101000111011100001110101101101101110101011011001010000011001001011011100010010000101111100111010110011011000010100100011;
#1 $display("%b", po);
# 1  pi=207'b011101000010110110000100110111110011110010001101110000100110110101010001010000000001010100010000111001011100101100110000110100100110010111011111100101110110101011011011010011101001001100101010100101101001100;
#1 $display("%b", po);
# 1  pi=207'b011010010111111000011101010110011000010110001110001010001101001000110010001111010111100110101001011101101000111011011000100001100001100111010110010010100100011000010110111110011000111110111011110000000011110;
#1 $display("%b", po);
# 1  pi=207'b111110101101010011111001000110101001000110111011110111000111001110011010110000000100000100111110011110010000011110011110010010100001000100000000111100110110110001010000111010000000101011011011111011110110101;
#1 $display("%b", po);
# 1  pi=207'b001100000101111111011000100110100111010010100100110000010101001011001010111110011100001100110100101010011101011011001101111100011010110000111000000000100110001100011010110000001000110000011011100101010000111;
#1 $display("%b", po);
# 1  pi=207'b110100001010101010101010111101010000101001100110100110010101110000001011011010110100111000111110010001101101010001010111110000011001101101100010000011011011011011111001011001100110001100010001101010111010001;
#1 $display("%b", po);
# 1  pi=207'b011001010100001001111001001101011011001101000101001101100110100101010110000101111110111100011110001011010011011110000000101110000010010000011011101010101001000100001010100001010111110000010101000000100110011;
#1 $display("%b", po);
# 1  pi=207'b000101101110000001110101010110000011000101111110101010100111000110101100000101010101111111001101100110101111000001001101010010011010000100000010011111001111110010001010101101111010110000000101000100101001011;
#1 $display("%b", po);
# 1  pi=207'b101000011011011011101011000111000001100110001111000111111011101001010001111010111100110110110011111010111001001000011100110100010000100010010001110101011101000011110000001111110100010100110010010111111010011;
#1 $display("%b", po);
# 1  pi=207'b110011010001111100011100011101110110000111001110111110010111111011110000101011000000111011110110110000001000110001101101001010100111100101000110011100100000000100000110000100010010111100010011001100100111001;
#1 $display("%b", po);
# 1  pi=207'b101111100000010001100001011011011110100100110000001110101101011111011100010110001010000111111100001110111101001001110001001110110101100100000101111010000100111100100001001101001010000101111000001100001010101;
#1 $display("%b", po);
# 1  pi=207'b100100101111100110010000010101110101101101101100100000110100000110001000011101010001110100001000100110001100001001100011011011111110011111000001110111110100000010010011001111101110011111010011000111110101111;
#1 $display("%b", po);
# 1  pi=207'b010100111111100011011011000101110101100000111001001000001011010010000101010110100011110110001000111100000111111110110010001000001100001010100010110111001111011110000011110111100000110100110101100111000010101;
#1 $display("%b", po);
# 1  pi=207'b001110101010100000100100111111111000000100100010110101101101111011000011011110001111110111000000011010011000100011110010000000101000101010101101001010101001110110001100110001000100001111100001001011110001100;
#1 $display("%b", po);
# 1  pi=207'b100000001111111111101010111010101111010011000100100110011110001001100010001101000101110100101011110000101100011100110111101000001111110101110010111011111000000110001101110101001101100011000010001101011001111;
#1 $display("%b", po);
# 1  pi=207'b101000101101100111000111011001111101011111111011011001111001010000011000000100100010110100100011111111001000100000101100101000011001000110110111011110000000101010001100011111111101000010011100111010101001011;
#1 $display("%b", po);
# 1  pi=207'b111001110101000000101100111101101011111011111101100000001011110111010011100100011100000010100010100101001110010010110011111001111101111010101101101101101101100111110111100000001111100011000011001111110110111;
#1 $display("%b", po);
# 1  pi=207'b010010101100110001001101000011100011111000110000000001101101111111001101101100011100100001000101000001011010010000101100101101100011010010010110101111100100011000100001000111101110000100111001011101111001100;
#1 $display("%b", po);
# 1  pi=207'b000010111010001011000010111100101111101011111001100001100101010000001101111100011011111101000100110100101110100110001010100100100111011001111111000001000111001000011001011100010100101010100000111010011101010;
#1 $display("%b", po);
# 1  pi=207'b111110110000101001001001011001111000101101011110100111111110110000010101000000110000001010011111010001011000011011110010101101101110111010111110111010001001000001000111001001100001110110111110001011101001111;
#1 $display("%b", po);
# 1  pi=207'b001110110011010110010110001011011110110100111001110101110101110010001101010100111100001001111011010101101001101111001110111011101101100001111110100000101110000010001111011100110101110100010011101100000011011;
#1 $display("%b", po);
# 1  pi=207'b010010010111000001010001110111100011111011001100011010110111110111001001000011010000011000011001000100000011110100110011011111011011001100101111011001100111000001101010100100011011000100111000101010100001110;
#1 $display("%b", po);
# 1  pi=207'b001101101110100101110010100010000001001110101000110101101001110000001110100001100100101001110001000000011111000101100000101011011111111101111101010111101010011100001110000101110010111101011101000011011101110;
#1 $display("%b", po);
# 1  pi=207'b101100111100000001001011101011000110010100110101010100100000010111001000111101011111011101110011011100010100011111101101111101110101110010101111011110101111110111000110001110111000110011011000000011000111101;
#1 $display("%b", po);
# 1  pi=207'b111010010101011000011001010101101111101000000111100100110010100001011001010000111100001110011100111100111110010010011110110101100001100011001000110100001011110010000101110100000010110000101100100101010010101;
#1 $display("%b", po);
# 1  pi=207'b100101001100100011110011011001000010000110111110000100111011011111001111011001111001100011011001011111100100101101100011110000000011001100101001011011111101110001101100001010101000011111110111010100101000000;
#1 $display("%b", po);
# 1  pi=207'b000101111111101010110000011001011000100010110011101001011110010111101011100010011110101010000001010010010101011001010011000101010001000101111000000010110001001000001110010000100001101101100111101100111101101;
#1 $display("%b", po);
# 1  pi=207'b100010010000100000101111110010010010011011101101100101000001111011001001111001011101011000011011111010111110000010001101011001110100010110111001100011000111000101001011010011001011111111001010110110100011011;
#1 $display("%b", po);
# 1  pi=207'b000101000001110110000111111001000111001101101101010100101001111001100001000100000000010001101011111101010001100110100101110010100011011100010000000100001110011001101011111110010000010111000110000111011111010;
#1 $display("%b", po);
# 1  pi=207'b010010110000100001110100100011000011100010101010010010111011110010100000100011110100100100110110011111010110101111010010110101101011000000010111101011010100100001001001010000001001010100100110111111011101111;
#1 $display("%b", po);
# 1  pi=207'b110110110110010100001111100011111101011101010101110000011000010011010000001001111000111111010110000010110000100000010010101010101110000010110001100001000101011111010110100100111101010010001101101001111000000;
#1 $display("%b", po);
# 1  pi=207'b011011000010000010100000110000101011010000000000011010001100010101010011101011100101101100000100111110001111001011100100111111111100101101010100000001100001100100110001100001000110110110011101110110010000101;
#1 $display("%b", po);
# 1  pi=207'b011111101000001101001111000001100110001011001101010010010010001010101111100001101001000111000000010100101000000001101001011111000110011111110110000000011011001111111101001010110110100010100100001000100001001;
#1 $display("%b", po);
# 1  pi=207'b001111100101011010101001101000011001101010101111110110100101111001111111100000010000101111111111011110000000100100110111100001011100010110100011100001000010000001110101101111111001101111011111101101010010001;
#1 $display("%b", po);
# 1  pi=207'b010111011100100000111100000010011010110000011101111001111010010001100110000000001100111110010010100111010100100101111101010101001000100001001000100001011011010101011001101010101010000111010111000001011101000;
#1 $display("%b", po);
# 1  pi=207'b101001111001011011101110000101011001101111010010000011000110110110001011110111101000111100101101001010101010110100011101111011111101100101001100100000110011110000000001000001011001100100000000001110110011001;
#1 $display("%b", po);
# 1  pi=207'b100110110100011000111111101111110100111001101111011111100100010010111110111000100011001001011100100001011101100101111010100100110110100001000011001111110001111000111010001110110011001100101010110000100101100;
#1 $display("%b", po);
# 1  pi=207'b101110101011001011011011101011101011111001000001101000100111010010010011101001000101011011111110100100010001011010111011010010010000110100100100011001010001111110101110010010000000000011010100101000110011000;
#1 $display("%b", po);
# 1  pi=207'b010100111011011001101110110000110001010010011010111010100000110110101011100010001011110011100011111111111111010101000111001001100011001111110000011100001011011111111111000011001000101000101101110110001110100;
#1 $display("%b", po);
# 1  pi=207'b111001001100001110100100011100101011010010100010000101001010011111110010101111001001011010010111101100101111001100101100100110011110001010110000110000101100011100111111111110011011011100110110001001000010010;
#1 $display("%b", po);
# 1  pi=207'b111110001110100101111000111011101001111000100111000100100011101000000111110101001110010101001110111111000101000001101110100111111101011001111100001000100011011001010101110111111111100111111010100111101000110;
#1 $display("%b", po);
# 1  pi=207'b001011101010110100000011010100011100110011111100000100111101110101000111111111110011010001110010110000101110010011010111110110110010000110000010010111000100100100000110010100100001011001011010110100010101010;
#1 $display("%b", po);
# 1  pi=207'b001100101001100010010011010101100001011111001111100100010001101111111101011010010000011010101010110010001101101100010001010000111100111001111111110100110001111000001010110000001101000000000001100110101000011;
#1 $display("%b", po);
# 1  pi=207'b010001001010110110101110100000101111010111000101000001100100001111100111011111100010000110101100111010000001110001011001010011000110000001010010010110011011000001111101011110110111101000001101001111001100111;
#1 $display("%b", po);
# 1  pi=207'b110100000000011100000001011110110100110011110010010010100101001111001010110001011011111001001101010100011010010110110011111010110000111010000011100111100001101000111100011000000100010000101001011100010011111;
#1 $display("%b", po);
# 1  pi=207'b011111001010001001111000001101011101100010101101100111110001101010001110110011011011100001010000011111001010101001000101110101110100010001001010101000001111100110101100011100001101111100010001010100001110001;
#1 $display("%b", po);
# 1  pi=207'b111010011001110000001001010010110001101001001010001101100110010001101010100011110011110011000110111010001011110101110001011011110100000111011011001001111101111001110000110000010110011100110001111110011011000;
#1 $display("%b", po);
# 1  pi=207'b111101000111101000000011001011011100100010010110001000111101010100111001110010000100111001100110100110111111100001001001001111001010001000011001000000001011010001000000010010000100101110000110110101111010111;
#1 $display("%b", po);
# 1  pi=207'b011110110010011010000111110000110101101001000101000000101010101101100111001011100111001011101000011011000000110000001011000010100110111000100100000011001001001110011001011110010001111111100110000001001100110;
#1 $display("%b", po);
# 1  pi=207'b000110101000011000101111101101010010000010100110000010010101010100000010101101010011011011110011000111001001011001100010010110101000100100101111010001011100000000101101000100101100110101010111111110000111011;
#1 $display("%b", po);
# 1  pi=207'b100111011011011111101111111111110010000100000001111001011110010011000001101111100100101010111101001110010001111111001111011111110001100100001110010000000011110010001100000001000100001100000011111111000011000;
#1 $display("%b", po);
# 1  pi=207'b000111001000110110010101010110011111000001001011110001110101010011101000000101111010000110000101101010000001011111011110011010011000111100010111010110011100001111101001011010100110111001100111000111010010010;
#1 $display("%b", po);
# 1  pi=207'b110001001101000001010001011001011011111000101111111101010000011000111011011010011001101000010101010010111010100111010111100011101000001001101000001111011111010000010010001011111111000010011101111011000111010;
#1 $display("%b", po);
# 1  pi=207'b000000111011000100011011000001101011001110000100011000010100001001000100100011110101100111101110110010001010110110011101010111010111101000001101001111011010111110010011111011001010101010110100010001111010101;
#1 $display("%b", po);
# 1  pi=207'b010010011101001000111100110110000110101000011000111110011010010110010010010001110110100000001001000011101111001110001111001000000111110000100010001110001010001111000101000010000101100001110010100010010111000;
#1 $display("%b", po);
# 1  pi=207'b000111010101101000111011110001001101000000010111000011011011100111111001110001010010100001001110111011111110001101011100110011110111100011010010001110100000101100101110000100100010001111000101101111000111000;
#1 $display("%b", po);
# 1  pi=207'b000110101001011101001001011011100001111110011010010011111111110010010001110100010100010010010100111000111000110011101111111001111101001100010100010101111111111111011110001001001010000000100111101101110000110;
#1 $display("%b", po);
# 1  pi=207'b001001100001011100100001000000101100111001001111001100000111011100101100010000011011011111111011111111101100001110010101000011001111101011001000010000110101010110100100001110000000100110011101011011111110101;
#1 $display("%b", po);
# 1  pi=207'b110100101011000111011100001100111001111000100001010110101000001101000011011101001001100011010100000111011100110100010010110101101001111100010110011001001010010110011001101101101011101111010011001001100101101;
#1 $display("%b", po);
# 1  pi=207'b101100100111011101010001001110000100001010001001010000000011111010011001011110010101011110010000011101101011001000000110110101111011100101101100101001111011110001111011011000001001011111010001001101011001011;
#1 $display("%b", po);
# 1  pi=207'b110100110000111100000011010001110010001111011101101100111000111110111001010010001111001111110000000001010000001111100100111111101111010000000010110001010010001011011100101011101111110101100100000011010101111;
#1 $display("%b", po);
# 1  pi=207'b110000111000000011111111011011010101111101000110001011101100101000001010111011010110001010100011001101010001110011111000101101011010001001101101111000110111011111010000101111010011101010110011100101111001100;
#1 $display("%b", po);
# 1  pi=207'b011101100101100000100110100100010110100110001010010000011011100111011010010000101101011101010011110001001110001111110011100111110101000011101101000110010110101010101111111110100110110111111110101111111011011;
#1 $display("%b", po);
# 1  pi=207'b011000000111001000101111001010010000010010100000011100010111101010110010010001100111100100110111100010001100010011111111011000110011100001000011001110111101111011111110001111100110000101100101001101111001111;
#1 $display("%b", po);
# 1  pi=207'b101011001010101010100100011100110000001010110100100101010111111010111011111110011010000111111001101011011101011000111001101111111111111011100111010101001110101001110011000111000101000011110111110111110100110;
#1 $display("%b", po);
# 1  pi=207'b101011111011001110111110101111100001111100010110100110001111110101100101101110101110001110010010011011000101011010100011100011010000011010111000101010010010011100011101110110011010100011010011110001111110111;
#1 $display("%b", po);
# 1  pi=207'b010100100000100001111110110111101001111000111000111110010110011001111101011011100011100110100111010100101010001111011111100101010100000000000001000111000011000111001110110110011111001001000001100010010100010;
#1 $display("%b", po);
# 1  pi=207'b010001000010111111101111100011111111001110011111100000110101001110100110010101010111111101010111011111010010001011101100111100000111001000101111010000000111111100101000100110011110111111011011101101111000100;
#1 $display("%b", po);
# 1  pi=207'b111111100000101001111000110110010001100111101011001001110001011100100101001111100101111110110100110001101110000101011111011001111110001110010111000010110000100010001010100001100100000011011100101000100010000;
#1 $display("%b", po);
# 1  pi=207'b110101011010010010111101101001000100110000000100110110001010010100100011110110011011100000101101000101111111100000100001010110100100000100011110111100100110101101010111110010001001010111111010010001111101110;
#1 $display("%b", po);
# 1  pi=207'b000111000111000101011111111100011111111000101101011110101101100011001111100011100110110000110001001000001100011011001001111010100100000110101010011010001101011001111000011000001110101101001100001010100100010;
#1 $display("%b", po);
# 1  pi=207'b111010001100000010100001101100101111101111101100110001010101101101010111000010110000011100001100110000100100100011111101010011000000100000110011001000001101011101001100011010100101010100011110010000100000110;
#1 $display("%b", po);
# 1  pi=207'b000001101111111110101111000111001011111001011001100000100011111101100000101111011110100110111111001001110100110011101111011011010110100110111011010010011011000111100010010111110101100101011110101101000100111;
#1 $display("%b", po);
# 1  pi=207'b100100010101101110111010110000000100100111101000110011010010101000011001000100010001101111000010011011000111111111111110000101111110000001010010011011110110100110100010100011101000000101010000000100101001011;
#1 $display("%b", po);
# 1  pi=207'b011001100111000011011001011111000100110101101011010010011011110101110000100101010110110111010010110101001010101011101001101011011100001111001000000011001010000101110000001001010001000001101111001011100111100;
#1 $display("%b", po);
# 1  pi=207'b100100011101000001010011111100011011001001011010110111111101101110000111001110101100001110000001110100010111011000100100101100100110000101111110010000111000110001000000110101101110001100010000100111010101010;
#1 $display("%b", po);
# 1  pi=207'b000010110010111000110101000111110111011111110000100100011111101100100011111110010100111101111101011000001110011110110010011011011110001010101010011111110001111001011011111011000110101000010011000001111101111;
#1 $display("%b", po);
# 1  pi=207'b000001000001001100101011101110001000001010011001110110110001100110011100010111101110000011010001001111000100101111110001010100110100000010110101101011110101000011010110101001000110110010011100100111011100010;
#1 $display("%b", po);
# 1  pi=207'b011000001011000001001000001000010111001101110110110111111100111101110110111000110100011010111100110011001000010000011111110100001000101101110001101010110000111101000010000101100110001011000101110011101111000;
#1 $display("%b", po);
# 1  pi=207'b101111110110000110110010000110111100010110011010001100010110010100101101011001000101101000011101111110010000010101011010010100001001110111010001110010110100001101000100001011001001101010011100111111001001010;
#1 $display("%b", po);
# 1  pi=207'b000101011011000111100100111011111101100110001000001010001011011100111100111100100011010101100010110001011000001111100100100001100001010111011010101110100101110000110010001110011101111011010110001010101111011;
#1 $display("%b", po);
# 1  pi=207'b111111000110011111111001001111000000001110000001010100010101001001000000010011001001110011011000101000101000110111010101101011110000011011010101110010000000110110001111110010111110010011010000110000111110001;
#1 $display("%b", po);
# 1  pi=207'b111010110001010110010101111011110110001010110011101010010111001100101111011100000001101011110110011110101100101011000001010110111010000010110110000111110110010000110101010101100001011100000011001000110010000;
#1 $display("%b", po);
# 1  pi=207'b001000011111101011101000011011011110110000000011011100111001100010110000000110011100000110001101110000101010101100001001000100101001101110000000100111001001111000000001001100111011111010000100000010100000111;
#1 $display("%b", po);
# 1  pi=207'b001100100010101011001011001100101111011001100011010100100011001100001111010111010011001101000000001010100110010111111001100001001101011110000011011101100101101111110000011000011111001000100000010000111001011;
#1 $display("%b", po);
# 1  pi=207'b110111000101000101000001111001101111111101101101001101011010000010110011001011101001001011110000100000011000101010010101101101011110111100000000011001010011010011011000100101011100001100011101101100000111101;
#1 $display("%b", po);
# 1  pi=207'b010011010101101110100100111010110110101111101010010110010010001000010001001101001010110101001101010101001110111010101010001011011000011101110000010001110110111101110100010101101000110010000101101101010101111;
#1 $display("%b", po);
# 1  pi=207'b000000100001110110110011111011001001110001101100100000010101010110010000000100111001010010100110010101001110111110101111110011000001101110111110000110101101111111010010001001010111010111110111010101110011110;
#1 $display("%b", po);
# 1  pi=207'b000010101100111101010101001011000111111010011010010101111111001011010010010010101111011110011000010000000011001111100011000101110010011100000000001010011101001101000000010101010000110001010110000000000000100;
#1 $display("%b", po);
# 1  pi=207'b010010011001110010100001110110101111000110100100010110001001001100100111110001101110011101111001000101111000000100001100111100010011011000110000110111101011000111001001010100100111001101000010101011110111110;
#1 $display("%b", po);
# 1  pi=207'b001011011001110100011000011000110011100010000001111101111000001111001010010000100011000001001010111011001000111100011010101111011110100101101010010100001101111111111110101100111010111000000011011011110011111;
#1 $display("%b", po);
# 1  pi=207'b111000000011101000000011101001001111011100010010011111001111010011110000111000011101011111100111000101000101101000001111010111011111111101111100000011101001000101110001100100110110011101110111011110000110101;
#1 $display("%b", po);
# 1  pi=207'b001001001010010011110111000110000101010101101001010001001001100100101101100010010000010110111100011011111011000001111010000111011001001100010100100111011100001100011101011111111011001111010110000101011011110;
#1 $display("%b", po);
# 1  pi=207'b110111100101001111101000111110110101011010001110010100001101010001000001101101010001101111010101110100001010010110011111011001010100001011111001101011000111100110110011110100111000101100010101111010100110011;
#1 $display("%b", po);
# 1  pi=207'b001010010000101111000101111110000101010110000001100100010110000100111101101000110100110100101110011010110000101100110100101111110010100101110000011010111110011000111011010111110001110010110100101110110001010;
#1 $display("%b", po);
# 1  pi=207'b011000100111001001001100000011100001001010110101101001001110010101111111101000111100110111101001101100011010010110111100001010011011110110101001101000001111100111111110010001011100001010011101111011011111000;
#1 $display("%b", po);
# 1  pi=207'b110101100001111100101111110000111110010011100000101000110101011000100100001110101000010100000001111110000001010111000111111000010010001010011010100001011011100011111001001011011101011111010101010100000011001;
#1 $display("%b", po);
# 1  pi=207'b010000010011000110000111001010101110100010010011111101000010111010100000001110100001100111000111111100000011111111100100110011101001010001100000100100101111000110001011011100111110111111111110001110101110111;
#1 $display("%b", po);
# 1  pi=207'b100101110111101000001101001111000000001001101111000001111000010010100000011001110110100101000101001001001111001000101111101000010010011110111110011001101001000110000010111000111011101011010000010001100000010;
#1 $display("%b", po);
# 1  pi=207'b001000100111100110010100010110101001110101101011110111001101010101011101111101110101100110000001111111111000101001000010011010101001001000111110010101100010100101110100010001001111010100001011101001000100000;
#1 $display("%b", po);
# 1  pi=207'b101010100111101101110111011011111101111001000000000010001110111111001011111101000111011111001001001110110011010101101111101100000110010101001001000000010001110101101010011000101001111100111011101111101111110;
#1 $display("%b", po);
# 1  pi=207'b101101011010111101101111001011001111101101000001100000011110010100100000100111010001001110100110110011000111001010000110100010011010101111100101010111100011011100000100000000000011000110110101110010000011100;
#1 $display("%b", po);
# 1  pi=207'b011101011001000101110000000001011001110100011010101100110100101011001011010111001101110001111011011001110010010001011011100100000000111000110111000001000101100101000010001001110111000001000110110010001110001;
#1 $display("%b", po);
# 1  pi=207'b110111100010101111100101111010101000101001100000100011000100001011001010000110000111100101011000110010010001000010011111100000111111110001100110101110100000010000011100011111110010011100011000100111001110001;
#1 $display("%b", po);
# 1  pi=207'b111000101010110111100101011111001010010001110110111100100001010101010100100000010111111100000011101000010000011010101100110011100110110110000110010000001011011010101010010010001010001000101011001110010010110;
#1 $display("%b", po);
# 1  pi=207'b101111111110101000101000101011101110000010011101111101111110100001011111000010001100010001011011000100011011111000010010001000001011110101011101100011101000000011110101001110010010110001001011110111001101001;
#1 $display("%b", po);
# 1  pi=207'b011100110111011011010000000010111101100010010110010100001100111100101100110000110111010010000101001100100000111100101111100110100011100001011110001001101001100110100001001100010100011100100100101001111001001;
#1 $display("%b", po);
# 1  pi=207'b100111111001010100011110001001110001011011000010001110111010010000010011010100110000010001111101110101100111001100110001011011010001100001001011101010001000010101011111001111101101111101011110110001010100110;
#1 $display("%b", po);
# 1  pi=207'b111110110010110111011110010001001010101111101101110001000101100010110000010100100101011111100101100000001110001001100010101111011010100001010010101001101010110101011001100111010010011100001100001111010010001;
#1 $display("%b", po);
# 1  pi=207'b010100100001000111000010000101011011101100000101011101110111010100111011010101011101011111111101010110111001111010001101111000000110111100000010001111110111000110000000000100110000110111001110100111100110101;
#1 $display("%b", po);
# 1  pi=207'b101000010111101000010011010110011110001100111111111110111000000111101010000110101001011011100110100000011111101111001100011010001100100010000111110101000010001100111100101000111111111111111101001100100111101;
#1 $display("%b", po);
# 1  pi=207'b011001101100110111100100101110000111011110000000001001001111001100111110000011001100010111110011001111111100000010101011011100011100100000100111101000011111100011010010010010110001110011010011111000011101000;
#1 $display("%b", po);
# 1  pi=207'b010000110010000011011010001100110010011110010000001011111100000101100010000000101001011110100011001010000001010010000001101011000001110000011010001101001001101001010000111001001000010010001011100111001000111;
#1 $display("%b", po);
# 1  pi=207'b100101100100100111000111110110110010010101100111000111010011011101001100001000010111011110101001110011101000110000100000000101001110111010111010101101110100110101110000011011111110111010001000010111001001001;
#1 $display("%b", po);
# 1  pi=207'b001100010101010001000111010100111001101110101111111000010001000110000111011111101100000010000101010111110000001001011001001011000111100100000000110010001100011100010010101101001100110001001000111100010110111;
#1 $display("%b", po);
# 1  pi=207'b101001000001100001001010111101011100100000101111001001011110011011010111000100100101101110100010110101001110100100011111101010111110100110011100101100010111100110001111110000010001100001000111000100100101110;
#1 $display("%b", po);
# 1  pi=207'b011101010011111010100111001111110000001101011011100010100011001111101110101011001100001111000011010101100101110000101001000010011101000011000010101100000000010101011000010010101001101111100101111001110110111;
#1 $display("%b", po);
# 1  pi=207'b011011010110101010111101000011010100001001100101100010101011110010110001110101110101111111010101010110011011111001100111001001000100011010110101000000111111000110010100110011011010110011101001110000111100010;
#1 $display("%b", po);
# 1  pi=207'b100010111100010011100001111011010010000000110011101101111001010100011100101111011101010000010110000100001110111000110000111101011111111011101110101010010001110001001100100000001110111011110010001101001001010;
#1 $display("%b", po);
# 1  pi=207'b011101010101001100111000110011010111001001111111000000101100101111010010000001100000000011010000100001110011011100111011111101011001001011000111001010110011010101001000011001000011100111010010101011000110100;
#1 $display("%b", po);
# 1  pi=207'b001100000111011100100000000011100011011011101001111101101000001110000001000101100010110010100100100010010010010111001000000011010010111000111100011110100001001000110101001111011011010011110110110001000111000;
#1 $display("%b", po);
# 1  pi=207'b001011011011000001001000110000011011000111000100100011001100000100111010010100101110111010010100010001010010101011010110010111010000011101011100101111111110010011000110100101101011010100010000111001110101111;
#1 $display("%b", po);
# 1  pi=207'b100001100001111011110110010110111100110100011110100000010110111101000011111011110101011010001010011111111111101000001111010111001001100001111011000011000100110111100110110001101011100101010111001111111010011;
#1 $display("%b", po);
# 1  pi=207'b001101101101101001100010011011101111000010000000010010101001010011100111100000011011110110110111011100100101011100110110010101001001100001111100111111011011100100111110110011000111000110010010000000010001000;
#1 $display("%b", po);
# 1  pi=207'b001000010001100010000110101100000001100111100011011101001000000111001100011110101011110111111001001000010101001011101000001110100000101110110011000101000000100000100111000111111111011111101011010000010001100;
#1 $display("%b", po);
# 1  pi=207'b000001100010010111000110000101000100111111110110010001100111010101001100011111110110010111000110100011000100101010000010111011110010101010010111000010100111110000110110011110011100000110001010101100110100111;
#1 $display("%b", po);
# 1  pi=207'b000001111100001000001111000101010011001111010111001000101111010100101101110011111000111011010011010100100101001001101011001111001101000111011010001011010010010100101111000111010010010111100101111011111000101;
#1 $display("%b", po);
# 1  pi=207'b010001110110110101101100100100001111000000100001010111000001100100110011001100100011110101111100100001100011010011000000100011111100000100101110101010011000100100000100110000111101000001111100010011100000110;
#1 $display("%b", po);
# 1  pi=207'b111000010111100111011001101010110011011010001010011011111110000101110010101101011010011110001111101000100000000111000110100110011001000111100110110010101110001011100001100101101110110000010111111100010000010;
#1 $display("%b", po);
# 1  pi=207'b010010011010001110110010000001110001001111010110010110111011110100001111000111001000000011101000000110110000001110010001101100100010110111111100110110010000100000010101100110101111011100000101010101101101101;
#1 $display("%b", po);
# 1  pi=207'b011010111111010000000111111100011101101111000001111000000111110101111011010100011111010110111111101101101010101100000101011011101011010110100011000100110010101001001110111101011110001001011101001110010001100;
#1 $display("%b", po);
# 1  pi=207'b111101010000001011101011111101101000100000000001000111100010001010011100110101010001101111111010101110111011001000101000110100010011001010111110110111110110111000001111001100010100000010000010011010100000110;
#1 $display("%b", po);
# 1  pi=207'b000010110000000101100000000000110011100100100001000011010111011011111110011001000000010011111010110111010100111010111000100001010000001001111001000001111111001010111000110101001101001010100010111000100010101;
#1 $display("%b", po);
# 1  pi=207'b000000100101000100010000001100111110010101110110001111011111101010011110000110001011100101000111010001010011000001101110110001000000101111011001010111110001100110000010101010001001111001101100010100011101110;
#1 $display("%b", po);
# 1  pi=207'b110111010110101010001101101011001000100110011101001110010001000110100101101010000101000100010011011111101110001110001011001111100101111001101011000000011101100001010111111100011010000100101110000001111000010;
#1 $display("%b", po);
# 1  pi=207'b101111011001000011000110011000101001101001000000111100111000011010001011010010111100011011001111011010010111110010101011100100111101001101000111100111001111000000101010111011001100101001111110110001111101010;
#1 $display("%b", po);
# 1  pi=207'b011001100001111000110001110000101001100110110011111000001100101011100010000000001110011010101110101101011110111110101111000111010010000001001011000011101101110110010010011000110111101010111001000100100010010;
#1 $display("%b", po);
# 1  pi=207'b001001111100010001111100010010011100100001011100111001110101111110110100100001001001011010110110011100101111110100100111000101010101110000100010011110011001110101110110101000000000111011001100011001100101001;
#1 $display("%b", po);
# 1  pi=207'b011111011111001001001000110110111100101001110111000010110110010101111000110000000011101011010100001101100110010110100001001000100101010111101111000110101101010010011110110001111111101100111100001100110100000;
#1 $display("%b", po);
# 1  pi=207'b101110101010000010001100010101110001010001101010100011101100111110110010000011000011010101000110010101000101111100011110001011011011100011011100110011010101010100111111001000101110011111011000001001101011101;
#1 $display("%b", po);
# 1  pi=207'b110001010000010000010100110100110101011011000011101001000010011101001101001000100101010010000010011010001110001000111111001000100010101100101110100101001001111110011001000011000101001001010011001011010111110;
#1 $display("%b", po);
# 1  pi=207'b110000110000011111001011110110111110001011010011001010100100000010011011110000101110001100011100000000010001010000111010110010010110100000111101111101110110001010111110010110000101101000010011110110110001001;
#1 $display("%b", po);
# 1  pi=207'b001001010011110000010110000110110011000011000110001000110011110001100100100101111001101110010011111011001111001110011001101101010100011001111011110001000010010111110001011010110010000111111001110000100001111;
#1 $display("%b", po);
# 1  pi=207'b101111001001100001011110010100011000110010011011000001000111010110101001101100000101111010001110111001110011111001101110000000100100110100011100101010111101011000010011111101011111000110110110101010100010010;
#1 $display("%b", po);
# 1  pi=207'b101000010011011011000011110011010100010001100011100111101010101100011000010100111001010001001101010001111101001001110100101100100000011101110110010100101111101101010010000011101101001001110001010100001100011;
#1 $display("%b", po);
# 1  pi=207'b101001000000001111000000101001101010000000110101001101101111010101111000001111110111010010101010110001111101000000001110111000100010000100000110111000010111101101000011000111010001101001111110011000000111101;
#1 $display("%b", po);
# 1  pi=207'b111011011001100111111110001101111111110011000000111010111010000100001011011111100001101100011000001110010111000011001000000100111110000000011011100010111000011101000110010010001110110101001001100110101000010;
#1 $display("%b", po);
# 1  pi=207'b000000100100010100010001110001101011101100011011011101111101100000100101000110001101011010101001010001011101111111100000011110010011111100011101111101101001111101010010110001010000110110111010010110011011111;
#1 $display("%b", po);
# 1  pi=207'b010111011000111001010010011110010100110101111101011110101000110110100101100100001111110000110000001111101111010010111011100000010000101011101100110000001100001010010100110111111011100000101101010011001011011;
#1 $display("%b", po);
# 1  pi=207'b110011011101110001101110111101111010100011001100111001010110101000001111100111001010110001111001010000101111001100110010101000110111010011011001000101101101010111100101111001011001000010101110011101101011110;
#1 $display("%b", po);
# 1  pi=207'b110001110000010010101111110110001000011100001000101100100011110010001010111111100010111101110100001111001011101111111100011000101010110111011010001000101111010011010100010111100011001001010111001010101100001;
#1 $display("%b", po);
# 1  pi=207'b110001100010111101000100111011110010011100010100110111110000011001111011110000001101000111101111100110001000000111001001111111111000101110101111000000001111101000101110011101111101010001010000111101000011000;
#1 $display("%b", po);
# 1  pi=207'b010100110011011011111100011011010110010010010000100101111110001101000000001101011001110001100101111100110111101110111010010111100011010010000010101001110001000000110111111010110001100010110001101011000110100;
#1 $display("%b", po);
# 1  pi=207'b000011001010111101111001100110001110000111111110000100110100101011011100111111111011001011101100000010000101110011110011111111110010010111001111110010100100010111001101101111110010100110001101100100110100110;
#1 $display("%b", po);
# 1  pi=207'b100111010000100100011011001011001101100101110111101100011001000110001111001101000010100100010001001011100011001111010010110010101111110100100000001100100110111001010111011111011110111100000111111110000100111;
#1 $display("%b", po);
# 1  pi=207'b000101110101001101000010001101101011110001000111110001001100101011011111110100010011101010001010000010111001100011000000000111000100111011001101101011100100001100000000110010001110111011000001100111101100111;
#1 $display("%b", po);
# 1  pi=207'b101111111010110001001010101110101000000101110001101001011100100001101110000111110100001000100111100010010100000101110100001011110101111101110011001011110010100001011011011000001101111111011101100101111010010;
#1 $display("%b", po);
# 1  pi=207'b111111101111111010010011000101011001101000001011001101011001001101101001101000101101010000000011100100000101101100001110000010110101000011101011000011000110001110000110010000111000110011100110000001001101101;
#1 $display("%b", po);
# 1  pi=207'b110001100001001010001110011111110110101000101111011100111111001011110001110111010010111110011010000100000010110100011101101110110001101101111001000100111010011001000000001001110011110100010000101110100011000;
#1 $display("%b", po);
# 1  pi=207'b110111001010010001001000101010010100101001011011101011100101000000011111101010000100101101111001010011001011011100100101010001111000100000101110010110001001111100011000110001001011101000100001100110100001101;
#1 $display("%b", po);
# 1  pi=207'b000100110011100110111101101000111010000011011101101111111010000000000001011100001110110111001101100100101010001101111010010100010011100100011011101111000011011010000011110100110101101111010111011011101101001;
#1 $display("%b", po);
# 1  pi=207'b011110001110000101111101111000100110110001010010100001111110110101111100100111110011000110110010001110011011010010110010110110010111011010000110111010100010001001001100100001000111101011100100000000101101101;
#1 $display("%b", po);
# 1  pi=207'b010001111110110110110000010110001101010101010111001111110011111011101101010001101101001111011000110101100111101101110101110000011111000101001000001001010101100100111011000101110011110101011101010011101010001;
#1 $display("%b", po);
# 1  pi=207'b010001100111011111010011100011010011010000010100110011010101111100110101001100100010000010000101100001010001010001001110010010100011101111011000111101101100100111010101010111110111111101001000111110000001101;
#1 $display("%b", po);
# 1  pi=207'b100101011001101010011101110111001000110010111011111010001011110000010101000110000100001010111110110111000111101101111001000011011001011111110010011111100101101011100111011100001110111111001110100000100011000;
#1 $display("%b", po);
# 1  pi=207'b000000010000001001111000011101101010111100011000010011000100001010110001101001101111101110100010011010011000000010000010111110111111010100101010101011101111111000011011010111000110111110010100000000010101111;
#1 $display("%b", po);
# 1  pi=207'b101110010100010011001000011010100000001110001000000010001011010101111111111101011000101100111010101101100110111100110111011111011100011011000111111111111000100011011111111000100010101110010011110001111110001;
#1 $display("%b", po);
# 1  pi=207'b011011101110101111111001111000010000011000101010110111010111101001111010001010010011110011000000100101110000010010010001101100111100000110001001100110110001001100111000101110100100010111100010110011000010101;
#1 $display("%b", po);
# 1  pi=207'b100010000111010101011011011011111000110001011101010111001100111011000100111101011010010001001110110100001000010001110010100011000100011001100110110000001100000111001001101101010001110010111000000100111000001;
#1 $display("%b", po);
# 1  pi=207'b110100010110100110010111001000000110011011111100110101010011100000101001110100010100000000111001101001001011110001110101111011101011111000101100011010010011111111101001001001011001011011000101000010000111000;
#1 $display("%b", po);
# 1  pi=207'b000101011011001010111100101000001111000011111001110001101000100100011011110101010010101100000001001011110011100001101011101101111011100011111000101001011000101101100011010101110011010101010001001011000100010;
#1 $display("%b", po);
# 1  pi=207'b100110000101010011000010101110010001100101011100010110001110100101111001000111100111000101101011101110000000110000100001101100001010110101011010101000001100001001010100011000100010100011100110010110000110010;
#1 $display("%b", po);
# 1  pi=207'b001110111100100100111010000111000100101000110000111100001011100110111011001111101101001101000000010101110001100000100010100100011100101110001111010110001011000001001001001010110010001001001110100110001010100;
#1 $display("%b", po);
# 1  pi=207'b010101100110011111000010001011001100000100111101111101101001100111100110001101110100001000111010110111011101110111100101011111001111110001100011011101011111101101011011010111100110000000010010001000010000010;
#1 $display("%b", po);
# 1  pi=207'b001001000001101110111010110000010010111100010000110110011111010100110001111110000110010010100010010010111000001001011010010100010000101110010101000001111001100010010110011100110001101011110011011100011001000;
#1 $display("%b", po);
# 1  pi=207'b101011010011110010110011110010011111100111110010100100110010110111111010010011000110010000011010001000001110111011100000110001001000000011101011011011111101011101000100011110001011110001000100010101010101010;
#1 $display("%b", po);
# 1  pi=207'b000110110111100100010111001110100010111011111011001000010000000001111110100001011001100111001111001011111101100001111001110111010111011001011001100000000100110110100010011010001001000001101111010011011000100;
#1 $display("%b", po);
# 1  pi=207'b110110000111100001101001010000101000110010011111010110100000110101000110100100100100101000011111111111101110001110000010111010001000010000010001010011101010100000100101110011001100101001111001111010010011000;
#1 $display("%b", po);
# 1  pi=207'b111001100110111010011111010101111001101111000000000000010111001000011011110111111110101110001010101000110000001110001111001001110001001110101100000001111001101001100010101100000010010010010001011011100110100;
#1 $display("%b", po);
# 1  pi=207'b011100111011101000110100100101011101001011101100100100111010010011100101110110111010011000001001100110100000100101011010110001000100001010110101001100000011101101110001001100101110110011000001111110000110001;
#1 $display("%b", po);
# 1  pi=207'b001010011000100010011011110010000100011100101100001011111001110000000110111101010101101011111011111011111110111101101101000000000011110110111100100011001111101011110110000010001010010010101000001100101001101;
#1 $display("%b", po);
# 1  pi=207'b000010001110111011110111111110010111100010111010000101110010001101000011111100000110100000011010011100110001011010000010010010001101010100101110101100000011010100011111110010000110001101100110101001110110110;
#1 $display("%b", po);
# 1  pi=207'b011010001010001101100001110001010000000000000010000101101100001011001001010111011010001001011010110011011101110110010100100111101101001111010011101111100001100000111110100110110010100101000110111100011110101;
#1 $display("%b", po);
# 1  pi=207'b101001010111010111101101010011001110011101001001001011011110100011001111101101110001011000111011000110001001001010110010101100000100111000110000100001011010101101101101010000110010111101001000111000011001101;
#1 $display("%b", po);
# 1  pi=207'b110100110101111000100011011101110101000111010101101000111101101110000101011011000001001111111011001111001010011000011100010000110110100111111010001100110110101000001001001000101110111011011000010011010010011;
#1 $display("%b", po);
# 1  pi=207'b110101001110110100011101010010111101111100111010111011011000101111101100101000000111000111111001001110100010100101000101110010011010011111100000110110010101011000101001001100100001000111111110100001101110011;
#1 $display("%b", po);
# 1  pi=207'b101100110110001100111101110001001001110111101000001100101100010111001011101110111011010100110001110011111011000111111010011010011001100101110000110100001101010111010101100011101100000010000001110001010101100;
#1 $display("%b", po);
# 1  pi=207'b010001101111001000010110110111000011100011101110111000010101100101010111010001011110100000011000001111111111000000001000000000011001000100010101001110000110110111011011100011110001000010110011110001000110111;
#1 $display("%b", po);
# 1  pi=207'b010011001101011000111010000000101010110011010101011101000101101101000111101111011100100110100010100110001101001011110011011111010010101010111110000111111001111000111011101010011001111010000010110001001111110;
#1 $display("%b", po);
# 1  pi=207'b111101011010110011001000100101111100000100111001111100010011001011110001001101110100010101010101100110110000111100110010100111010011011000100101110101010000111000110110001110000111011101100110011111111010100;
#1 $display("%b", po);
# 1  pi=207'b111100101001100100011101101111111011001110010000001000011101110101010101111010111001010110100011100010000100010110100111110001111101111001011000011000011100001100010011111111101001111000110011101000001010000;
#1 $display("%b", po);
# 1  pi=207'b100101011110111100110000001111110101101010101100001101010000010101110101010110100011001100000101111010011001010100001110000110111100110010011101110100000000011111001000110101001010011000010000010010101011000;
#1 $display("%b", po);
# 1  pi=207'b111100110000001010100010111100000001011011100000000001001110110001111111011100000000111011010111010010001000110011100100010011010111000110111101011110111011100010010011100000100101010011000101100001110110000;
#1 $display("%b", po);
# 1  pi=207'b001111110001000110101001011100101110010111110101101101100100001000100001111110011000101100011000110111001011001010001001111111011111111011010110001001111010011111100111100011101001110010111010001011011000000;
#1 $display("%b", po);
# 1  pi=207'b100101011110011101000111111100110001111010001010110101001000100000000111010000000011001111010000101110101110101101001001000011000010111011111110101000101100000000111010011111111100011110101000001000110001010;
#1 $display("%b", po);
# 1  pi=207'b110000110101110101010001011100100111101010001001100001101010101100100110000011101001001010101100110111110001111101011000001000101011100010001100110010011000001010001011101111101100010010111010100110101110101;
#1 $display("%b", po);
# 1  pi=207'b111101001001101011110100011101010100001000101111101100000010100110110000011011010011001011011000101101110011110001011010101001001011000100101001100000000100000111110001111100111010010100111100111011101010110;
#1 $display("%b", po);
# 1  pi=207'b000010011010011000010010000010110001001011101110101101101101011010011001001101100000100010111000001010111000110101100100111001100011010000000110001100101011101001000100010101111101000011100101001110111110010;
#1 $display("%b", po);
# 1  pi=207'b001101001000100010010100010100110001001100000000011011110000110100010001110010001000101011000101100010110101010111011100010100101110000111001000101001110100001100110011010101111111100011101001010110100000000;
#1 $display("%b", po);
# 1  pi=207'b111101111100110111001110010000010010111001110101111010011011100100010110100110000100001100100000111000110111001001001011011100000100000001101100000001000011100001000010100011111011010111100111010110110101101;
#1 $display("%b", po);
# 1  pi=207'b101010010000110101011000001000010101010000110001000010010010001111110010011101010111010010110110001111101110101000100011010010010101011100110011110010011100110011100101110111110000101101000101111110110100000;
#1 $display("%b", po);
# 1  pi=207'b100010110000011101111101000100000011010110010011101101011011100100100011101101000101011000001100111010011000000001010010101011011110101000011110000100101101100110010100000110010110111100100011110110001100011;
#1 $display("%b", po);
# 1  pi=207'b110111000000101110000001000110010001111100000111100011101000010101100110101101111100010100000010010001111100111001001110001100100101100011111001000101011011011001001001001100001011000110101111000101001001000;
#1 $display("%b", po);
# 1  pi=207'b010010001010011001100011011010001000111101000000001011110000101000111011001000101001111110110010011110000111111110110101011010010011100011000010000100110101110111100110100111100101101101000110110100100110010;
#1 $display("%b", po);
# 1  pi=207'b110000001101011100010010111010101011010101011011100010011111111100010101001110000000011110011011011000001101110110111011001011100010101110011011101111011111110010010100111000101100111010010101111001011000010;
#1 $display("%b", po);
# 1  pi=207'b100110000010110101100111000000010100110111001001100001010000110111101110110100010010011000011011010001111001001110000100110100101000111110000010001010100001100010010001110100110111101100010110101100000001111;
#1 $display("%b", po);
# 1  pi=207'b010001000100110000111100100101101101100111000111011111111011111000110010001101000110101011100010011000110110000000111101010011001011110001111110011000011100101111000010101111000001010110010101000101110100101;
#1 $display("%b", po);
# 1  pi=207'b011110100100011101000001001110100010101101001110111011011011101000001010011110011001111000110100101111110011001011111011100101100000110000001010101011010100101001110110101111100010000110001110111011011110110;
#1 $display("%b", po);
# 1  pi=207'b100000101010000111000100100011001100001010111101001000110111000110010001001000011000111100111000011011110010101110100111110101001100100000000010010111011101010111001100010011011011000011111010011011111100110;
#1 $display("%b", po);
# 1  pi=207'b000011110000010001111000010010101110111101000011111110111110001011101111010010011011100000010000100001101011100110111010000101000111011101011110001010110110101111010110011000111011101100111000110010001000100;
#1 $display("%b", po);
# 1  pi=207'b100001001100101110100001011000011001001000101010000110110110111110111110110101011001101100101100000010001101001101001100100001101001001000011011101001001110101111010000111001111000110001111010011101111001110;
#1 $display("%b", po);
# 1  pi=207'b110000000101010000111100001111101001100100110011010100110001000011110000110000010111101111011110000100011111001010101100000101010010010011001100011100111111001001000111000010100000101001010010000001100100010;
#1 $display("%b", po);
# 1  pi=207'b000111011000110111011100111011001111000110000101100100000011101101111000101001000011101000011000101101101111101110101110110110111100011000010110100011000011011001000100011110000010011111101110110001011011010;
#1 $display("%b", po);
# 1  pi=207'b101110101111010101101011010001111010110110000010100000110110100001000000100101110000111001110010100011100011001010100101110111100001001001011010000100111100100011001100110111101100110010001001100001010111011;
#1 $display("%b", po);
# 1  pi=207'b100100011101011100101101111010110010101001010110110101001010100111001001010010110011011001101011000111111000101000000001000101001010111111101011001001000001000011011000100100010001010011100011100001011110100;
#1 $display("%b", po);
# 1  pi=207'b101110100001011010011010011011010010010001010011000000100001110001001110001000011000001000011010011001111000000001111001111110100111001010111110111000010111100101011111000010011101110111000111110001110100110;
#1 $display("%b", po);
# 1  pi=207'b010111100101101110101011100110100110101101101111011000000011110000000001100011110110010001101011101111100001000101000000101000111000100101011010111011000111001101010101110000100100110001001001000001110111100;
#1 $display("%b", po);
# 1  pi=207'b100111010100110110111101110111000000100110110111000001111110010101111100100001110011011001010100111110000011011001110101110000110111001100110001011001001011111011011111000011011001101110000111000001100100000;
#1 $display("%b", po);
# 1  pi=207'b101101111111010010011011000111101011100000000010101111101110110000101011101100011000010001011010101001100000011111100100000010101001001010111010001010011111101010110110110101001100011000111111100110100001111;
#1 $display("%b", po);
# 1  pi=207'b011100011101010010011110010101000100100000101000000010010001000011101111011110100101100110001010010001101001011000110001101000001010001100001001011001110011000100010100100000010001001011011111000101011010110;
#1 $display("%b", po);
# 1  pi=207'b101111100101000000010000011101111001010101011001110011000001010110111111101110101000000101000111000100101000010001010000011010101001010001000111001100010100000110010011011010000100110101000101110010111101111;
#1 $display("%b", po);
# 1  pi=207'b011010011001101111111111001010111011001000000001011010001111110011110111110011001000010011111111110101001110110001000101000011101011011100110011000101010011111110111101111010011011000001111011111011001000100;
#1 $display("%b", po);
# 1  pi=207'b001001000010110100100000011111011110100111010100111100010110010001011000110000101101011000101100011110101110011010101011000100101011110101101010111000111011001111111101011101011111000000100001000000100010001;
#1 $display("%b", po);
# 1  pi=207'b110001011001001100000011000001001100000111100111111110110011011001010111001110100001101010011110010111001110100101110011111111000110010010111110011111111100101110010011110100101111011001100011110110000100000;
#1 $display("%b", po);
# 1  pi=207'b001010100001111100010100000111111011100100010010000111001111111010101101100001101100010110111101001100011010000011110001010011011101001100011000100001110010000001001101011111101110001011010101011101010100001;
#1 $display("%b", po);
# 1  pi=207'b101101100111000101111111000010110110101101001111010101101111101000101100111110101010101100001100001000100100110100101011010110010110000000000000100101000001000001100111010010010000011000001100000010010101001;
#1 $display("%b", po);
# 1  pi=207'b100011000100011000111010001110010101100011111110101100000110010101011110101111101110101100101100111000110000111110001010010001111011010110010100011111000010110100011011110001110011010110011101011000101000101;
#1 $display("%b", po);
# 1  pi=207'b110010001101001100111011010101110001011000110010000001111010111010111001101010100111001001110101010111100110001101101110001111101111010001010011000010011000100101111111001011001010111101001101111000110000010;
#1 $display("%b", po);
# 1  pi=207'b010010001101011100010111101011111000011100011001111111100000111011100111001000001001111101101100111010011001010110001100000101000000111111101110101110101000001111010111100010101101101000011011100111000010000;
#1 $display("%b", po);
# 1  pi=207'b100001001001100100000011000100100110111011000110101100000011000010001100000010001010100000001011100011100111111010000100001010100110111100110011011111111101010111111000010001101010110101111001000111001100110;
#1 $display("%b", po);
# 1  pi=207'b011010100110110011000111101010110000101010111111101010110101011101011001001101100000011100100000100000111011101101101000010011100001111001101011101100100001000011100010001101100011010111111000001010010111101;
#1 $display("%b", po);
# 1  pi=207'b000000000010111101011000100101111001110010001000110101000100100111001100010111000001000011111101001101110010000101101100111000010101100100101101100101000101001100011010111010011111001100000000001001111011001;
#1 $display("%b", po);
# 1  pi=207'b010011111011100100011110111101100001001101001100001011100011010011010001000111100110010111100000111010111010110110111101000100101110100100011011111101111110000001101010000010010001001010001000100010001100000;
#1 $display("%b", po);
# 1  pi=207'b100011101010101011010001011101010100000000010010000101100111000111001001101110101011111111100110011101000001010001001101010100000010100010001100001100110010110010100101111011011110001010010010001001111110101;
#1 $display("%b", po);
# 1  pi=207'b001101110111011001000010011011110100001100110111001100010101011111011011000110101010111111010101000011000110111011001100011000101101110100100011110100010110000001101100101100111100111010011110011000101011010;
#1 $display("%b", po);
# 1  pi=207'b011110100101001100101011001101001000111001001111110100001110011100111011111110101110011111111100111001001100010011000001010001010000111010011010110000000001100001101110100111110000100101110110110011011110011;
#1 $display("%b", po);
# 1  pi=207'b110000101001110110001011110101001101101100001100101111110000001111101111001110111001100101010110111100000111001010000100010111000110110100001011001001000110000110001000111110011111010101001100110101110010000;
#1 $display("%b", po);
# 1  pi=207'b101011010001011001010000000111101011000000001011011011001101000111010001000100011101010100011100111101111100111101010111011100100001110001110001010000100011111110000101000000001110100011000011110001110111111;
#1 $display("%b", po);
# 1  pi=207'b100101111010000001100011100000111100001010010000001111111110100011100001111100000000101011100000110111101001101110001010001001100110010100101100100101111010101111110000111111101001101010110111101111011001101;
#1 $display("%b", po);
# 1  pi=207'b011000011011011110111101110101101010000111110111010110100011101000010001010101011000010110101111001010010111100000101110111011100101100101011110011110111000101110110100001000011110001100100101110101010010111;
#1 $display("%b", po);
# 1  pi=207'b111111011000110110001001101111100010111110010000011110000010111101000101000111101101000001011010111110010101101010010100010000111111110000110001000000001001110101001110100001101111110100010001100110001110110;
#1 $display("%b", po);
# 1  pi=207'b011011101101011101100000010110110001010100111000111010100101011000110010011001010010000111101111011011001111100011110101001101011011001001010000101010101010001010100100001101110100001110100001110101111000101;
#1 $display("%b", po);
# 1  pi=207'b010101110110010100111000001101100010111110011001100110010100001100001101111010110101110010010001100000110111010001001001111110011111111101100110000100001011011101001111100110101001011110000101111010110000001;
#1 $display("%b", po);
# 1  pi=207'b110010101101110011010010110100101010100110011111000100000111111110101010111100110000010111110000010001000010001000000011110011001010111011111111000001011011001100100100011001000110011101110001001110110101010;
#1 $display("%b", po);
# 1  pi=207'b011001011001010110001001111100110001111100001001111111010111110101111001010101101011000010111110000010010101001110111001000111010000101010110000001100100000100001001110010101011101011010110001100000100100101;
#1 $display("%b", po);
# 1  pi=207'b111001110111000101000110101000111011110110100101010010110111001101011001100110011010100100100110110110110010110001011101100110110010100001001110100010010000000001001011010011100011110010100000110111110100110;
#1 $display("%b", po);
# 1  pi=207'b101111111010111101010100110111101010011010110000000111111010100101110100011011111010100101001011100010100110110101111101101011001110100111010110001010100100110001101101010000001101101000110001001111110010111;
#1 $display("%b", po);
# 1  pi=207'b111011001000001010110100101001100000010001110111111010001011000001110010100100110111110111110011100101111111110111100110000001010111001011001001100010110010011101000001111110010101100010001101010101000111101;
#1 $display("%b", po);
# 1  pi=207'b110000100011101110101000110000011100111011100100101101100011110100110111001110010010011101101111110101001101111000010111000110010110001101011111101010101111100101110101101101101000001110111101010000000110101;
#1 $display("%b", po);
# 1  pi=207'b000110111101110011101011100111111011101110100111111101110101011010000111101000100011011101000111000101110110011111101111110111111001111100001000111110100000110001101111100110110100110111101111100000110001100;
#1 $display("%b", po);
# 1  pi=207'b010100101111111101000000100010010000101110001111001000100111110101100001011010111000001011100110111110101101101000101111110110100010100100001101111110000101000101011101010111101110110110000110111001000000100;
#1 $display("%b", po);
# 1  pi=207'b001110011000110110011111011110110010101111000110111001101000110111010011110000110111111110011011001111100010100001100110100101110010100110011011110110101010111001001111000010111011000101011011010001001001111;
#1 $display("%b", po);
# 1  pi=207'b100010101011010000101110001010011010000111011001101010101001100100101001100000101100110000100001001110101010100111110111111010110100101011000101000010101100111000010001100110111110111011010010111001000010100;
#1 $display("%b", po);
# 1  pi=207'b100101000011110011110010000111000111000100101001011101110000101110001100011110011001100011100010001001110101011000001101010111010000101010011111101000001011110100000101110110000010100011111111000001010011111;
#1 $display("%b", po);
# 1  pi=207'b011101011000011111001110101111110010001100100100101101010001000011100101011110110010100010011101100011010000000010110101010000010001000101100000000000011110100111111101101011101000110101101010010000000010101;
#1 $display("%b", po);
# 1  pi=207'b011000000101111010101111111111010011011001011100001000111101101100010011001110010100111000100011011000110000011110000011110101111000010101100100010111011011100001111011111000110100101000010010010111111110000;
#1 $display("%b", po);
# 1  pi=207'b100100100001001111011110000100110011111111101110001001000100000110110010100001000010100101011000010100001101010000100001111110001110111001111100000111000101110010011001011110110010000111101001010010100001111;
#1 $display("%b", po);
# 1  pi=207'b011111111011010101100110101000110011011111111000010011101100100001101000001101000000101100111001110111110011010011111111110010010000101001101101010100001101010100111000010011010100001010001011111000000011011;
#1 $display("%b", po);
# 1  pi=207'b111001001110111001011101100111101110111101110010000100100000101001011100110000111001110011110010001011011111011010110010100101010111100000110111110110000111011010010011010110011001011001001010000101100010000;
#1 $display("%b", po);
# 1  pi=207'b001100011111000111000011111001100000001000010100010110001100011000000111000100110010010100000010111011101000100110100100110010001000100011101001000101010011111100101111100001100101111110100111011000101001011;
#1 $display("%b", po);
# 1  pi=207'b011101000000001010010110010011001001000001100110110000000110011000110001101101010101011111011100110001010100111110110111010111011110011001001001010110100011011010001011110010001110001001100010100011000100110;
#1 $display("%b", po);
# 1  pi=207'b000011100111111111000001010011011001111000100011101000110101010011111100101000010111111011100101010010000001010100100100101010100011000110000110100101111001011110110010111001011000010100101001010111111101000;
#1 $display("%b", po);
# 1  pi=207'b010101110110110001010110000111001000010011110110010011000110010001110110011000110111101100101101001100011001110001001111110010010010001110100110110010100011011011011010110101001011101101001101111000110001110;
#1 $display("%b", po);
# 1  pi=207'b001111001100110111101010100010001110011100110010011100100011111001000110101100001101001010110000100100110101111111101011001000110001010010100101101000011100101100101100000010001100000110111000001110000011001;
#1 $display("%b", po);
# 1  pi=207'b010010010101100000101100101100010000101101101110110001010010111001111001010001011010101101011110100100110111110010111011000011001010010011100011001110101110111111001110110110111110001001011110100011000001111;
#1 $display("%b", po);
# 1  pi=207'b110011100000000011111101010001111110101110100110011111110000101001100100001111101100011100000100111110100100000100101111000100101111011000000000011010000100011111011111011101111110011000000101000100011010111;
#1 $display("%b", po);
# 1  pi=207'b000111100000100101110000100000110001100100000000101111110111101111001001111010100011100000110101000110001011110001110110010010100011100010001000111111001101000011110010110000010001101011101101101010100110111;
#1 $display("%b", po);
# 1  pi=207'b110110001000001011000010000001111011101101011000100001100100000010001100101010111011011000000010010100110111111011110111111011000100010101010001011001111111100000000100001110110111110110000010110110000110001;
#1 $display("%b", po);
# 1  pi=207'b011100001101100110101101001001110100000011100110101001100001110100001100101101010110111000011101111000010100001110001000011110110110000000010010101110011010000111111101111000001001000011011111000110111110101;
#1 $display("%b", po);
# 1  pi=207'b101100001000100000101011111010010010100100100101101000010010100001100110110110111111101101011111000010011001001111010010110010010110101111110110001010000001001110001011010110000110011000111010010001010110011;
#1 $display("%b", po);
# 1  pi=207'b111001101010101110111101101000100100001110010111111110101011111100001010001101010010101110011010000000001001100110011111100101000101011110100010000000111010111111000100000100110101100110011101110101001001011;
#1 $display("%b", po);
# 1  pi=207'b001111110001100110110100101011110000111110011111011100110001000010100100010001111001100011001001101000001001100100010001001101000111000111111100111100101001010111010011010000010011001011000011111101001001001;
#1 $display("%b", po);
# 1  pi=207'b110001110100001001101001101100000000000011100100111101001101100001000100101011001011010001100001100001101111010100011000111011001100111010110001011110100110100111110110100011101101111101100011100100010100010;
#1 $display("%b", po);
# 1  pi=207'b000101111000101101001011111000001111111011011000001111010000100001110100111000011001011010011101010001010001101101101101101110001110101111101001110011001000001001110100111010011011010101101101100101101011100;
#1 $display("%b", po);
# 1  pi=207'b011011100100110000001001011100110101101101001010100001110010000001000110011011000101010101110001011011101000000001010011111111010010010101011110011111111001111010010000010010110100110010100101101100100101111;
#1 $display("%b", po);
# 1  pi=207'b010000101010010011101110111001111000111110100101000100000011010011100100001110000111010011010110110111100011100101011000000100110010000000110110101001001101011110101101110001100111011101110101000010001100000;
#1 $display("%b", po);
# 1  pi=207'b000100000100000100100110101001000000010100011001011001110001001011100000001011010011101000101001011111110011011110010101100011111010000011011100011101011010110000011110000101100001001010111000110101011101000;
#1 $display("%b", po);
# 1  pi=207'b011110111011101100010101010000000010011101001010001001101001111111001110111011100010111100001101000010111010011001100110010101011011101110001011110111101011011011001010100111000010110101111101010100111110001;
#1 $display("%b", po);
# 1  pi=207'b000110001100101001011001010000011110001010011000010011101011010101110000101101001110011101011111010011111111010011001111100110100111101000101000100000001110000110001010100011101100111010011111010111001000000;
#1 $display("%b", po);
# 1  pi=207'b010011111010110011110110011000100101000011110100110001000111000101010010110000011100110101100001111001111101001000110010001110111100101100001000011101010000101101010111110110101000010101111111100010101001011;
#1 $display("%b", po);
# 1  pi=207'b000100000011101110111101011011100010010011110011111000011011100000111000011110111010110100100110001001010000010000101001100000000101010011110001100011010100011111011000101110011100000010110000101011000110101;
#1 $display("%b", po);
# 1  pi=207'b000000110011011001110011010111101011100010011100101100111110111011100001001100110110111001111101100100100001111101111001010000011110100100101100111000010101000011111101100010110101001010111010011100000001110;
#1 $display("%b", po);
# 1  pi=207'b010010010001101000010111000010100010110001001000111100111001011100100010100100101110101010100000000101100110110101110000001010101110111100010110000101010000101010100110101000111111100000000111001010000100110;
#1 $display("%b", po);
# 1  pi=207'b100111010010000100111111011010011011100110100001110100100011010001110011111110110010010100101110011110011000111001000001111111111110111100001011101011101001001100000001000011110110100001100011000001110001110;
#1 $display("%b", po);
# 1  pi=207'b000100000011101111011101010010010100101110000111100110000100111011000110100001000001100001000010110110010001110100101010110011111101110000101110110100100001011010100001100111110010110111111110001100111000001;
#1 $display("%b", po);
# 1  pi=207'b110110100101110011011101111000111101110100111011100000011100001011000100010111101111010001000010010101100101110010010001100101100101010000011100101010101111110010011001101010000110001010010000011001000011010;
#1 $display("%b", po);
# 1  pi=207'b111000010000000100110111010010010101001111010011001010110110100000000110100101001001001100110010001101101101101010110010010001100010111101101000001011000011000100101100001000011001101001110101001001110111111;
#1 $display("%b", po);
# 1  pi=207'b011100010101010010000010111000110101010111001000000010000001010001110010000010010100001101101011111111110100100010100100000111000010011001100000011111000010010010100101110000001101110000011110100001100001010;
#1 $display("%b", po);
# 1  pi=207'b100010010011101010001010010001101101110011100101100110001000000100110000011100101011100000011000111110000011100000011001000111110100000100001001111100010010100010001010100111010001011001010101111000010010000;
#1 $display("%b", po);
# 1  pi=207'b011011000011010100111001010000101111111010110100010001101000010101010011110101011010001001000001000110101101000101101111000000010110100101111001110011100001110111011000110000001100001100010000010001010001101;
#1 $display("%b", po);
# 1  pi=207'b101111001011000001111101111000000010011111010100101101111010000000000011011110001101010111111011011001001101011110101001111000010010111000101100000111110010111000100110011111101111001100110110011011111101010;
#1 $display("%b", po);
# 1  pi=207'b111010111111010000001110010010110011011101011101011010100100000100011101111101100111101101011001100011000101000101101101010110000101011110111011001010010000111011110110110110010001010110100001101101110111110;
#1 $display("%b", po);
# 1  pi=207'b010001101010011000101100101001000111011010101100001000011111000111110101110111001001011101111010111100110110000100010100010000111000111000100001110000000001000010111110101001110001110011110111011011011010010;
#1 $display("%b", po);
# 1  pi=207'b110111100001011010110110100111010000010111000100011111011111001010110110100100010001011010000000111010101001010000001101011010000010100001100111010100100110110010011110010111101111110011100111010101110010010;
#1 $display("%b", po);
# 1  pi=207'b011110010111010101101100101101011001110101011110111000111010111010001010110011010001101110100101101100101001010111100011101010010100100100001000100110100110000110011100101101101011100011010101001101101010010;
#1 $display("%b", po);
# 1  pi=207'b011101110111010000011111110010001001111101000110010101001110000011010010110010110011111111001101100101010101100100010110010100011000001010111100000111011110111110100011110011111011110011110111101001001101100;
#1 $display("%b", po);
# 1  pi=207'b111110110001010100011001101100000101000101101001111100000001000100011001000101011100111001111010001001000100000010000111001111001010110101010011010101101100110101001101101101100010110001100011111101110111011;
#1 $display("%b", po);
# 1  pi=207'b011111110010110010110010011100101011001110111000010101110100100011101011000100001001110111010010001001110001110111001010010111000001010111010011011101000011001100110100111110000111110010111001111000100010011;
#1 $display("%b", po);
# 1  pi=207'b111100000101111100011001101011001100110001010000010000001111100000110101111111001010101110101010110111110000101000000111011111111100001000011100000101110001010111010100101110001110001011001011100011010111100;
#1 $display("%b", po);
# 1  pi=207'b000110010001011110111001100011001111001111100100000111100010001011010011100111100101110100001111010100000101101110101111101011000010001001011111010110000010101010000001000100010001111001001010100100101101101;
#1 $display("%b", po);
# 1  pi=207'b011001110011100001100010011111111000110010100001010110010001101010111100111101100001001111011000001110101101010100010110100011111110111001011111110010101001000000110101111100011101010010110111000000110111010;
#1 $display("%b", po);
# 1  pi=207'b100011111110011010100111101000100111111100110011101000110001110001000111101111110101111111001100000101101110101111010100100100101111001000100001000100011001110111110110100111101100111001000101010101011000011;
#1 $display("%b", po);
# 1  pi=207'b111100110001010110111010110001000110101001111001101110101000000111010100000111111011000101110011101000010100000000111000010011011110111001011011011111100000100111101100001000101100000011011000010111111010000;
#1 $display("%b", po);
# 1  pi=207'b110111101100010010010010010000000001111111001011101111000000000100111111000110110111110000100101001011001110010111100101111011110111010011010101110011111100011110101001111100101110111000111001101100010110100;
#1 $display("%b", po);
# 1  pi=207'b000110001001011000001110110110010111101101010110111101110011111000111011100111010010111100111101111100111110000111000001000111110011101101110011111001101101111101000011111111000100100111101111010010000011110;
#1 $display("%b", po);
# 1  pi=207'b001100011011011000001100000001101000111111100101001001011000110111011110101100010000110100000100111011001111001101010001001111000010000001000010100011100010000101000011001011100100110000000001100100101100001;
#1 $display("%b", po);
# 1  pi=207'b011010101011101101110110100111011010011010111011000011010100110111011101001110101010011001000000000101100000110101110111101110110110110001100010110110011000010110001110110001110001101010101001011010011111111;
#1 $display("%b", po);
# 1  pi=207'b001001100111001100000010001010001101110111110101000001110001001001010111000110010110100010011010001000011100101101010010000110001110000001101000010111110001100001001111100100011010011100010000101101000101010;
#1 $display("%b", po);
# 1  pi=207'b011111100011001111111011110100111111101101100011000000011011101010010111010110011101001111111101111010111111010100010111101100001111011110111111000100011001111110110001111111001110111110000111000110000000001;
#1 $display("%b", po);
# 1  pi=207'b101010000111001111110000000110101010101000110000111111000101000110001010010000111000011111000110100110101100000001011100010111100011111110101110110000011000100101110101011010011001100010001010011011100110110;
#1 $display("%b", po);
# 1  pi=207'b001110010101100101110101000110111101000011000101101001001011010000001010000110011010110001101111011001110100101000110110000111111110010100110110100000010110010101101101100110011000101000110001000111100001011;
#1 $display("%b", po);
# 1  pi=207'b011110010000000101110111011100100001101000001100011111001100010010000011101010101100010110110011110111010011110010110111011010110110101010111110111100110000110001001100110110111100000110110000111111111101010;
#1 $display("%b", po);
# 1  pi=207'b100000100110101101010101010001000111011011101001001000111011001100000001001011110100101111100111010001100101000111001101111111001010100111110111000000000110111011101111100011000001011010110110011110001100001;
#1 $display("%b", po);
# 1  pi=207'b011000011101001110001000100011101101001000000100010111000110110010111010010101000100101011011001110111001001010011001010011011001100001000000011100011011011001011101111101111000111101011100011011010011111101;
#1 $display("%b", po);
# 1  pi=207'b110000000001111001011100010010101000111001010100100101111011100100010010101010101100111101011100110011101111101101100100111111001110101101000011010010100001111001100001101011110101001110011101011101111010110;
#1 $display("%b", po);
# 1  pi=207'b010010000100111101010010001010100000100111101010011001010110110010001100011000011100001010011110011111000111100110111100000111100000010001001100100100110100101110101110111011011011111011100000101111101101000;
#1 $display("%b", po);
# 1  pi=207'b011101000110001010001111101001001100011001000000111101101101010000000100011101001101110010101111010100100100101001101011111110110111011001000101010001000011111001111111110100111111010100010001000101001000001;
#1 $display("%b", po);
# 1  pi=207'b001101111100000001010110001110011001000110100000001010100011111001011111000110111010100101101100110100000110011001001110100000100010100111010010110010011101010100000101110011111101110001100110011101100110000;
#1 $display("%b", po);
# 1  pi=207'b010001010000011001010110001111001010000100111000110010000110100100111011011000100100001010111100000101100001000001111000010001001100010011111010101111000010101100011100100101100000110001011110111111010010110;
#1 $display("%b", po);
# 1  pi=207'b111101010110011111100110101110010000111011101000010000011110100110100011001111000100101100011101111101001110101011011101110010010111000010011010000000100000011000000101110101000011000111001111000011010110011;
#1 $display("%b", po);
# 1  pi=207'b000100111000110011111010101100111111011101101100101111101110010101111000000110100001001000100010111110110000010001010111000001111000111001011001001011000011100111110011111000011111111011001001010000010011000;
#1 $display("%b", po);
# 1  pi=207'b010000000100111011110000010110110011000101111000000101001000111010001111011111111000101101011110110011101010010100000110110100001011001011011000000000010010101110110010110110110110001000110110111101011111011;
#1 $display("%b", po);
# 1  pi=207'b001110001100100111111010001110010111011110010000010011111011111100010110110010010100100111100011010101101101111110010001010000101000100010111101001100000110101111001001010111111010111101001110101011101111010;
#1 $display("%b", po);
# 1  pi=207'b100011110010101011000011011011011100010101000001111001100011111011111100010110111100000011111011110111101101100111010000111111100010110100011110001111010000101001011100010001011100011101000101100110100000110;
#1 $display("%b", po);
# 1  pi=207'b100110111011010001010001110010101100000111110000111011001111110100010101000110100011011000101001010101110010001110110010100001100010100000100011100101001000000010110011100111000000101001101001110001100111010;
#1 $display("%b", po);
# 1  pi=207'b000100100011111000100010010001100011101000011101010111100011001110100101111110101010011001100111100010000111001001110101011010000011001010111101101010010000000000000001010010111111010101000100011011011111010;
#1 $display("%b", po);
# 1  pi=207'b101100001000010001010011010100100101110011101010001111111110111001000100100011001010101100110011101111101110010111000101111110001011111010111101010000001100001011001010100010110010010010110111101010001011001;
#1 $display("%b", po);
# 1  pi=207'b000110011111100010100001000000011110100001101001000011100000010011000010001001010001000011011010100100111001001000100110001010101101000001101001001100011110011111110101111100100100010101110100110000010111000;
#1 $display("%b", po);
# 1  pi=207'b100101111001001001000110100000001011000010010100110011110000100101010100011001011000001001011111100011010010101100111001111010001000000101101101110011001010011101100101111000100001000000011000000011001011101;
#1 $display("%b", po);
# 1  pi=207'b011001001010010011111111000001001110100110101010101001101011110001101101110100010110101111101001100101100111010001111111001100010111111000010001011110001000010100001011011010101110100010011001101010010000110;
#1 $display("%b", po);
# 1  pi=207'b110100001111100110100000111111111001111011100001000001000110010010011010000010111110110011000010101101001011001110100000111011100010100110010110100010101011011110110000110110000001000011010010100110001101000;
#1 $display("%b", po);
# 1  pi=207'b000110111101110010001010100100111000100101010011111110110110110101010011110001100001111000011110101000000000101001110010111001010100111101001011000000011101110110111110101000001100011100101000011000110010111;
#1 $display("%b", po);
# 1  pi=207'b011000101111011011111110011010011111100101010011001011110011101001111010011011011000010010001100011110101111100101111110000010101001001110000000101100110011000100010111110101111010001101011100110011110101101;
#1 $display("%b", po);
# 1  pi=207'b011101000001001110000000100100100100000101001100101111111101110010101001011011001101010011101011001101010111010011110110001110101100100010001111111100001111101111110001110100000110100001010011111001011101110;
#1 $display("%b", po);
# 1  pi=207'b011100000010101100100101001110011111110111111000011110111010101000010110100101011101110000010101100101111110100010011011011100111110011011110001100100010001100111000011100101011000010101100100110010100101101;
#1 $display("%b", po);
# 1  pi=207'b001110010110101010101110000000101011001011010101111000101010101010011010100110010111010101100010011110110111100010100000110010001011011001010010011001111010001001000000011000000001101010011010100001011010000;
#1 $display("%b", po);
# 1  pi=207'b101001110110101000001000101000101010011011001001101100100000110110001001000111100000001011101111111010010100100000011001010011110000111100110000100011010011000011000111011111001111000001000111011110001110100;
#1 $display("%b", po);
# 1  pi=207'b001100000001100001001010000000001110000011001101110000010011011101010110000000100010111111011111101001111011000000110110001001100001100111111111101010100101001100010001100011100011010001110111010000100110011;
#1 $display("%b", po);
# 1  pi=207'b000111101000101010100001111010110110101011100011000001001011011101010010001000100001011001000111100010101000101101110111011001101011110111101001001001111001001011001100110011101100110010111111111111110101110;
#1 $display("%b", po);
# 1  pi=207'b000101001110101011100110100000110111100001110000111010010111111001010010100100100001111010100010000111110001101110001111000000100011100100010000000001001110110001101100001011010100100011111000000011000011111;
#1 $display("%b", po);
# 1  pi=207'b001000110001000100010000000011010000100000010101110101010111001010111011101110110100110110101100101101010000111110010100011111100101010111110111111011010100010100100100100101010110101111010100110000001011111;
#1 $display("%b", po);
# 1  pi=207'b100100000110110010101101010000101111000001011100110001101010100011001111001111100101000101101001110010101110000100111011110110001101110101100100001110110011000101101110100011011011001000001111110011101000000;
#1 $display("%b", po);
# 1  pi=207'b001111001001111000010101100110000001011011011010011111011000001101100100111111011101111010101101100010100111001001111010010000011001101110011000001010100110100011110100101000011100100001010011101011001100000;
#1 $display("%b", po);
# 1  pi=207'b000110101111000001010001011010110000100100001110110100001100110111010000011110111010010100101011111010010011011101100100011001011110111000011011100010001101010111001111011110011110011100101110100100000100010;
#1 $display("%b", po);
# 1  pi=207'b111010010011100111110010010011110100111010100110111100010111100100010100101001000110110010110111000010110011100110001001001101011000100010101111001010011100010011011100110000101001010001100111111010000101010;
#1 $display("%b", po);
# 1  pi=207'b101110011100100101010101100010110010111011001011111010110100011101001111100111010100100001100001111010110110111110011001000011011101001101101111001111111000010110111000010000001000000111000100000001111000111;
#1 $display("%b", po);
# 1  pi=207'b101110101000111110000111011110000110111001011001011011110010011111001001111100000011001001101111011001110011111111001100101110000000101000001111010110100001000000101110000011000111111111101100110000110110000;
#1 $display("%b", po);
# 1  pi=207'b110111010011110001011100110101001011010110100100000000100010010101110101110000110000000011000011010100111011000101001101000010011110010011001110011000011010111110101100110100110001000011010110101110110000010;
#1 $display("%b", po);
# 1  pi=207'b100011001011011010010001000100101010010101110000011010001111101000010010011000101010100000110000101001110101000101011000011111000011100111001101111011111011111000111000010000110110111110001001101111101100111;
#1 $display("%b", po);
# 1  pi=207'b110000111010001011100011101111010101101010110010011101000000101100100101111001110000111010110011001111100111010110000001010001100011011001000001001010001101100010010111100000111101100010000100100000010110100;
#1 $display("%b", po);
# 1  pi=207'b011101011010101101000111000110000100110001100010001000001111010001011110000111101111110100010001100101010010011001001001001110001010000001111101000110101111001000010011001000001101110100110100100110011111111;
#1 $display("%b", po);
# 1  pi=207'b011011100101101011100001111001111100100011010111101000101111001010011000111010111000010110111010000010101001000111111010111100110000110111011111001000101011111110011010111011000110111111010011110100101100100;
#1 $display("%b", po);
# 1  pi=207'b001100011110011010111011111100000110001111000000100001100101001010010001011111010110010010111100001000101000100101110111010110100101010001100001110111000111001010110100010000101110111111001111001010000100111;
#1 $display("%b", po);
# 1  pi=207'b001100110110101110010010010010101100011001010110000010010011001111110010100101011111000011111000000010110100011110000100001100110101111111011110101001100000111010000110101011001111000000101010010011100100100;
#1 $display("%b", po);
# 1  pi=207'b000011110000011111001001010001010011101101001101101110111110100111110101010111100010000110111111110101000001010010000111010110000100000110001110011111110101010000001001110011111001110111101010111101101001011;
#1 $display("%b", po);
# 1  pi=207'b011010111010111110110111111001111100101100101010011100011011000111011110110001101000011010000110101111001010000010001011101001101100010011011010010110001000101001100011110110110111110001011011111100000101111;
#1 $display("%b", po);
# 1  pi=207'b100011010011101010010110010110110111100101111110100111111111010100000111000011010011111110111010011101100010011000001001010011111100011110010111111010010100111101000000011110000000101100011100001001010011100;
#1 $display("%b", po);
# 1  pi=207'b100000000111000011010001011100001101010111011100000101001001010001001111011011110100111100100101010000110010010000011011010101111000001001111110110111110000110111110101010111001011111101011011111011110000010;
#1 $display("%b", po);
# 1  pi=207'b000010110111000000101111001011010101100010110101100110100110010011001001110010011101000110101110000101000011110110011001001000111000111110111111011110101101101111100000011110001010010000101011010010100000101;
#1 $display("%b", po);
# 1  pi=207'b001011010011110011001100000111011101100111100001010000000101001011100110011010111010100000011111011110100001111000101111111111111011111100000110011110100001010000101011001000001110011110111011011101001100111;
#1 $display("%b", po);
# 1  pi=207'b111100111001101110001011110110001110111011010110111111010001010101111110000011011010101100111000010001011001101000011010011001110011001110111001110011011110010010000001011011011001110110010011110110000111000;
#1 $display("%b", po);
# 1  pi=207'b100101001001101101000010100101101011010000110111110101110000010010000000001010000111101010101011111001111011101100101101000011000110101100011110010000000011000010010001000111011000111000010101111100010110110;
#1 $display("%b", po);
# 1  pi=207'b101110111111101111101010001011010110110110101000011011111001000000010001111101011101001100101101010111000001000111110111001001011010110100001001000010110100101101010000110110111000111010011111011010101011100;
#1 $display("%b", po);
# 1  pi=207'b100111010000011000001100010011001110000011100010100100000000010000111011000010101101011110000011101101010000101101100100011101000001001111010011001101001110101101100010100101000101010101011010010011110100100;
#1 $display("%b", po);
# 1  pi=207'b110101100110100010010110110111100101101110110010111111000101110001010011100011100010001100011011111010111101010111110000000100100101100111001110010111010111100010011100100111000100001011001001011101000001110;
#1 $display("%b", po);
# 1  pi=207'b000010110000001111100010011011111101111001110110101100100001110011110010000100010111010000000110101011101100010110000111000001100101111110011100111000100110100001010101011100011011100101101011000101010100000;
#1 $display("%b", po);
# 1  pi=207'b101100100011011010101010101100001101101001000100110010000100101101011000110011000010000100100000001010000101101101010101010111100111001110010101100000101001101111001111100101111000100110011101000110100111100;
#1 $display("%b", po);
# 1  pi=207'b110000011000111111001100111000110010111000111110111110000100011111011011011110100000000110010001110010100011010111111011000100110011111111100010011010110101101000010111000011111001011011010000000001111001010;
#1 $display("%b", po);
# 1  pi=207'b100100111111101100110110010110000101100111110010000110011000011100111010111001100001100100100010000101111100001101100000101101011001101110110010010111000101111001100100101110000000101101011111100011000100000;
#1 $display("%b", po);
# 1  pi=207'b000101100101010001011111101110101001110100111010111101010100110101000101111100110011110000110110001011000111101100110001110100111101010100100110111101000011001101110101011000110100010011010111101000100110111;
#1 $display("%b", po);
# 1  pi=207'b100000110001010100010010011111111101100100100000001111110101101110101111011110101110100110111111101011001100110010000000101111001110101110010011000100001001000011110101111101011111101110000001110101001100111;
#1 $display("%b", po);
# 1  pi=207'b001001100010001010010001010010101101010101001100111001110011101000110110101110101010000010000101000010010111110000001001100111010001011101010110111101101011001100000100000100100001011101011110010101010110001;
#1 $display("%b", po);
# 1  pi=207'b010000101101110110110011101011100000010001101011010010111100011001011000001011010101010111100110011111111001010101001101011011110101001100000101100100101010110001111000001100100000111010110110101001001001001;
#1 $display("%b", po);
# 1  pi=207'b100101001000010011010110110111010010101100010000100001110000000110110110011110001010011010010001100110101001011000001101011110000111110011111111111101011110011100111111001111100000111110111111100001101000011;
#1 $display("%b", po);
# 1  pi=207'b100110001001011010000101110011000100001101100011000101111110011011001010010010101101111110001100100100110110110010001000100101010111010001101111000011001111001100001010101010101000110010010010001000001101100;
#1 $display("%b", po);
# 1  pi=207'b111000010011100110100111111101100010111001100000001000101010001110110000111010011110111011011011111000101000110110111100101101110111101110101011110111111011101101000001011000001101100001111101100000001010011;
#1 $display("%b", po);
# 1  pi=207'b000011010100000111100011110101110010001000110000110001101011101101010110100101001111111110100100000000010010100110101001010001001111010011110111001000110100000110000110011010111101011001011101000001000000101;
#1 $display("%b", po);
# 1  pi=207'b001010101111011001110010010011100000010000110011011010011010010000111010111111011111010010001011111111001011110110101101100001011010100000100000110010101010101101001011000000011001100010100101011100110100011;
#1 $display("%b", po);
# 1  pi=207'b101101101011100011010101001010011101011111111100000001011011110011101111111000101101001000000111011110000100000011110100111001001010011001100011111000111111101101010000101100011010000100010011110100000010111;
#1 $display("%b", po);
# 1  pi=207'b101100111110000001010001100010010110010001010101000000011000100100001000011100111010111001011100010011110100001001011101001101100001101111110111010001001001000011101110001000000001010111010011100011111110010;
#1 $display("%b", po);
# 1  pi=207'b011010011001010000101101101000101000000001011100101001100010001000011101001101101110001010110101000010000010101010010101101010010001100010001111010000010011100010101000111001011001110000001011000100110111100;
#1 $display("%b", po);
# 1  pi=207'b110111010111111100100100101111100101001110100000000110000111111000100010110000111100100111111111101110011011110111010101011101011000101001000100100110110110010101000110011111101100100011010110010010001111101;
#1 $display("%b", po);
# 1  pi=207'b111101110110100100000011111000000010110001000100010110000110011001010111011000010001000100000101001001001010110101001000011101101000000101001111010101100000101011100100111100111011101110111110001000111000001;
#1 $display("%b", po);
# 1  pi=207'b000110000111010010010011010001000010000111001001001111100100101110000001000111101100110111110001110100111101010101100010011001000000100101111100101111001100110100010110000010100110001010011001101000010101110;
#1 $display("%b", po);
# 1  pi=207'b001000010100101111111001001110011000000010100001000011001110011111000000110000110010101001010010110011111000011010101000101010100001100010010000110100111111001111111000100111000000111101001101000001111011110;
#1 $display("%b", po);
# 1  pi=207'b101101110011101100000000110000000001111000000001101010111000010100110111000001000001100100101101010010010011111101011111000011100111111111100000100100110011110111000010101001110110110011011001001011001111001;
#1 $display("%b", po);
# 1  pi=207'b000000101110110001110110011110111000110110101011010101101101011011100001110001101101000011001010111111110110101110000101011011100111000010010110010111000110000100011101010111100110011110111010111111101100011;
#1 $display("%b", po);
# 1  pi=207'b010011111110010101000000010001010000001000110001010000110000110101010110010010000000000001001101101001010011000111011000100001100010000110101111111011001000010001100001011001001010101011110101101011010110100;
#1 $display("%b", po);
# 1  pi=207'b101011001000110110011011100011110111111101000101000011000101111010100111010111011001110011101010111100001110100001000001000010111001011000011111110111010000011011100000101011101110111110000110010011001110100;
#1 $display("%b", po);
# 1  pi=207'b010110011110111111000001111001000111000010010101111010001011111101101010111011011101100011100000001100111100111001001111101101111101011000011100000110110100101010100011001001110110001100000111101010011101110;
#1 $display("%b", po);
# 1  pi=207'b100100111111110010100100110010100001100100101111000010000011011110100010110100000010011010010001010011000110111111111010000000011100111010110100110111000101011101111101011100000111100101110001000000001011101;
#1 $display("%b", po);
# 1  pi=207'b111011101100010000010001000111110110110000011011000010001111000010101101110010010101101101011101100110011110011101010110110111101111010011100001001011011000010101000100000111000011110001111110100001010101000;
#1 $display("%b", po);
# 1  pi=207'b010101010111101101111011011001010000000011001000101100110001110011100010010000000001100010101001000011100111000000010010100010001101111000100001000111101110111000010110110111110000001100110011000110000101100;
#1 $display("%b", po);
# 1  pi=207'b100110100100000110110111101011110111000110010100000010111101001010010110100110010100101111000010101100100111011111111010000010110111001000000011111000111101001111001110010000101100101000001101000011010111111;
#1 $display("%b", po);
# 1  pi=207'b100101010101110011100011111001101101100000110010100000001011111000010011111000000000111100101111011011110101010010110010111100011000111101110111011001010011010000101100110011000101110001100010001100011010011;
#1 $display("%b", po);
# 1  pi=207'b100100001011100011110000101101010111011110110000010101001010111011101010110000111011000110010100101100000101100110011110010100000001111011110111001110101000001111110111110110101001010010110010010010001010010;
#1 $display("%b", po);
# 1  pi=207'b110110010101110111000001000111011110010000100011101110000000101011010010000100000001101100001111000100000000110001011110001111010111100100001110001110000000111001110111010101011001110100000110111010100110110;
#1 $display("%b", po);
# 1  pi=207'b101010011011111010001011011111111000011100111001000101010101100101110011100101110110101110111010011000010001011100100010101101011010000110101011001001011010111101001011001001011010110010100011010001110101111;
#1 $display("%b", po);
# 1  pi=207'b010110101100001110110110010010001001101101110110110001101111001011000010110111001110110010001101101001000101101011000110000010010001000010111000000001100000010001001111011110111010001000011100111100110111010;
#1 $display("%b", po);
# 1  pi=207'b011101010101011101011010110010011101001101011001001110010101010101110101111000000001111001001101100010011100001100011011111110010101111100111101101100110010001011111010110110001101111101010101000100011011010;
#1 $display("%b", po);
# 1  pi=207'b110101110000101011000000101110001001110011011110001000111101100000100011101110010000010101110111100100011000000010111011111110001111011001001001101001110101110110101110000100001101101110111111010011000111001;
#1 $display("%b", po);
# 1  pi=207'b011101101111000010111101001101001000000010110101100110000011111011010101011101101001001111010100000010100110110010011111001001111011000111010011010011000100000000000011001001101110111000011110100111001110110;
#1 $display("%b", po);
# 1  pi=207'b111100001001111100011001101110000100010001101010110111011100001000101111110011110110101100111101011101000101011001000100011000100011010111101101110111101011001000101001101010010100010100101010011111000101001;
#1 $display("%b", po);
# 1  pi=207'b011100001100001011000010010111100100111011011100101100110000000001110111101101100010100001100001011110110101011111101110101110001000111111111001101001111011001000110101111101111001010000011110101010100000000;
#1 $display("%b", po);
# 1  pi=207'b110000011000001000010010001111110100101100011011000100010110000111100101001100001101100111000111100101110111111010011001100111000110001111100111010110000110110101010101011101100011100111001100000011111010011;
#1 $display("%b", po);
# 1  pi=207'b101000110111000011111000001110011010110111001000110000001101000010001010110010110100000010000111000111110111100001101001100000010000010101011101000101001000110010101110001000111111011010100101101010100100001;
#1 $display("%b", po);
# 1  pi=207'b010000101011110110011001100111111010001100000011011000000011000111110010101101111011101110000010001110000100000101100001110110000110010010000011110000111010000100100011001000110100001110110000101011001100001;
#1 $display("%b", po);
# 1  pi=207'b001001101100011101101101010001111010111101111100101001001010100000100000000001111001011001010010011001011010100010000010110110011001111010100001011100010011100000001011110110011000010001010001101011101010000;
#1 $display("%b", po);
# 1  pi=207'b100001100010010111110000101101101000110011100101101110111111001010001010010000110010011110111001000010011101101110011111111111101010100101110111011110110111110011011011010110111011010100101010101110111100000;
#1 $display("%b", po);
# 1  pi=207'b111110110011011011010101011010001000110100011110111000111100111111111100110000000101011000000001011011110100100010100010011011011110101000011010000111100110010100110110101111001000111010110011000001100011011;
#1 $display("%b", po);
# 1  pi=207'b011010010100000111110111001001000101010110101100101101000011000111000111000011101001110111100100001011100011111000110101101001110001000110001000010001000011111110001110101101110010111011100000111110000100111;
#1 $display("%b", po);
# 1  pi=207'b001100110010100011011001010101111001111010011000100010101100100110111001010110010101010001000011010011111001110000100111111001110111010100010110100111000101011000010010001111110001111001101101000001000100011;
#1 $display("%b", po);
# 1  pi=207'b101011110110111000001111000010011000110001110010110110111110110110111010110100100010010110000001001000010001000100101110110001011010110111000001001111100111111000110001111010010101110101000111000110010110001;
#1 $display("%b", po);
# 1  pi=207'b100000111010101111000100000011101100001010001011011110000101101011011111101110010000001110011100111010010111100010010111100001100010010111011100111001100011001110101000000011111010100010001011000101011100001;
#1 $display("%b", po);
# 1  pi=207'b101010101100100000000101011110110100111010010000010001001111001101111101000111001010101101110111010000100111110101100000100110111100001000110111011010100100110111000100001010101011000111011010111100000111100;
#1 $display("%b", po);
# 1  pi=207'b100111101011000001100010110111000000110010110001001101110111100001011100010100111000111100111010001100001000001111010111010010011001110011000100111101011000111011010000001010000010011000110000010111100111100;
#1 $display("%b", po);
# 1  pi=207'b000110111011000011011011111101101110101101110010100111101010111111100111110000100101010000100110110101010010100111000100100100011000101101111000010010110100010100101010100101110111001100111111010111010110111;
#1 $display("%b", po);
# 1  pi=207'b111101101010110111111101110101010011101111000001100000100111111001011110110000000011100011011010111011011100111110001111100111111100110101111011101111110010100001011110001111001110010000110100110110010100101;
#1 $display("%b", po);
# 1  pi=207'b011111110110010101111100101100010011011100100110101011101110010001011101101111101101000011001000000001011110101011100111110000000000001101100110101110100000011000101001100011011000100101100001101111001101110;
#1 $display("%b", po);
# 1  pi=207'b001000001110001010001101001011011110010001110001010011010100101110110111001001000011001001000000010101010101110000000111101111110100100100110110111001111010111100101010001000001101011101010101001010100000111;
#1 $display("%b", po);
# 1  pi=207'b110001101111000010111001011100011010000100101010000110000001000011101000001101011010111110101001111111001001010011110010001001100101100111010001100010100011111000101001001110010010100000000111001010111110101;
#1 $display("%b", po);
# 1  pi=207'b010011000100111010011000111010111110100110101101110101100011000100000011110000110101100010001111000000111010100101010110001111000011000111000000100000111011111100000000101110010011001011000000011010010110101;
#1 $display("%b", po);
# 1  pi=207'b101001100001111101100000010001101101001111000010011111110010011101110000001000110100101010111110101001110000000010000011000100110101011110010010011100100101101011010011110100100010100011001000001001010011111;
#1 $display("%b", po);
# 1  pi=207'b100110110110110011000100110111010000010010111101011011100100000111100111100101110001111110100011011011000010101111000111100110010100010010000111110011011100011000110110011001001111001010011001100100000110110;
#1 $display("%b", po);
# 1  pi=207'b001001011010101111000100100110101110110100010111111001001001110111000000001000010101100101101011011000001000000000001110001101100011110100010110010000001110100010110001010001000111001110101110001001000100100;
#1 $display("%b", po);
# 1  pi=207'b101001101100010000110011011101011101110110011010111000110001111011000010101100010100001110011011100101011101101110011011110010100000111101110101011000000011100001000110100101010111010111011011011101010101011;
#1 $display("%b", po);
# 1  pi=207'b001101011101011010001001101101011011011100111011100000101011111000010000100111110100011011101110000000101010101001001011100001100110000100100000110111000111010111101000111111100010001010010110001100101101000;
#1 $display("%b", po);
# 1  pi=207'b001001010011001100100000010001010001101001111111100001010001101110000010011000001001001000010011101011101010011100000001010010000101110110011000100110111010000110011110110010000110101001010111001011000001010;
#1 $display("%b", po);
# 1  pi=207'b101001101010101110010010001011001001101111010000110010100011000111011110000011110110010101100100000010000100100001001001000100011111100100010001100101001100101011001001000100101011110100011001101101101000101;
#1 $display("%b", po);
# 1  pi=207'b101011101010010101000100110010100011001000000100101100010000010010100111110111001110000100110010001010100010001000011110110001110110000110100010111001001100010110001010100101111110010110101100111001011110110;
#1 $display("%b", po);
# 1  pi=207'b011001011111101011111010101000010010111100000000001111011111101010100001011110100001001011011010100001111000101010111101100001011000011100001111001000001011000010011001000100110101000100000111111000000101010;
#1 $display("%b", po);
# 1  pi=207'b011010100011100011110001111010010010010010011000110000111000110111100110100100010010101101000010101101100110000111001000101010110111011100101011111100000111111011011010101011001011010101101100000000111110010;
#1 $display("%b", po);
# 1  pi=207'b100101011110010110010001111110110111010111110001011100001001000111010100001110111110000110111110011011010101011110000110111110110111110110001001010010111111100000001010110001010011101110111110101010111000110;
#1 $display("%b", po);
# 1  pi=207'b101101010100011111101010000110101011111101011100010100011111010011010111101111101000101010000010110111001110101100100010010011001001000100000001000100101100101110100111110000101000110010110110010001110101001;
#1 $display("%b", po);
# 1  pi=207'b110110110110011000100100011101101100100000010101110110000010111101110010110110011100100001011111010100101101011111110010101001100000010111101100011100001110100101101000111011000101111010011111011101000011000;
#1 $display("%b", po);
# 1  pi=207'b110010110110001000011111111110111000111000011111110001111000111000000000111001110011001000111001001001110001001000000111001011100110010010111000111001011100010000111011000001100001100110111111000100100111010;
#1 $display("%b", po);
# 1  pi=207'b101100111010011010101110101111010000001010111001011001011010000011011001001011011110111010010111101011010110110100101111110111110111100111100101010111011010101101000100110000100110011000100111110001100010111;
#1 $display("%b", po);
# 1  pi=207'b011010010011100001111011100110001001001001100111110110110011000011011010100100111100111110101001110010100101110010010010011100000111100111011011000001010000011011010110101001000100101111100001100101000001000;
#1 $display("%b", po);
# 1  pi=207'b011110101010010101010010011000000100111100000011011111010011100101000011100111001010110001010110011000110100110101111111000000011001100110100011001001001011010010010101001000011111110001000111101001011101110;
#1 $display("%b", po);
# 1  pi=207'b010010101110001110000010010101111000010101000010100001001011001000010011110001001010010000000011011101110110101110111110001001000110000011011011101100011000000110010001100000010010001100001011100101110010100;
#1 $display("%b", po);
# 1  pi=207'b001100101101001110101011110101100001110010100101110110001001101111100100100001111110000001011011110100010001111101111110101000101111111111111011011100101110111101110101100001110011001010000010100110011100101;
#1 $display("%b", po);
# 1  pi=207'b100000001100111000110100111110011000101110001100101101011001001100111011011001110100010101100000010110010110110001011001000111110000000101000101111111000001001100111010111001010100011100101001110010101001011;
#1 $display("%b", po);
# 1  pi=207'b011010011011011000010101011011100011001100111010001011100110100110001110110011000000101111010100101100101010110010001100110101011001011101001110110010100110111011110111010100111000000000011111011111001110010;
#1 $display("%b", po);
# 1  pi=207'b011000101100101100110101001001011101111111111001000101101011111110010110100101111111110111111011011010111000101010111011101011100011101011111110110101111110010011010110001111000101101001000111011011111101101;
#1 $display("%b", po);
# 1  pi=207'b111110010110001001001110000111101101101101001101111010110101110010000110101110111111000010011001000001111011110010011010011100100010111001110011110010000110110110110001011001111011111010011100101011000011001;
#1 $display("%b", po);
# 1  pi=207'b001100011101100100100001111110001110011111110010101100011001000000000001111110101111010101111010011100111001100110110011011001001011111111001001001110110110110001011010001001011101001111000001100011000100100;
#1 $display("%b", po);
# 1  pi=207'b110011010101010100001100000010011011001010011000001000110000010010111001100001101000100000101110111110111001100000111111110010110100111100110101000111110001011100110010000001011111100110100111001010100010001;
#1 $display("%b", po);
# 1  pi=207'b001011110011010100010110001001100000001100101000001100110011101010001101100101001101101010101110001100011101001101000100100101011111101100000000001110100001000100110011111010010100111110001000001111111111100;
#1 $display("%b", po);
# 1  pi=207'b001111001111111100010001010101011111111000111110100111000111111100101010110010000001110100010110111100111111001011011111111100001010011000101010100101101100000100111110100110011100110111011010110001101100010;
#1 $display("%b", po);
# 1  pi=207'b011000110110100010110110111101111011000110000101011110011110011100001001001111001101100110110111010100100101100010010100001010101011001001011100010110110001000000110111110011100100010011101011101110101101001;
#1 $display("%b", po);
# 1  pi=207'b111100001001100000010001001110010101000010011001111101100011101000010111110110001100111101001001110100010101111110110100011100111000111111000100011110110111001010000111111011011000010100000100101100011001101;
#1 $display("%b", po);
# 1  pi=207'b001100010010100101111010110001010001100001101011111110100101100011111000111001000011001010011001110100111010001000101101000000111001100110101101011101101100010001110100111010100110101001001011000010010101001;
#1 $display("%b", po);
# 1  pi=207'b011001010100100101110110000101000111101111001010111001001000001011011011011101010001001001010001010011000111011110101010011010100101111001111001000100101100010001010101010101111000001110010000111010010110001;
#1 $display("%b", po);
# 1  pi=207'b011100011000001101110111001111011011111101100000011010011100100101100110000110011100110101010010011000000100001100011011001000011101010011011110001001100010110001000100101100000101110001100000001110100101000;
#1 $display("%b", po);
# 1  pi=207'b011100110100110011101000100111110100111001010100110001101100111100000010000000011010011101101000011100011110010000011111101101001000111011011011001000101111001010110110101101000101110000010111000001111010101;
#1 $display("%b", po);
# 1  pi=207'b011000100001111101111011101001101100111010011101010001011011010110110110101001111010011001010011010111011100000101110010011110101000000100010111011110110000011011000001001111101000010100001001111101011111101;
#1 $display("%b", po);
# 1  pi=207'b010100011001101001000000100000101000110010010001101011110011100010001110011010000011001100110000001011101000010010000000010101111110010000010110111000001010101001011001010111100011010101011111111010001111111;
#1 $display("%b", po);
# 1  pi=207'b101110101111010110011100101001111000001011000100100000110000010011011010011110101000100000100111001001110010011000101001110100110100000000001100101101011101110010001101010101100011000100111101111000100100110;
#1 $display("%b", po);
# 1  pi=207'b010101100001010100111001101111000100101000101101101010000011110100011011011100101100010110001011010010011010010010001100011001000000110010010100101111100001100011001001111110101110111110011011101010010100100;
#1 $display("%b", po);
# 1  pi=207'b111001110011101111111100001101001011100001110001101111101010011100000010111010110011001010011011000101000101100011000111011011010100000010000100100111101101010011111011110100010011101000111110010010001110001;
#1 $display("%b", po);
# 1  pi=207'b000011000011001000000111011110000101010110110011100110101000011110111111100111010000000000110100000011011011101110000001110011000000000000100010000110000000001000101010100010101001101010010100001100000101010;
#1 $display("%b", po);
# 1  pi=207'b010000010001000110110011100101110001100100011001100001011110110110010101110111011011111100000010010100110101001001001110111101101110101100100011111111100001100111111100000010111101100111011000000100111001000;
#1 $display("%b", po);
# 1  pi=207'b000100101010010001010101011011110111000001010100111001110001100000001101000010011111111110110111100011101100000010101111111110101001101100001011110110011110100111010001010010101100000111100101011001100101011;
#1 $display("%b", po);
# 1  pi=207'b010000111110110011000100100000101100010001111100011010011100011011010101001100100001010011111011110010000101100111010101101001110100001010000111010101100101010101010110000111001011010000111000111010110011100;
#1 $display("%b", po);
# 1  pi=207'b000110000001111010011011011111010011111010101011001001101001000001011110000111001111110100100111000110011110010111000011011111010101000101101111011110110110010000100010000001010110100001000011110011111010100;
#1 $display("%b", po);
# 1  pi=207'b101111110011001110110111110111111101010010111011011100111001001100101111101110000000010001000101101010010001010110101001010101010110111111111110101100100000001011010110111111111000110111000011011111001000000;
#1 $display("%b", po);
# 1  pi=207'b111010011111000111100111000001110111110110110111101110100010110101101100000000010011101011100110011010011110010011001100001111101100000001011001110000000011000001000010000000110011011100101111000001000000111;
#1 $display("%b", po);
# 1  pi=207'b111010101110010101001110101100001110100101000010000011101101011000010011000001111001101000101100011010000010001010101100111010101111001000011111010000011000011101000100011100100000010110110111111010010011010;
#1 $display("%b", po);
# 1  pi=207'b001111101001111010100101110101100101011000011100000001001001000110010100001101101000100111100010111001101111111100100001110010011011010010000101001000110011010000110001100110100011100010111010111110101010011;
#1 $display("%b", po);
# 1  pi=207'b000101111001101110111010001010101001100110101111000010101011110010100001000101000000111101111010001100001100110001100101000111001011110010110111111110010101010000011000110110111101001110101100010111010101001;
#1 $display("%b", po);
# 1  pi=207'b011010010001011110100100111011001101011111000110010010000011000000000001101001011110011010010011111110011110100110101101010110000100000100010101110000110111111101000011110111111010111010000101001111100001100;
#1 $display("%b", po);
# 1  pi=207'b110000100011100011010111100111000111110100011110111011010101010010010000011001000111100001001010110101010001000100010011101111101000011000101001101010010110111100011000011101100100001001000110101100110111111;
#1 $display("%b", po);
# 1  pi=207'b101011110010011000011110010110010000101010101011110001011101100010111111001001101010110111000111001100100010100101111101101001100000110110111111011100110001000111001010010101000110111111111001100101010100100;
#1 $display("%b", po);
# 1  pi=207'b101010110011100010010110110011100000110110110000010010100011001001010011001101000010010010011111101001010001010101010101000111101011001100110111010100011111101111011111010010101001111110000001100011010100000;
#1 $display("%b", po);
# 1  pi=207'b110110011100001100111010010101110110101101100001000000000000011101010110111111001110000000101110100110100100000011100000010010111100000110010000010100100101100101101011000000011010010011011100010000011101011;
#1 $display("%b", po);
# 1  pi=207'b010111111111101111011110000100101101101010100001011100110010011111111110010010110100011111000010111110011110101001000101101011011100001000100110011010000100011110011111101110000001011110101011001011111100101;
#1 $display("%b", po);
# 1  pi=207'b111010010111011111101011001000101000100001010000010100011111111000111001101011111010011001011011110001110001001011100010100000110110001100110110001010100010010101011000010111111011100110110010101101000111001;
#1 $display("%b", po);
# 1  pi=207'b101011010011100101111101000101001101100010111101110000101000111111000110101011010100000011111101110110011011001011100100100000110100000110010111110110101011000100101101100110110011000001010111001110000011101;
#1 $display("%b", po);
# 1  pi=207'b111010001011101110010100110100111101000101110111111001100111011100100001100111001001101011110111110100000110011000011011010110011001001111111010010011010111100111000110101001001011011000001101011011011001000;
#1 $display("%b", po);
# 1  pi=207'b011111100100111001011010001000001010111101001110001010000100001101111010101101011000001110100010011011111111001101100101000110111101111111000000101110010100001010011110111101101011001110011010011011011000111;
#1 $display("%b", po);
# 1  pi=207'b001110011111100111001001110101101100111010101011001011101011100111010000101010100011111100011100110111010011000101100110101010101110011000001101011001010111111001011010000110101101011100101111011101010000110;
#1 $display("%b", po);
# 1  pi=207'b101010010010001111111010100100011111011001111011111011001001110111011100101001110111100111011000011101101111101001001010110110011100100110001011001001000110111111110100001111001110101101100111010101001001111;
#1 $display("%b", po);
# 1  pi=207'b101110001000010001001101010000010010110010110101111101000011100001001001000111011101011101001010010000101110101010010011110111101001011010011101010000011111000010011001110100010100111100101011010110000000101;
#1 $display("%b", po);
# 1  pi=207'b000111100100010001001111010110111100101001101000111010100010011111100011010010101111111001100100100110001110001000011010001101100110000101111110001000100111010110000100001010110001110000011011000100101110001;
#1 $display("%b", po);
# 1  pi=207'b100000011101100100011110010011010100101110101000011110110000010001110010000101100010100101010010110100110110001010011100010100111111000011000000101001100001101110010110011000111100011101011100101101010110011;
#1 $display("%b", po);
# 1  pi=207'b111101010001101111010101000110110101011001010010100101000100110111101110111010001110101101110101101000011110011101011111100100010100010111100110101010000111010100100101001001011010111000000100111111100111011;
#1 $display("%b", po);
# 1  pi=207'b100001100011000000001100011100111011000011011100001001000110010100010110000101110010000101011010111100001101010001110110110000000000011101111111100111101101111100000101110001010110101001000110111011110000111;
#1 $display("%b", po);
# 1  pi=207'b011000101110111011111111100100010111011001001101101111001101010101001001010111100100100010111001111100110001000001110000110000101010001001111101111000100011001011011010010100111111000111110011101100010101100;
#1 $display("%b", po);
# 1  pi=207'b100110111100101000001101101010100110010010101100001100010001010011000000001110101001100110111110001000001001000010110100100101110011000001110110110101001100100010101000001011000011001010011110011001000001101;
#1 $display("%b", po);
# 1  pi=207'b100010100010110000010100001011010001101001011101100110001011100100001001010110000111110001111001111100000100111100011001011100010000101010101110001011101111101010110001001100101010010010011000101011111000010;
#1 $display("%b", po);
# 1  pi=207'b100111110011101111010101101111011100001101101011000010100000010111111100010100001011100010000001000100101101010101010000011011000111000111000100100000010001110001110000110100000001011101011111001000011000100;
#1 $display("%b", po);
# 1  pi=207'b110101100101110110111100111011010001000110010000001100010011100011011010110110001100011101010010001100110010000110001000111011111100011001001111011110001100100100011111111101010000011101111000001001101000010;
#1 $display("%b", po);
# 1  pi=207'b000111101001100111110101010100111001101000111011010100111101111111001110011101001111111100101001111101001001111100101011010000100010100110110100101010111011111111101001100000111110100110101110101100011110000;
#1 $display("%b", po);
# 1  pi=207'b111011001000000110110010011111000001101001000001011110101000100100110000110010001111101001000101100001000111100011011110110011010010111010010100011011111100010110011000011101000000001110101110011011100000000;
#1 $display("%b", po);
# 1  pi=207'b111110101110100010000100011000111111100010001101001110001001010111100111100101010010100111100110110000111111110010000001111100110001010011111110101101000111110011100010000010100010110100111111011010111110011;
#1 $display("%b", po);
# 1  pi=207'b111010010000001011110101000010011100101101100100010100110110110110010011111001010100111001000010100100110100010110101010000011110110001100101101001001111011010100100001000000011101010101000011010110000100110;
#1 $display("%b", po);
# 1  pi=207'b010110000001010101010010111011010011101010011001111000010000000011010110111000000010001111010100010110111111010101101111111001000010110000010010110111110011011010100110110101111111010001101110111100111101000;
#1 $display("%b", po);
# 1  pi=207'b010110011110011010011100000010110100000001110110001100101000001000000110000001010110100000000010111000100011101101110100110110000001101110111101100101000111001011001011001111101100001010101001101011101001101;
#1 $display("%b", po);
# 1  pi=207'b111110101011000000001111101100010011000101111111111111000011111011101101001101010011101100010100111010101100110111110101001110110001111111001011010101000011011010110111000101011110110011000011011000010000110;
#1 $display("%b", po);
# 1  pi=207'b100100011101100110000001101010111011001000011111011001001100001100000110101011000101011101111110101010011101110001010001111001010000101000100000001000000001001101001000100001111011100000001110000100000000001;
#1 $display("%b", po);
# 1  pi=207'b111111011000011000000100000100110111010010111110111000100000011011111101011100011011010101100110110111111111101000111011011100011111100001111110110010001101011110101011100110111101011010001001100111011000000;
#1 $display("%b", po);
# 1  pi=207'b100011011110010010001011010101011100100100001010011001100111110010110000001000101100010001110010111001101101110000010000000111010000101011101001111011101111011011101111110111111010001001110000101011100010010;
#1 $display("%b", po);
# 1  pi=207'b111101000010010001001000000101011010101011011101001110111110101001001010100011110010010110000101101100111100010000011010000010101110111110100101000101100100011111000001100111110101110010100110001010011000010;
#1 $display("%b", po);
# 1  pi=207'b111100110000001101100110101110001001110000100010001111011111010111101100101111110100000111111100010001100100000111010001010010100100110111001100000010010111011011111011001001110010111100110100011110011110100;
#1 $display("%b", po);
# 1  pi=207'b010111100000011011001101101011000001101110100011000110011011000001101000100010001111111001110101101111111111100010110111101011010001100100010110111101011001011100110000111110000010011110010101011100111110100;
#1 $display("%b", po);
# 1  pi=207'b010011111001111100110011011010011000110011011100111001010100000011000111111101100100000111011100010000010011011111111100110011100111101110001010111101110110101011110101000100000001111101001100000100101100010;
#1 $display("%b", po);
# 1  pi=207'b110100110111110010001010010101011111100101111010001111010011001001010011110101111111000100010101110111001000000010100001000011010101010011110000001110101001001101111110101000001000100001010111010101001001111;
#1 $display("%b", po);
# 1  pi=207'b001110111010100100000010110110101000010111000110101101101110111100101001101011100111011101011110111001110101101111100101100110010111100010100011111010100100011000011010001000100001101011000111001101101010111;
#1 $display("%b", po);
# 1  pi=207'b111110010011011000100111010100001100010101011000010001011001011001110001011111111010101010100010111111011111011011101010111110000100010000011001101010111000100010011001010001011001100001000000111000000011111;
#1 $display("%b", po);
# 1  pi=207'b101011011000110000111000100111111011001010001111100110110011000101100011001110000001010110010000011001010111111110001010001001011100011010110111101100111101010000111111111110010000000111101101111100110000000;
#1 $display("%b", po);
# 1  pi=207'b001001100010111101110011010111010000110001011110111000011111011110000010110010000010001011101110010001110101111000111101110001110101000101100000100110010010100110011101101111100111111100000100101111101111000;
#1 $display("%b", po);
# 1  pi=207'b011000011000100001101010000111100011100000101010111010100001001101011100000010010110110001100101000000000000110011000000101001111000001011110110001010100110101110011100000000010000010111101010111000101110110;
#1 $display("%b", po);
# 1  pi=207'b110000110011111001100010001100100100100011011010111011110000001001010110100000001010101100100010110000101111000010111111001111100001000000000010100101111001010101000011001111011001101000011100110000011000101;
#1 $display("%b", po);
# 1  pi=207'b000011111100100111010101001100011001110100100001001000101101110000100011011011010000001101111010100100001111000111100011100011110000001010001010010000111000011111101110000110100111101011110101011000010000010;
#1 $display("%b", po);
# 1  pi=207'b000111110111101110010100100010000110010110100111001011011110101000010110011100100110011100111110110100001001101100100110100100010000001110110001100011000101110000010111111000000010011010001111101010100010000;
#1 $display("%b", po);
# 1  pi=207'b011001001011010011001110110001001110010100011001100110110010010010011101110110011101001000010001001101100011011001111101000001110101000101000001111001111011110010001000010000000011101100111111110010000111001;
#1 $display("%b", po);
# 1  pi=207'b100100110011011101001110010100110000000011000000001010011111110001101011000111011010101001111001110001100010110010111000101001110100101101100101010011100010111100010101100010111101001100110001000001001010001;
#1 $display("%b", po);
# 1  pi=207'b000100001110010010010001100100111111111010100111011001100000010011010000000110010101101101100110010010010110011100111000101011100101010110000100101111100100011111011011110011101010110001101100010111110101000;
#1 $display("%b", po);
# 1  pi=207'b111101010111110101100111011111101011111100001010100110111001100101000111011010011100100001110111101001011000000101011111011111101001000100110100001100101100100100010010011110010011010111111100011010010100010;
#1 $display("%b", po);
# 1  pi=207'b100111001001111001101111111010000010001110011110001101101100010001100110011110000111001111110101100001101010000110111111011110010100010000110100001010101110101001010000001100101101011001001010011100011100011;
#1 $display("%b", po);
# 1  pi=207'b000011110011101010000011001101000100111111001110100001011101101110010011111010011100010010001111111111100100001111000010101001000100101100000110110010110111011011101101100001100011011110011010110001010000010;
#1 $display("%b", po);
# 1  pi=207'b011000010111101000101101110011110101111011010110000001111111100010001011110111011000000100111000101101000101001011000101100011101000000010011001100111011000000101000011010001110001000110010010010010100100110;
#1 $display("%b", po);
# 1  pi=207'b111001100110111100000100111110100111000011110101000101101010111111010110001000011011111110000100111100110011010111111110010011010001001011011001011010100101011110010110000110111001000111111000110110110101111;
#1 $display("%b", po);
# 1  pi=207'b111101000110101110100010011111000110001101110000110011010010101110101101100011010001011011100101100111010000010010111000101001001000001000010111011111111010011011101100100010010010000001000101010101111010000;
#1 $display("%b", po);
# 1  pi=207'b000010011101111101011000101000100111101001111111000011100001101111001101101010100110001000000111001001000111000011000101010101010000010010010001110010010101000010010101011101001011101000011101011110111100001;
#1 $display("%b", po);
# 1  pi=207'b010001011110001000001111000011101000001111101000000111101011111001110011010100101101110011111101100000101010010010111111110111101001100110011110110010100011000101001110100101011111000101110100111001100111010;
#1 $display("%b", po);
# 1  pi=207'b100100000001000110000100110101110010101100000101001101001011110000100010000000100000010111010001010100100100100010001000010001100100000110010011011010101000010100010000100110011111000101001010011011101000100;
#1 $display("%b", po);
# 1  pi=207'b101011101110110111000000011011111110000000001110101101101111010110010101010111010100010000001111111111100011111110111011000101011111100000100010010000010011010101001100010110111100001111011010100001101110010;
#1 $display("%b", po);
# 1  pi=207'b010011110010000110011101011010110010110001001011001111111100010100111100000111100111100111010011110011011100111011110100001001111100111100011101011000110101110010111010101000111001000101001000001101011011110;
#1 $display("%b", po);
# 1  pi=207'b010011001001101111100100000110111000000000100110100011000000001011110000000101000111111001011110010100001000100110011110010111011101011101000111111000100111011001111101101011100010011111001000100100110010010;
#1 $display("%b", po);
# 1  pi=207'b100111001101011110001011010101110001101010100010000000001010000010101111011001100001110111010001111110011011101001000010110110111000010011101111000010110000111110001001110110000000110111111101001011001101101;
#1 $display("%b", po);
# 1  pi=207'b110101100110110000011101111111000110101101011000100001000000110011101100010101110011111100001011100111111011110011101010100101110100000101001011010100000011110100001010000011100010110011101011101011010011110;
#1 $display("%b", po);
# 1  pi=207'b111001110001101110111111101111110011111000100111000101100010111010110111111011001101111100010101001111101011101011001101111001010100100010110101100010011010010011000001010101100001011001010000010111101110100;
#1 $display("%b", po);
# 1  pi=207'b011110011111111000110111101101010100000010011100111011011001011001101111110110001110001011100000001100001011101000111111110101001000110000101111010111011110011110101000010100111100111000000011110111000110101;
#1 $display("%b", po);
# 1  pi=207'b111011100101011001000100101001010000011011000000011001101110001111110001011100110001100001000001110010011100110001000111001011000001010000101001110101000111111011001111001101100011010100110010101101110011011;
#1 $display("%b", po);
# 1  pi=207'b010011001110111100001100001011101101111111111000000001101101100101001111100111011111110111101011011001000111010001001000101100011000000110001111111000101101110010110000111101010000010111100110101010001011010;
#1 $display("%b", po);
# 1  pi=207'b010101011010010111110001101100111011001111101111111010001101010001101100111001010001100111000110001011000001111111011101110100110110001001101101101100101110100011010100101101011101111101010011011111000101101;
#1 $display("%b", po);
# 1  pi=207'b101100010100111101000100001010110010110011100101101101000111000011100101110010101100001000000011000011011111010111001101011010110001000100011001110100111101110011100000110001010111100000011111010001001110110;
#1 $display("%b", po);
# 1  pi=207'b011110000101000001000111110010110000001101111100100100110111100110100000001111000011100101100111111001100111111111010110101010110110011110101101111011010100010010011100110011010100011010011111101100000010010;
#1 $display("%b", po);
# 1  pi=207'b110011101100011000101100100101100110010000101100000100011111011001101110111011010000111101100101110010000001010000000010000001010010110010110010011100011111001111000001000100110011110010111100000101100001010;
#1 $display("%b", po);
# 1  pi=207'b011100100100111000111000000101100100011001000100011100110110101001011110111010101000110010101100001111000110011100011010110011111001000111110000111011000111100001111111011011100000011010000011011101001100001;
#1 $display("%b", po);
# 1  pi=207'b101101001111001000111101001000111100000011010010010100100111110101110111010001101110011001100111111101000000101101001100000111111000010111001000010011100100110100100111000101110111101110010001100110100111100;
#1 $display("%b", po);
# 1  pi=207'b011101011110111101010010011111111010110010111101100101010011010110011001101100110101100101110100101011110101001011100010111010000000001000110001111010111110110010111110110000010100000111100100010111111011010;
#1 $display("%b", po);
# 1  pi=207'b110000000110010101110001101011011111110000000001001011011000101001110110001011001101000101100111101111111010001000001110100011001010110000011010111110100011101000011011001000111000011100101101111000101010111;
#1 $display("%b", po);
# 1  pi=207'b100000100000011011101110110001111100000110110000010110001101001101011001100101000101100000101011010111011101000011101101011010000011000011110010011000001011111100011111010111000100111011110011001001110010011;
#1 $display("%b", po);
# 1  pi=207'b111011001000011100101000101010000000101100011011001111111000011111111001101111011101011000110011110010001000011011100111111101001011110110101000100001011001011110001010001001101100000011001010101011111111111;
#1 $display("%b", po);
# 1  pi=207'b111111010100111010001100001010111101111100100010100000100001100000010100010101100000100001110000000100101000011101101000001011000100000101001000101011100101101111111010010010110011100110000110111001011011111;
#1 $display("%b", po);
# 1  pi=207'b110000011101101100110010001001100000111000000110110010110001010001101100011011010011011011101010010010110011010111100011110110011101101000110100100010111110100001001101101010111011110101100000010001011111001;
#1 $display("%b", po);
# 1  pi=207'b000101011110111011000011110110001111111010111101011000011010101111011110011010000011010001110010001011001100001101000100100111101011101111010010100100001011101100101000111010001010000000011000010001010011100;
#1 $display("%b", po);
# 1  pi=207'b101101101010110110001111110010000101000110001100101000011000111000011101010111000001011101110000001110101000111010010111101101001000100100100110001000001100000011001010011111010011001110010100101101101101101;
#1 $display("%b", po);
# 1  pi=207'b000110000110001011111001101111110111101101011011101011101010100000010110000000110100110111000111010010001000100010011100101001100111010111011110010100100011111011011011110110010010101111110100011001011111101;
#1 $display("%b", po);
# 1  pi=207'b101110101000111100111110101110011100101100010110001010000111001010100000111001011001111111011011110010000111001111001010110100110101111110110110010001100111111000101110111010110011110110000111100111000011011;
#1 $display("%b", po);
# 1  pi=207'b110100111011011010000011011011000001010010100010110111010100010000101101011111011110100111110101011001110010000100011111111110100000110001100011010010001001110110110110011000111001111001111110001110101111101;
#1 $display("%b", po);
# 1  pi=207'b011000101011110010000111111010100101101011100101000000101010001100111000111000000100011101101010100000101001101001000111111001100001110010001110001111000101100100001010111100001101000111111000010011001000100;
#1 $display("%b", po);
# 1  pi=207'b110100000001101101110000011110100000101101001010011011101011111011111001111010100101111010001111010000100111010100110010111000011110101000101100000101110101111001100100111101110011100111111000100010111111001;
#1 $display("%b", po);
# 1  pi=207'b100100001110010110001010010100100001000111101000011000100000011100001010011000001010100010011000001100011101011000010110111011100000111101000100111111011011110001110010101000010010100101101001010011001110011;
#1 $display("%b", po);
# 1  pi=207'b011000111010011100010110100010101001100011100100100111010010010111000001101101110011111011010110010100011011011110101000010101100001010111100100001001001101011110010010011001011010110010011011111100100101011;
#1 $display("%b", po);
# 1  pi=207'b011011010000000101101111001101101111000100110101110111000101001101111110000100000000100110110010101111000100111100101011000101010001010111101011010000000100011001010010110111011010110011010100101010101101011;
#1 $display("%b", po);
# 1  pi=207'b101011011100011100100010011110111111011110101111011010011001111001111001110010100110011010010101001110010111111010001110110001010010000100101110111101000001101011101001000101100111101001111110001001110111001;
#1 $display("%b", po);
# 1  pi=207'b010011110011100101011010011110011010111101010001000011101100111010100101000000000010011100010000110000001011011010010100011101101000011010110001000111101000000011111101001000111110000100010110001000101001011;
#1 $display("%b", po);
# 1  pi=207'b101110011101001101011101100101111011111000101010011100001101001001100100011000001011110000101100111010100010010011111111110100111000001011010010011000010001011001101111000011011100110000010011110001001101000;
#1 $display("%b", po);
# 1  pi=207'b101001011100010111101000110101101010111110110000000101100010110100111101101101101010110010001110011111111011001011101111010111111101000011101100101010000111100110110000000001000011010110011010000011110110110;
#1 $display("%b", po);
# 1  pi=207'b001011000110010111110111111110011001100000010000110100110001101011101001001101011001110101011111100000011001000100111000011111011010111111110011110011101101000011000100101100101100000110110010111010100001011;
#1 $display("%b", po);
# 1  pi=207'b011101110000011001011010010101111011000101010110001011011000011001101111000001100000111111000101000110100100110111111011101011100011110011101010011111101000111101001011101101001110101101110011101011100101101;
#1 $display("%b", po);
# 1  pi=207'b111111001100111110111100100101111101101101010111100010000101101111100101101100001000101100110011001011111011100110101101011100100111101010011111010111010011111000011010111000010010001111101110110111001000010;
#1 $display("%b", po);
# 1  pi=207'b101100011111000101101110111110111010011111101001010101011010111110101000011001000011011110001101101001000101101000010100000011110010111010100110111101010000100000101100111001110110110111111000001001001100000;
#1 $display("%b", po);
# 1  pi=207'b110101110111100110110001110000011110001101111110011011100001001001001101110111001110100100011100101110101000101101111010001100000011100100000001101010100000101011011101110111001110101110000010000110001100001;
#1 $display("%b", po);
# 1  pi=207'b000001101010000100001000011110011111111000001110101100000000011011000111001100000010010010111101101000001111100101100100000110110100100100000001010010011001101010011101011011111010110101101000100110101001101;
#1 $display("%b", po);
# 1  pi=207'b000110000011111101010100101001101000110000001110010001000111100100000011001010101111101011010110100010001010110000000001011001101111000011111111111100010011110110111101101101011010000111101010101001001011000;
#1 $display("%b", po);
# 1  pi=207'b000110010010110001110001010010001110000100101101010011110000101101010111111001100010100001100100111111101010000101011101000010100111010011011010001101111011111110010010000001000011110111001111101001100100010;
#1 $display("%b", po);
# 1  pi=207'b110110000111111111001010011001010001101000001001001111010010000110100100101010001101011000111010100111110000101000000101101101111111111101110111011010010000100111100000111111110101111100011101001010100100110;
#1 $display("%b", po);
# 1  pi=207'b001100000011101010000000000101001000010000100000001101100110111011110111100100000001010110010011010010101010011101101110011010111111000000001101000000010000010110100011110001010000010110100101000110010011110;
#1 $display("%b", po);
# 1  pi=207'b110000110000100100001101001100010000100011010011000100010111111111110010000001100101010100000010001000100101000011011111011001010100000101010011000011011111111101111011010101010100110100000011111011110111001;
#1 $display("%b", po);
# 1  pi=207'b100001011010010011100000001011011100001010100001111111010010110001101110101111001010110011110001001111010100011011001101101100001000110100101011001011011111101000001000011101100011000110010000100110000001100;
#1 $display("%b", po);
# 1  pi=207'b111011101001011010111000100011100001100110101011110101011110010001011000011111101101111000111110011011110001101110000010011100000111011110100010100111011010001100001010111100001101011100100110011101101001001;
#1 $display("%b", po);
# 1  pi=207'b001110111110010001111100001110110010011011010001010010001011111101000011100010000001100111010111001000100001110111101111011010011101001111111110100011100010011000110010001001001111001010011101010111011010001;
#1 $display("%b", po);
# 1  pi=207'b010011000010110100011010100011110001101100101001100011100111100101100101000111000010000111010010011010101100100001100001011100010100101001101001010011010010001110110010111000101100110000100110101010100110001;
#1 $display("%b", po);
# 1  pi=207'b100001000001101101101011101001001010001011010001001011000101010001100101000011011011110010110011001111110001001000111001001000100001100011100010000101110010001000000111001100001000101001110001001000001101000;
#1 $display("%b", po);
# 1  pi=207'b111101100111101110100001111101000011101011011000011011011110100111101101110011000011110011011000110000101111101110000000101100000110011011100110100101000101111110000010001100111111010000100111011000111001000;
#1 $display("%b", po);
# 1  pi=207'b100111111110001110110010010001110001110000011110000101101001010111101001001010100110110011101000000100111011100010111011101011110101101011111010111111011001110011011111100101010000101000101010101110000000000;
#1 $display("%b", po);
# 1  pi=207'b110111000000011010100001110001111011111100110110000001111110000110000100000011011100001000100111001100101000001001100010111111001100011011011010101000101010111111100100111001010100010101100000111000111010001;
#1 $display("%b", po);
# 1  pi=207'b111110001011101000001000001110010100100110100010110111000100000101001010000000000001011011001000100110010011101000111010001011000011101100010010111111010010000101110101001110111001010111000101101000111111000;
#1 $display("%b", po);
# 1  pi=207'b110111001110101100000001010000111011001100100111100100000000011001110111000000000001001001001010001010011110001100111110100110001001001100101110111101111100101100111111111010010111000111110010100110001110111;
#1 $display("%b", po);
# 1  pi=207'b110101010010110110100110100111110000101000111110101001001010111101111101101111010010000101101110101000100101011101010111010111110100111000111100101001101011111100010110011000110000011001011001110100110110000;
#1 $display("%b", po);
# 1  pi=207'b101110101111101000110010011100101001001110111011110101010010011010000001000010100101011100010110001011101100100100101111101111001001111011010010110000100110111010101111110011000110000110101101100110011000111;
#1 $display("%b", po);
# 1  pi=207'b000110011101001011100000010010001010011010101110110111111100010011000111000011101100011100111011111110110100110001010000010100011010001100101001000110101001110010010110011110010001110100100100001101110110101;
#1 $display("%b", po);
# 1  pi=207'b110011010000000101110001110001111110101001001000010101011011001110010100101011001001101000111100111000011011011100100101101111100000011011000010001100110111010011011010101010010001000110110111101011000111010;
#1 $display("%b", po);
# 1  pi=207'b111100000001101111111100000001010001111010001100010100001101110100110101101101001110011101001101000101010001111100010100100000111111111100110101010110110100011110011101100000010000011001110001000101111111111;
#1 $display("%b", po);
# 1  pi=207'b100011000000010110101111010001010100000011000011001100100100001010001100110010111000000011100001111001011010011100101001100000011000101001000001111110001110100110010101101000100001111000110110001100101100011;
#1 $display("%b", po);
# 1  pi=207'b000101001101011001101101001000100110101011010011110000111000111010001011101010001000011110000001011101110110111001010010110100000101100100110111010011001100000000111000101111010111001011101010011101000010000;
#1 $display("%b", po);
# 1  pi=207'b011011011110101111110011011010010110101001101001111100001010110011101011001110111100101100010111111110100001110010011011001110100101010110000111111000101011101011011101110000101000001110100011101000100011110;
#1 $display("%b", po);
# 1  pi=207'b100011010001111110000110011001100111000100110010010011101000101101100010011011101001010100100101111100111101111001011100010001001010001010010101010111101011000101110100111001010000001011111011001011110100110;
#1 $display("%b", po);
# 1  pi=207'b000101110010100110100011010011011000011110100011000101010110001110100001011000011001001111011110111010100100101000100001100000100000010001000100110011011010000000110110110110001110100111011111000001001001100;
#1 $display("%b", po);
# 1  pi=207'b111110011010110101110110000011101100100101001010110100000101010010100100111001001001010001000110101010111011101011111010110110101010111110000110101100000010100000001000001001010011110000110001010101100011001;
#1 $display("%b", po);
# 1  pi=207'b011100010010101001111001001011110111010110100011001110101010011110110001010000010000010110110001101111011001010010010010111000010011011011011101011111100110101010100100100100011110011011111100001111111000111;
#1 $display("%b", po);
# 1  pi=207'b101001011001100010011000010000000100111101100110100000010010001000011011101101101001000001101001010110000111001001001011010100001100010010101100100100111101100110010110011111010000111010010101100101010100010;
#1 $display("%b", po);
# 1  pi=207'b101100000101011000011111001010110101100001001110111111010010011011101010101101100011011111110010111000010101110001010000001010001100111100101001101001111111000010001010001011010111110011010100001010010110100;
#1 $display("%b", po);
# 1  pi=207'b110011011101000100000101101110110001110011010010101010001110111001010001010110110100001000001010010110000000110101100101010001010001101101001110111001011011000010100011001101011110000101100110101000000100111;
#1 $display("%b", po);
# 1  pi=207'b101010011000100110000001111010101000101101001100011000110101101111100100000011010011001101010000011101011011110000110010000010100100101111000101001010110110000100100001010100101101111101011101111111100011110;
#1 $display("%b", po);
# 1  pi=207'b011000011111100101000000111011010000100101011000011111000110110100010111001111010101100101011000000100010000010111110111110110110111100010110011101010010001111010100110001100000100001010110010101011010110001;
#1 $display("%b", po);
# 1  pi=207'b110100110110100011111010011110001010111111110000011001101110100110100000010010100111000001100111001000001001110000100001100010000100100000000000111111010010110100111110010101100011101000110011100011000011010;
#1 $display("%b", po);
# 1  pi=207'b011101101101000111001110010001001100110101001100111110110010011001110110111111001000111000011100111111110111111111111101000100010001000010001100111010000111110110010100001100001000110111110101101101001110101;
#1 $display("%b", po);
# 1  pi=207'b001101001000000010110110111010110010100101011010010010110010100010101110001100111111111000000001110010011100011111010101011111101111100110000111100110001100110011101101111110110100100011101001101001001011010;
#1 $display("%b", po);
# 1  pi=207'b101011101011110010001000111111110000010110101010101001010100110101100011000001010100011001100101101101001111000000111000001010101101111001111100110111010111110111011111000111011000111111010011011010011101011;
#1 $display("%b", po);
# 1  pi=207'b011100111001011011000010010100011001101001100101111001100000000010101011111001011111011101100010111111011101101101010011100010101110100001000010010010000000011011100000000011101111101010011000100001000110000;
#1 $display("%b", po);
# 1  pi=207'b110001010111010010101010010001111000111000110001110011011100100000010000011111000100001111011111111001110010101100100010100011111110100110011001010001101110000010000101111010100000001101010101100110111001001;
#1 $display("%b", po);
# 1  pi=207'b101011001110110001001100000010100101010100000000101101100100101001000010101101110011111111100010011011001010001001010111001010000101010111110000001111010000100010000101111010010010111100110100010001101101001;
#1 $display("%b", po);
# 1  pi=207'b011111111101011000101010100101111010111100110001111101101111101101101111000010101010011001110001001101100010011101011101011110000111010100011000010100011010000101001011101100100111101110000010110111100011101;
#1 $display("%b", po);
# 1  pi=207'b010100101011110111010100111001001010001010001111111101101111010110000001111010010110011101111011010110011000101011110110001101010000101000101100101010000011011100001010101111000011111111110110000101010001110;
#1 $display("%b", po);
# 1  pi=207'b000001110111010010001011000111101011111100000101011000111011000101000010011100101001011101000000110010110101001101111110011100111000110001011100010010011011001011111101100110001100001001101100010101111011000;
#1 $display("%b", po);
# 1  pi=207'b110011110101111101110111000010111101010111010110011111011110101100011101011110001110011101010010010100011100110100000111011001111100100111010011010010010010010010111111011110111000010101010000011101010110101;
#1 $display("%b", po);
# 1  pi=207'b011011111110110011110010111001111101101101110010100111000100111100001110100011100010110100111111101100011110100010011100000000101011111111010101111110011011011010111110010001110110011011110110101111000000110;
#1 $display("%b", po);
# 1  pi=207'b010110111110101001001101010101110011100111001110110000100101101010000000111110111000111010100110110010011110111110011110110010010100110110111010111110111101101101011101011111010101101001101000101100110111000;
#1 $display("%b", po);
# 1  pi=207'b011000010111101011011111010100100000110101110110001011110001111001001011010110100000011100010101111001101100110100101001100101001001000111000010111011001100101000000001000000100000101101100111000001101010011;
#1 $display("%b", po);
# 1  pi=207'b010101111000110100000010011101001111000100011111001100010100000001101100010100010111000001001000011111010010011010010000001111011110011011010111010010010001011000001000011110011111000101010001111110001100010;
#1 $display("%b", po);
# 1  pi=207'b100110101010010110111101100100000001000100101111100010101000010111000010101011001000101100111110001001100000100011111010011110101001010101011000100101110001010101011101001101110011000111000111100100100011101;
#1 $display("%b", po);
# 1  pi=207'b010000000111111101001100011100101000000011001111001110010100001101010110100111010001101011001100100111000000110111001101100010110010110011110001000111010100000001010101000011000000011110010100110101010011000;
#1 $display("%b", po);
# 1  pi=207'b101011010000010110100010000110000011000101100100000000111111010011110101010011101110101010000011100001000010101101010010111110100100110010110110111100100010100011101010111100000100001100111101001100001010000;
#1 $display("%b", po);
# 1  pi=207'b011010110100010000010000010100101001010111110001111011000011010000101000000100011101011011000011010111001111011001100100000111000101101000001011000000000011010111111001001101111010110100001001011000000011001;
#1 $display("%b", po);
# 1  pi=207'b111101101101000011011001110110001100010000101011100011000000110101010010110101110010101110010011000001100000110000111000101110110000110110101011111011110110100100111100010001001101100101000110001101111110010;
#1 $display("%b", po);
# 1  pi=207'b001001001111010110000111001000111010011001111111001110111011100110110110010111011101011001110111111000001110101110001101101000100100010100101001010110011100110011010001000100101001110010101101110011111111101;
#1 $display("%b", po);
# 1  pi=207'b100100010001011000100110000010000010010100011011011101100110010100101001101111110001110100011011000100100110111010010110101101111000100110000100010111111101000101011110101000110100110110110000101010101111111;
#1 $display("%b", po);
# 1  pi=207'b011010100000011110100000101001110010011001001011001100010010110000111001000010110010111100011111101110110111111111001001101101010001011001011101101111001000010001010101100101101111000100000000010111111101110;
#1 $display("%b", po);
# 1  pi=207'b000100111000011000001101101000001110101010000110011101111001010010110111110100001011000011111101101111001111101101110101001111000010011110101011100101110001010101011110100010110010111011011010000111111011010;
#1 $display("%b", po);
# 1  pi=207'b010100001000110111100110000001011011110000100100100001100011001111000101010101010011011011010001100010100101110010001100110101011001110110010011111011001110000010100001111010110011011000110100100010000111111;
#1 $display("%b", po);
# 1  pi=207'b010101000001111110101001100001111010011000011011100111110111011110101011010101001001100101110011101101011011001111110101100010001111001000000001111101011000000000000110111110010111001100111110100100100011110;
#1 $display("%b", po);
# 1  pi=207'b111011011000000111111111010010001101001001001000110110001101010100011110110001010111110110011011010100101001010010110001110101111110001011001111011011010100000011110011010100010011010010000000011000010100001;
#1 $display("%b", po);
# 1  pi=207'b110001000100010100000010000110100010101111010011111100000000011010111111110000111001001110011001100110100100001111000011000001111000100100000000110010011011011100000101101100001101111010000111011011011010111;
#1 $display("%b", po);
# 1  pi=207'b111111010100011010001011000001110100011011110001100000010011001101010011100000101001111010111010100110001110110100110000000010010001001110001001100100111111100000110011110111100010101010101011111111101110111;
#1 $display("%b", po);
# 1  pi=207'b101001100101101011010010100110000010100001111001011000000101000110000101100101011100000100100001001001100101011110010001000011111101101100000010001011001001001110011110100011111110010111100001111001100100000;
#1 $display("%b", po);
# 1  pi=207'b101100111001100010101000110000011000010100101000111010011110000100110111010000011111111010111100010001001100001010111000001110000000110000111001100001010011000101011000011000100101110110110011111111001110101;
#1 $display("%b", po);
# 1  pi=207'b111111011010010101100000110111101011110010100111111001100011111111010010110111101000000001111110101001101010100000000110100011001011100011000011110000101111111010111000010101000001111101001111111000010100000;
#1 $display("%b", po);
# 1  pi=207'b001111001011011000001000110100110000111001010001100100111101101101110010101001000100011010100010101100000001010100111100011010011000111011001101010111000011110010010011000010110011101011100110010100000110010;
#1 $display("%b", po);
# 1  pi=207'b001101101100000111110011010111110111101111000000101010111100101100001011101001111101010001111001100000010001010011111000100011101110101110110100011101010011010000110111010010100011110111110101100100110011110;
#1 $display("%b", po);
# 1  pi=207'b001001100110100101010010111100000110011100011111001011110010111111000000010100010000110010010000000100000101100000001001101100010001101010001010111100001010110010010001111111000000011000100010011011110111001;
#1 $display("%b", po);
# 1  pi=207'b010011000111001101100111010101100111010101111110110111010100000010101100101011100011101001111001101011101100101110010110011011000001011011110001010010100001111001110101110110001110010000000100101101110000100;
#1 $display("%b", po);
# 1  pi=207'b000100111110010110010110000101100100000111101101010010111001000100011010100010100101100010010000100011100010010100111000100000011010000001101111011111100101101010001000101100001101001001100001110111100111011;
#1 $display("%b", po);
# 1  pi=207'b111001101011111011110001110111110000000110001011000101110011000110001110001111100001000110001101101001100111000011001000001010111111110101101101110001010101101000101110100010001001111111110001011011010011110;
#1 $display("%b", po);
# 1  pi=207'b000110110001111000101101111101111011001111101110000011110000100110100001101110100011001011010101101110001100111101111001001111100000111000001000100011111100010111000100010100111100001110010000100001101100110;
#1 $display("%b", po);
# 1  pi=207'b100101001100011011000100010110010111111100101100001011101101100110011110001111000100011001010110101000001100101111111100100111010110100001001001000010011011111110000001110011111101100011000011110110110110110;
#1 $display("%b", po);
# 1  pi=207'b001101001110111100101110100111101110110011001011111110101100011100010111101110010000010000000100010101101001100011011100011001111010110011101010011100011000110101111001010001101010110111111111111011001010110;
#1 $display("%b", po);
# 1  pi=207'b001011001110100001100111101101101111010011100010110000100100011111010000011011011000101011001100001010011110100011100100111011001001100011000010010000001100000010000110000010010001111011111110000010111000101;
#1 $display("%b", po);
# 1  pi=207'b000010100111101010011010010001000110000001011101110100000000011010111000000000001000111101100101101100111110011010110110101010001101011101010001010001100011010111000001101011101101010011101101101001010000000;
#1 $display("%b", po);
# 1  pi=207'b000111111111000011011110110011000110100101000111100111101001111111001011101011000110001011100101001011100010001010101111010011010000110110100101101000111011000011110000111000100011111000010001001101110010001;
#1 $display("%b", po);
# 1  pi=207'b110010010111101001110100001001010110011001111001010011100000101111010101111100111000101001000111100100111111000010101010101111001010110000000100111010001111110011011001110101111001101001000001101001110110000;
#1 $display("%b", po);
# 1  pi=207'b100111001011001011111101010111101000001000111111010011000001011001001010011011101001010111001001100010000000011010101001110100001101001111001000000100011000010110111000011000000001111000110111100000011101100;
#1 $display("%b", po);
# 1  pi=207'b110111101010100011001101010000010111001111110011001001101100001011100000011110010010011001100101011000011011001101110011100100011100010001010000000110111011100111010111001100011000100001101101011001100011110;
#1 $display("%b", po);
# 1  pi=207'b001100011001000011111001011011011001111100100001001111011010110011011000000010011010010010100001100100010011110110101011010000000110010101011101010110001000100101100010110110011000100100110000010011100001011;
#1 $display("%b", po);
# 1  pi=207'b100110101100001010100001001100100110100101110001000100101010111110011011110001010111110001110110111101001110010010111000110010000110011000101111100110011100010110110111010111001000100101101100001111110011100;
#1 $display("%b", po);
# 1  pi=207'b101010110110001101001000010110111100001001101000100011101100100100110100111001100000101101011000101000001100010100010000100010001010000001001101010011010100110011010011101000001010011111100111111001000101000;
#1 $display("%b", po);
# 1  pi=207'b011101101001101000010010011000111001000011001010000101111110100000001000110100001100110001100110111011010111110110111110101011001111011111001100011111101010001111001110001100001000111000010010101011111010000;
#1 $display("%b", po);
# 1  pi=207'b110000010100101011001001100000011110001101001101000011111001110000001101110101111011110101101100011100001011001110111000110111000001011110110010100101010111100010101001111001010111101011110010011011101100001;
#1 $display("%b", po);
# 1  pi=207'b101001110001010000001000100000000010100000110011100100100000010010110100101010011001010011111011111110111100001111100111110111011101111110010000001100101110100000001010000101010011011011110111010111111101001;
#1 $display("%b", po);
# 1  pi=207'b000000000011011001011011111110001110111000000010001010101011010011100101010101011100001100100111011111101101111110000111010011000101111001101110101101011100010101111111010110101101100010000001110100001111101;
#1 $display("%b", po);
# 1  pi=207'b000110110010011000010111101010000001011000100101011000010010101100111001011000100111111110001101100100111001110100011011010111001100000101101000101111100011110110000001010010011100001010000011001001000011011;
#1 $display("%b", po);
# 1  pi=207'b111100001010011101010101010001001010111110111110100101111101100001110101011001111110101000010110000011001010111010101001010101111101011010000000011001001010110010101101001011101010101001110101000110010000101;
#1 $display("%b", po);
# 1  pi=207'b001100111101110110110001110110000110001110000011010110111001001110101011111101010101101101000101100000101101011001001111111110111111010010000111101011100001000001010101001000111110011000010000001100001101001;
#1 $display("%b", po);
# 1  pi=207'b011000001000000100000011111000100001001100101101100000111010010111001100011001010011011001111010011100001000010100110111000111100011100111110000101111101111100010100111101011110110000111010111010010000001101;
#1 $display("%b", po);
# 1  pi=207'b011011001010111101000011010111011001111111111011100001010101110001111000100100010100000011000100110000100011110011001010110010101011110001000100101001101110100110100010011101111011111000101100101001000010001;
#1 $display("%b", po);
# 1  pi=207'b001000001001110011101110110101010110110011011101011110111000001110100000000100101000001011101000011000111000010001100001000110001010000001000100100011010000011010001110101001010110111011000010000110110000101;
#1 $display("%b", po);
# 1  pi=207'b111111010100110110111011111110100010000010011101100100010011111011110101110010001011011000101000000000111010100011100000110101101110010111010001001000001111001100100111000100101000001000000111100101001100110;
#1 $display("%b", po);
# 1  pi=207'b101011111111101010100000010101010010100111011001111001111000100011010010010101110100001001111010001111010111110010000011000001111101100011100100000101101110011111010000101100001000010111011110110000110111100;
#1 $display("%b", po);
# 1  pi=207'b010001011001000111110001110100000001000111110011001111101100010111010110000101001011111100011010111011101101100101001111011000001100101111001001100100110110000000000110110001001000100000101011011011001001101;
#1 $display("%b", po);
# 1  pi=207'b011001101000111111011011011111001110110000100010101100010000010100000110111100011100110100011100011110000110000110010001001011101110111100010010100111001101100101011000011001100011110000110000101000100110110;
#1 $display("%b", po);
# 1  pi=207'b101100000010101000001001111001101100000011110001111111100000001000110001000111101101010011000100111000101101011110010100010011011000111111100001111000011110011011101110101110110010000110011000000011001111110;
#1 $display("%b", po);
# 1  pi=207'b100111011011010000000010101100110111000100011010000101001000110000001000101100010000001111001010100100101001010101111110001000100010000110111111111100001110011110000100010010000101111000011110010011001111111;
#1 $display("%b", po);
# 1  pi=207'b100001101110110010011111001010100001010111011011110100001100100001100100010111010001001101011101001010000000010000100111101101111100101010010111010110010000010010010110000110110011000111011000101010100010110;
#1 $display("%b", po);
# 1  pi=207'b011100110000110010011110111110111111010101110001111000101100111100100101110010011100111001010000001000011110100010000111110011011100101010001110010001011010100100101101010001010111110100100000010101010001100;
#1 $display("%b", po);
# 1  pi=207'b010010101000001000111010100100110000100111000100000111000011101000001011010111111101000111000010100100100101110110111111000101010000010111110101010111111001000010101010000011110011001100001111100101001100010;
#1 $display("%b", po);
# 1  pi=207'b011001101100011111011100011101111100011111110111101100110110100011101010101111110110000010100010010011101000011011011101010011001110001010001100010100010001100010010101101101011011101000110111100100111110001;
#1 $display("%b", po);
# 1  pi=207'b001000111100101101111000001101011001001010010101000011000100010011101010110011101011011001000000001011101011000010001101100110000000101110000001111001010010010101110111011001011101010011111010110010001100101;
#1 $display("%b", po);
# 1  pi=207'b000011101011010100000100011000100100010011001110010111001010100010100110101010010101001110000001101100111100110101111110001001101101111110011000111000100010110000100111010000001011000101011011111110001101110;
#1 $display("%b", po);
# 1  pi=207'b111010100000110001100110000110100110110100110001000100011011100011010000010100110101000111100110110101011101100111111110101000000110100101001100111110111110110100110100110010001100101100011010011010101110111;
#1 $display("%b", po);
# 1  pi=207'b111001111010010011001000000111010001100100000001000110110111000001110111110110101001111010000011101001110110100111110100000010100100010001100001111110101110010100010111000100111011100001101011001001100000100;
#1 $display("%b", po);
# 1  pi=207'b000100110011000000111000110010111110101011011011001011001010011010011111101001010001010101000110111101110110011111001101011011100111001110000010100010100101111000101101111111101110111011100110111011010011101;
#1 $display("%b", po);
# 1  pi=207'b000010011011011111010000011010011100110000011101101101110101100010101001001010001011111000101111100111101000011010000110001100101101000010101100111101101010111010000110110011111010101000000001011100000010001;
#1 $display("%b", po);
# 1  pi=207'b110100101110001100011101011010101111001001000001101011001010011101001011100010110001111110011101111000011001011110101001100100100010110100000001001000110010010001111000010001001001101001101101101010111101111;
#1 $display("%b", po);
# 1  pi=207'b110010111010101101010011101100100000011100110010100101011011111101011110100001110000111011100101001010010110011110110011110001000011100011110100110011110100100011111000010100000101101111111101111110000011100;
#1 $display("%b", po);
# 1  pi=207'b011010100110101110000110010011010000000110111111011101010111111101010000100001111010100010100110100100110100110001111010000100100001011100111101001011011001011100011000001001001000011101100001000101111010011;
#1 $display("%b", po);
# 1  pi=207'b000000100111101111010101101100001011011010100011010100111000001001001101001010000010101010110000010010111011101000011010101111011000000011110111011100111000101111110111111101110001101110011100101010111111101;
#1 $display("%b", po);
# 1  pi=207'b010111010110000101110011011011000111111110011000111110111110001011101101101001101100000010101110111111100010000101011111100111000100111001100010001101011011101111000111100011010010001001101110111001011110100;
#1 $display("%b", po);
# 1  pi=207'b111011010101100101111011000110001010010101000101010110001111011100010001101111000011110001110011000101000000010001111111010100110101111010101110110001111011100100100000110111101110111010001110011100001001100;
#1 $display("%b", po);
# 1  pi=207'b100101111111110000100100000001011111111110000100101000111111011111000000010111101001010100110101000001001001110110001110111000100111101101010000000101101111000000111100010110011000101000000110010110001010010;
#1 $display("%b", po);
# 1  pi=207'b111000000001010010111010111100101110000110011000011111100100010010011011000100100001011011110111110011011100110000100110001010110110010011000011101111111101010111111110001111110010111011100111110101011010111;
#1 $display("%b", po);
# 1  pi=207'b010011111101000111000111000001111000101001011111010101010011000111010111100110110110111100111111101000011101110101110011001111111000111000110110110011000111100011001101110000110101011100111100001001001111101;
#1 $display("%b", po);
# 1  pi=207'b010011001000001000111101111001111101100011110101111000010000011011100000000011011011110100011001010001101010000110001000010000100100011100010111001100001011010011100001100111001010110001110111001001100011110;
#1 $display("%b", po);
# 1  pi=207'b110000001011110100101011010111111100111110110110110000000100101000100100100100011101010110001000000001010110000111110110001101011001110001000111001101010101011010010100101010001101000000101100101011100000001;
#1 $display("%b", po);
# 1  pi=207'b011000100010010001011011110100000110111101110111111101111101010010111010010110000110000101110101011000011000100100011111100001010100110111101000100011110000011110011010110010111001110011011010001110110011100;
#1 $display("%b", po);
# 1  pi=207'b001001101100100110011011001111001100111001011001001010011010000100100100101010011110000011101010101111011010000001011110110000000101011001011101010011100000111111010011111111101000110001011011011111100010111;
#1 $display("%b", po);
# 1  pi=207'b000101110000100001101101010010010111110011111111101000001011110101100100110100101111101010001000001111010010010101111101111011001001110011010100001000011011101110101010000010000000010001000101100000011000111;
#1 $display("%b", po);
# 1  pi=207'b110100011000100011111000001001011011000000110010001101001001111010101001011111101111000110100000101110101000010111101100011011110110010100000010011111001111010000011001100010011101011001111011010011001001100;
#1 $display("%b", po);
# 1  pi=207'b100001011000101010000000000110100101100001110010110110101011010000111001111010011110000111111100001110101000111101101010110001111111010011111011110001011001111010000100100111101010100000011010011000011001100;
#1 $display("%b", po);
# 1  pi=207'b101111001101000101101100001010000101001001000110110111010010010001110101000001011000111011110010101111110111011000001001100011111011111001011111110110111001011111100010001100101011100110011110110111011000111;
#1 $display("%b", po);
# 1  pi=207'b001011111000010101100111110101010010000101101001111100110000101001101000000101101001110010010111011111001010100001111001111011110101001101000110011000100100110100100111000011110000010010100101100001101100000;
#1 $display("%b", po);
# 1  pi=207'b001100011100111101110110111000011011110000111011001111010101010110111110011100001011101100100100100101010011000110011101000010001010100100111101000101011000000011010100011011111100011000110100111010110100110;
#1 $display("%b", po);
# 1  pi=207'b000011101101011101011111000000011011111001000110011001010001101101110110101101001000111010111000010100000000011100100110110100101110100101100101011001000010111000001010011101100101011101101011111000101000110;
#1 $display("%b", po);
# 1  pi=207'b100001101100000100100010011100100010110000011001100011010000101100100001000100001001011110110111011011110011010000010011000010010001110000101001000100010110000011010111011110000110111011010110101001000000010;
#1 $display("%b", po);
# 1  pi=207'b110100001100110101001011010110000100100100011100000111100000100001000000010000011000010111000110110111000110010100111111011011110011111011111010100001100111010111010110001100111101100001000011000010101110000;
#1 $display("%b", po);
# 1  pi=207'b101111011011101011011011001100011000100010010111010001000010101000011110010111000100110111000110100000100111101100000100111100100000100001001101011100001000000011110101000100101111001101111010111101110000000;
#1 $display("%b", po);
# 1  pi=207'b111000110010101111101000011111010100101011011100101011010001000101011101111010011101010010110001010011010101010101101011011011100010111011010110010101111100000010000101111111100111111100011010000001111011111;
#1 $display("%b", po);
# 1  pi=207'b000011101001111100111001110001111111111110010101101101010001011000100000100001011110111101000101011111001110011011000010111000001111110000001001000001111110110001000101010110001000010111110010111001010011000;
#1 $display("%b", po);
# 1  pi=207'b101111101001001111010101110100011000001100010110111111110111001011100101010110001001001110100001101010111100100110110000011010100011010100101011011101000001001101001111011000001010110010101011000101001010001;
#1 $display("%b", po);
# 1  pi=207'b011000101000100000111101111000001110000100011111011011110111110001111110101111011011101101110100110100100110001110001110011001100001100011010110111100010001100000001101000000100011000010101110001001100001001;
#1 $display("%b", po);
# 1  pi=207'b000010011110110001111100011001111110110010101001110111110010010001100111010010010011001010110001001010011000000010111111000011011110101111100101110110101000011001011111000101101111100101011010111000001010001;
#1 $display("%b", po);
# 1  pi=207'b010011111110111001101011011011110001100000011011101011110101000101001101100010000100001110010110100011110101001001100111110110000001100001110110110111000000001001000100110110101011100111000010000111010111011;
#1 $display("%b", po);
# 1  pi=207'b010101001010001110110101011000000010100111011111110100100101010111111001100101111111110110011000100101001101100110100100100010011001101010100111001000001010101110000000000010111000000100000010111010011110101;
#1 $display("%b", po);
# 1  pi=207'b110001100101101011100100110011110101001011010110110110110010100110000010100101111101011100010110011000101011111001110011000010101110111100111110110001100000100100001101010100111110000011000100000000101100100;
#1 $display("%b", po);
# 1  pi=207'b100110111110111110010000011010000110010101001100100010010000010010101001011010000110110111001111101010110000101000101100110011001111000111110011001011011110101001110001111100001001011011010101110101011000100;
#1 $display("%b", po);
# 1  pi=207'b100011001101101111100101101000110011111111110100000111000000000011000111011000100111011001010011111011101011000111100000110000111110110010010001011000101111011111001100011100111010101111111101110101110011000;
#1 $display("%b", po);
# 1  pi=207'b001101001110001110011000110010101001010111110010001010100100110001010110110011011010010110111101010000010101001101001111111000101000101100111000100001000010010000010100100110110101010101010110000010111000101;
#1 $display("%b", po);
# 1  pi=207'b100100100010111010011000110000000010110101110111111010010101101110010010100111111001111111001100110011101111111111101001011111011010001101100111011111111100000001100000011100001101001011110101010100001010101;
#1 $display("%b", po);
# 1  pi=207'b101111001110100000111001110011010101110111110110111101000000100000111100000101101011001001001000101101110111100100111011001100101001011110011011100110011000001100100110101011000000010100010100000110001111011;
#1 $display("%b", po);
# 1  pi=207'b110001111110110000111111011001011001000010011100101010111110110001001100010000111001110101011001000001011000100100011010010111000011101110101111101101011010011111110100100100000010011111101000010110011011000;
#1 $display("%b", po);
# 1  pi=207'b010010110010001011110010100011011111000001110111100011101000100110000110001010010011011010001000110110111011001010000010011111011011010100010101111001111011110010111111010001101100001101110110010000000000110;
#1 $display("%b", po);
# 1  pi=207'b000010011010100000101110010010111001111010001110010100011001000100111000011000101010000011000011100010100010011010000000000110101011110110110100011011011001100111110001111010111100000011101111101111001111010;
#1 $display("%b", po);
# 1  pi=207'b110110101100111010001011011100000101101101100001110101011101001011001100111100110010000000010110101011010101111000001111101011011010000001101010101010001100110010110011010101011111110001101101011110111101100;
#1 $display("%b", po);
# 1  pi=207'b001101011100001001101000011001011111000010110110101010001101110010011100101111001101001111011100100110111000101110111101011010001000001000000110110011111011101001111001110010011101001000001001101111101110100;
#1 $display("%b", po);
# 1  pi=207'b001111001010100000100001110100110011011100101011110001001010001011101000011110111011110110001100001000000000111101010101111100100101011110101100110001111110101011000101001100111111111011001110001101011000111;
#1 $display("%b", po);
# 1  pi=207'b000110111000111100100000101100000011001000110100001000001111111111110101100101000010110110111010000010101101000011101001100100111110111101110001011001000000101001100010011010100011101100001110111111011111101;
#1 $display("%b", po);
# 1  pi=207'b101100111010000010110111101111101101110000100001110010110101001001110011011011011101110111001110010111101011110110100110011001111010010101101011010111100101010010101001100111100101000100011000011001011011011;
#1 $display("%b", po);
# 1  pi=207'b001110110000001110010101111010000111110101100000100011111110111000000101000100111111010000100100011101000011111100000100100101100001110001110000001110100010111100111111000011000100101101001001001100111111000;
#1 $display("%b", po);
# 1  pi=207'b011011110100001001111011111001100011100101001010110100100011101101001011000101100100110001100011011101100101011010011101100110001000000101011000010100011101001000000111011000001000110101111010100101001000010;
#1 $display("%b", po);
# 1  pi=207'b100011111011011000011110110110110110010100110001010001100010101100010111011111101011001011010101111111000100010010100001100010000001100010000111000100011000101000010100010010010001000001001011100001101001001;
#1 $display("%b", po);
# 1  pi=207'b011111110001001001100111000110101110010100001100011000000100111110100000000011011001101000011111000010010010011111101111011011000101110000000110101111010110100000000001110111011111011010001010001111100001110;
#1 $display("%b", po);
# 1  pi=207'b011001111110011101011110000011101000101110010010100001111111011001001111011011011101000110011100001011101011010100010001010110101110111010011010100110101010100000101111111100010111111111011000010011111010101;
#1 $display("%b", po);
# 1  pi=207'b010100011100100011000101001000111111011000111001010011111110101010100111001100101000111011110000111011101001011100001110111010001001010111110010000110000010011111101000110011100100111011010000100111100100000;
#1 $display("%b", po);
# 1  pi=207'b011110101001011101101000000101001001000011001001010110000111100001001010010100010010111111010111010001001110101010011110110001001001000000010110100010011010111111111000011000001000011010101111001110001001101;
#1 $display("%b", po);
# 1  pi=207'b000001010001001111011111011001110011100111011001010000100100111011010110010011111110110111101100000001100101110100010000000010101100100110100010010010110010010101000001101011101010000001110110100110011111110;
#1 $display("%b", po);
# 1  pi=207'b011010011001111011011101100100000010101001011111011100100011111101010110100011110110110100100111100011110101110100001011110101111011000111011010101000100011100110110100100010110000010010000010100001110111010;
#1 $display("%b", po);
# 1  pi=207'b100011100001100110110101000111010100111010101010001111100001000000101000011111110001010010011000000011100100110010010101001001011010000010011001100100010010001101100011000101110101000011110010100100100011110;
#1 $display("%b", po);
# 1  pi=207'b110000011011011001011001100110101101010110011011001111001011110100010001010000010111111010111100011111001110110001010010011011000001000010010101000001010011100101110011011101111111100011001011111100010000001;
#1 $display("%b", po);
# 1  pi=207'b001010101001101110111101111001000011001001000010101000000100011011001111111011000010011001011101100101011000101100010111011011000111010001000011111100111110100110100001001000110111100001101110100110111101101;
#1 $display("%b", po);
# 1  pi=207'b011001010100110111001101111110100000101000110110110010110110001110111110001101010101000101000100001011110011100010001100011111110000001001011000110111001000000100011111010101001100001001100111010001001111001;
#1 $display("%b", po);
# 1  pi=207'b111011010000100011001101010011001010110111000110010110010001110000101000110111000101011111000000010001101100001011001101110111100111000110111101000011111011110110111000111011000000110101110010111011000101110;
#1 $display("%b", po);
# 1  pi=207'b010001001100101101001000110010011100110011111111100110000111010110100110001100101000101011101111100111100101001011111000000110111010000011110110100001001001001100101000011011110111111100001101001000000001000;
#1 $display("%b", po);
# 1  pi=207'b010100001011000111111101111011111000110001111011010110100000010100000010011101110111110111000000001011010000101011100000101111001001111011011111000101111111011111011110010011001000111011101000000011011001011;
#1 $display("%b", po);
# 1  pi=207'b010110101111010000010111101111011110100010111100101100110100000001000001110010000100111011101011001111100001000011110101111111011111011111011000010010100000101011001000011101011000011001010101110001100001000;
#1 $display("%b", po);
# 1  pi=207'b101110111101111010011100010011110111011001001011100011010000010000000001000011000011011011011100101110101110011100010100001110100101100111110010010111000111000010001110001111111001100000000001011111001001001;
#1 $display("%b", po);
# 1  pi=207'b110101110110101101111000010110001010110111100011100111000011010111010001000000100000100000001111101011001110110001010011011011100110101010100011100101110100101100011101011001101110101001000011110111011110101;
#1 $display("%b", po);
# 1  pi=207'b011011001010000001101101001111110111001101011011000110110110111011111000100101101011011001001011110100001101110010010110101101010100010111001100001101110000100001101101110011011000101100010101001010000001010;
#1 $display("%b", po);
# 1  pi=207'b010111111011101011100101001010111110110110010101000101111000100011100100111011110111111110110001011110101010000101001110110101010001111000001110000111101100110010110011110100011100011001111000101100010010011;
#1 $display("%b", po);
# 1  pi=207'b111100010010110110010101110111111101100010001100000000110011000010110001000100001100110110010010111101000011100111000001011110010111010100001100000110110010101011001001001000011110110110111001101001011110111;
#1 $display("%b", po);
# 1  pi=207'b011000100000011110001110111010110101010011011111110001101110010110010111000000101100010111011110110100100011110101100000101010100011110111100100001000100101110010000110101101101101000001001001110101101111110;
#1 $display("%b", po);
# 1  pi=207'b110010100011000000011010111000001100000101010001100000100000001101011110101010011001100101001001011101110110000001101101101100110100110111110101011100010011100110011010101011010111001110101110001001110101001;
#1 $display("%b", po);
# 1  pi=207'b011110110010100100100011000010101110000110100110001101110001111001110000010001001100101100001000000010111000101101101010000111100101110001011111000001111010111010011101111001001100100100110111011001001010100;
#1 $display("%b", po);
# 1  pi=207'b110011011111110101110111000010100000111101010001001100010001000111111010010100111111011010000000101000010100101001010001100111110110111111000101010001110100101100010101001000101000101110101011001111110111000;
#1 $display("%b", po);
# 1  pi=207'b010101010100001100111001111001010010101010001001011000010011000110101011000100001000110110011010111111101000001100011110010010010001111011011000011101011100010001111100001001011110000011000110111101111010010;
#1 $display("%b", po);
# 1  pi=207'b100100101111111111111100001001001000000011001001001010100101011110000000010101100011000101101011101101100001100011111110001101101001000110001001101010011001101000010000010111100110100111010101111001111001011;
#1 $display("%b", po);
# 1  pi=207'b000010010110100000100000010000010000101110000011110000101101101001011100011000011011111000100100000010000011000010100101100001110101000111100100000101110011100010001100010100001111001100110010010111000001100;
#1 $display("%b", po);
# 1  pi=207'b111111101011111110110101001001010010100001100110000010101000110110011101110110010101100111100110011000011011110011000001001001111010110110000111100101001001001101001110010111101101100010101100000000010000110;
#1 $display("%b", po);
# 1  pi=207'b011100011000010110100001101101101101110011010000010010000110101010100001001001100111101010001110111011000111111010010010001111110111001111010110001000101011110110000110101101100111000111000110001110011111001;
#1 $display("%b", po);
# 1  pi=207'b111111111100010011110011001010000001011110100000111010010100011010001010011000101110111010100001100101110101111001010000010100001000010100011000111010001001000011110000101010111101001011110010101011001111011;
#1 $display("%b", po);
# 1  pi=207'b100001010010101110111100011110000100000110001100100010110100000000011001010111010000010110111000001011011011110101101010100011110010101011010010011001000100010101111111100001010100111011011110100110110011000;
#1 $display("%b", po);
# 1  pi=207'b110101001110110101011101110010100100101100010001111100011011000111100101001100001011000110011011101101011101100101111011100011111100100110110010011010100101110100111000010100001011001101000110001100111100011;
#1 $display("%b", po);
# 1  pi=207'b001000010000100010001100101100010101110001110110011111110101011100010011101001000010100011011110010111101111011011111001010010001011100110001111011111100111101101101100010000101010111010011010100110101101000;
#1 $display("%b", po);
# 1  pi=207'b100011011000100001000000011000100111000010000010011101010100000000111111001000100011110100111001010101100010011010110000111001110011000000011011011001101101000010100000010011000010010110100101001110111111101;
#1 $display("%b", po);
# 1  pi=207'b001001011110110010110110100100001001011000111100111111100001000110110101010001101001010110111101100110000101011001101011111111100100000110011111001110000011000011111011010110111101110100010101100001000100000;
#1 $display("%b", po);
# 1  pi=207'b101011110111001010110001011001100001100100010111001010100110001011011010011111111101111001011001010110000111010110010000111001111011011000110001101110001010111011100100011011111101011110000111110000111010100;
#1 $display("%b", po);
# 1  pi=207'b000100100001101011100110111000000010101000011111110101100001000011110100100111010100100110101111101100010010001110110011110101011100101010001110111001111010111101011100110110010111010100010000110000101011001;
#1 $display("%b", po);
# 1  pi=207'b000101100000111100111001111001111100011110010110100010000110110001001010011001010001010110001001101101110111101001111111100110001111101010001010101011111100100000111011001000011111100100010001000011111011010;
#1 $display("%b", po);
# 1  pi=207'b001001111010001100101111011111100111001001000010100111010101110110100111101011001111101101011110010110101110000001101100111101001100000010100001000101101011100011010111001010100001111010001010010101111001000;
#1 $display("%b", po);
# 1  pi=207'b010111101011001010000000111010101100011100000000111011100110011101111111011010101110000011101010000110000111110110101001101000010011111001000000000101011000101000011001111001000110110000111110000011000011110;
#1 $display("%b", po);
# 1  pi=207'b111000101101011000000010001111110000100010010100111000100000110000000000100111011101000000000011000000010100100001001101100001100100001101111010101101101101000110111011000011001011010001110111001000011100111;
#1 $display("%b", po);
# 1  pi=207'b100010100011101000011110101011110101011111001110111110010011011110010001000011110111111111110110010101110101100010000101100001100001100111010100010100110010110100010111010111000010000110010100001100010111111;
#1 $display("%b", po);
# 1  pi=207'b010011000111001011101111110011101101010010110111001011010110110110111001011010001011000011111111000011110001001101010000110100000101000001110110011101100101011110011100101011111111001011110100100100110111101;
#1 $display("%b", po);
# 1  pi=207'b100100111000111101101000100001011011010100101011111101110000011101010111101000100101101101101001101000100101000110111111001111010001111000001100011111000110001101110010101110100011010101111010111111100001010;
#1 $display("%b", po);
# 1  pi=207'b001111010100010101000110110100001011111010101111010011110000111100101001110011011100110111111101000111010111101000101110100111110100101111101101011010101010110101111011110111001110101111010001010001000101000;
#1 $display("%b", po);
# 1  pi=207'b010001100101100011110100101111110111000110111110001101101010100001110001011000111101011100011010010100100110101011111010010010110110000000011001000111110100001110000011011011111011001010111011101010101100010;
#1 $display("%b", po);
# 1  pi=207'b111011100011110011110010001011111110111001101001001110101100100110101011001010101000011100101011001100010001100100000000011100000110101100111000101100011100101011000000101111001011110100000101110100111101101;
#1 $display("%b", po);
# 1  pi=207'b001010001010011110011101011101010010110100100011010100110101010101000011111001010011100110101100100111011000001010011010110100001011001001001000000111100110000110111001100101110010110010000001000001110001110;
#1 $display("%b", po);
# 1  pi=207'b011100000110101110111010010111010010001001011111111010011100011111001000110101111001101010010000111100111011101101110000001011010101010101100010111010010110110101100010000001101001010100111011011110000111000;
#1 $display("%b", po);
# 1  pi=207'b011001101111001001001110110010001111011011110110001001111000101010000010110010001101110101101011001001011011100011011100110001110110110111010110000111000110110100010100111111100011011011110100010010101111100;
#1 $display("%b", po);
# 1  pi=207'b010101000001000011001111110101111000010110100000011011111001101011001010011010110000101111011001011010011100000001010000110000001110111011010011110100111001010010000001100001110111010010110011001111010010011;
#1 $display("%b", po);
# 1  pi=207'b101110100111101011011001100011001101111011100100100010101111111101011001001100101001010011111000101111001010100011111011110110000000110111011011101110100111010000100011100010011011111000000011011001100011000;
#1 $display("%b", po);
# 1  pi=207'b001001111001110101101110111111000000101100110110101011010011101110111001101100101111110110010101100111100110010001000110111110111110110010101111100111110010100010010110010010000001000001111011011001001111111;
#1 $display("%b", po);
# 1  pi=207'b010101001011010001110110110011100111100110101000100001001010001101101111111010010010110100010110100111000010010101000110001011010001000001010111110110001101110001001111110001011110111111110101110000111101010;
#1 $display("%b", po);
# 1  pi=207'b111010111000101001111000000001100110011011000100100111011011001001000101001000011011010011111011000111100000000010001001001111101001111111001100111000001100001110010110100111000001011101101101001001000100100;
#1 $display("%b", po);
# 1  pi=207'b001000010001001110111001101010110110011111110000001110000011000011110000010001001111101100011001011101100001110000001110101001110001100110110011110000111111010001000001011111011100100101100000010000001100110;
#1 $display("%b", po);
# 1  pi=207'b001110101011010001101100010010011100100111101011011010010001110001001100100111000001001011000000101111100001000000011100111101110011010100001010001101101011000110111010111101011100000010010001001101011000011;
#1 $display("%b", po);
# 1  pi=207'b001010010110101111010001100110000110000100010100011000111010010101111001011110100000001010101111101100000000011000001111110011010110000011100100011010110000101100010110111111101111110111100100101111000010010;
#1 $display("%b", po);
# 1  pi=207'b010010110001011010001110011001101010101001110111000000001010010001101011110011001001001010110100100001001100001110100110111101111101001110011010000011101111001010111111011000110111011100011101011110010010101;
#1 $display("%b", po);
# 1  pi=207'b101010110110001100001010000010000110000100001011010100101011111001110100101011101001101000110001110101101010011001100011111101111111100001000110010110111010101011101000010001011001101101110101100111000010011;
#1 $display("%b", po);
# 1  pi=207'b110101100101001000011101000011001101100011101100001100010011101000100001011000100110101110001001011110111111111110101101101001110101101111011110011111000001110101111110100100000001000011110100100011111011101;
#1 $display("%b", po);
# 1  pi=207'b100011010101100010010010101111010010010001001110101011110100000010001000000010001011100001111001011011101101100110110010000110011110110001111111001000001101110111100001011100101100100000111010011000101000110;
#1 $display("%b", po);
# 1  pi=207'b010101100111010111000001000101010001101101011000101010011110000011001010110100101010110111001111000000000010110110110110110101110000111111000010011010000100010001011000010110010001111010110100011100111101001;
#1 $display("%b", po);
# 1  pi=207'b100001001001000111101011001001001111111010110010110000001001011010110100100010111111010101110001010110101100000110011010011010100110010010101011111001011011010010011010100001111011000010001100100101110101000;
#1 $display("%b", po);
# 1  pi=207'b100111010101101100000110111101100000000110111100000101011100101000001110001011000101001110100111101000011010110101101010110110000100011010001011101010100100011000001101010100001001101011110001010000000111111;
#1 $display("%b", po);
# 1  pi=207'b100001000111100000110001110011110011100110110101011110101100100110011000001000010010100110000011110000111010011001110100100001000011001101101010011011101110111011011111001001011001100111000111011101110111111;
#1 $display("%b", po);
# 1  pi=207'b110110101011101001100100010001111011110001011011111010001100110010111011010010111011011101001000000100100011110111101110000101011110111100010111011010011110111000001011101010111101010110111101101011010100011;
#1 $display("%b", po);
# 1  pi=207'b011110111100011111111011011011110011000111011011101111011000010011101100010111001111100000110010001011010011111001101011111100101110101000100110001001100000101000110000000100010011000101000100010110110110100;
#1 $display("%b", po);
# 1  pi=207'b000011101011101110000110111111100010000011011101100001101000110010000110000010101101001100110010011100100011101110011110010010110001111001111011110001001000011111100100100011110100111111100001100110001110010;
#1 $display("%b", po);
# 1  pi=207'b001011101110000000010100010110100101100111011110111010000011100001011000011110011101100111011110110100110101110100100011111100111010110100001011100010000011010011000010011111101100011110010111010110110000010;
#1 $display("%b", po);
# 1  pi=207'b010011010001100000101010011111110110110001111011011110100001111001001010001110100010110001100111011001000101010100101000101101110111000001111101000000111001011000110011101100001010111000011111110100100110101;
#1 $display("%b", po);
# 1  pi=207'b011000111101110101111101001101110111110011000110000111011000010001111000101010010011110000110000001011101001110100100101110011111110010111110110011010010101111101110101011000010100010101010101101100011100000;
#1 $display("%b", po);
# 1  pi=207'b100100110111010011001011011100011100000001000100011101111110010111110011110110001000100101101111001001101111011011001010000011000001100001001110010100100101110111000110110110100100000001000111000101000111001;
#1 $display("%b", po);
# 1  pi=207'b001101110111001000110111010000111101000110001011011111110000001111111011000111011101001110000101111111001011101110010110101100011000001100100100110001010101101010001111111011101000100001010010101111110101000;
#1 $display("%b", po);
# 1  pi=207'b001011100010001011000001110000000000000001101001001100100111011101101001111111110110001101000011111001101011000110000000000010010111101110110111111110101000001001000110110001010111100110010001100110001101111;
#1 $display("%b", po);
# 1  pi=207'b010111000100010000000101110000001000100000100100101101100011101011111100100111010001100110001101000110011100101001100000110101001101010011001110100110011110001101101000100011111100111011000001100111001001100;
#1 $display("%b", po);
# 1  pi=207'b001010001010101101010111000111111000101110100010101011101000011101010101101001010100101001100010111101101010010010010000100101110000101100001100101011010001000010100101111001011110101010101110010001100001010;
#1 $display("%b", po);
# 1  pi=207'b110000000011000000101000000110000011000001110000001000010100000010011110010100101111000000011000111100001011000110110101110110001110001001001111010100111001101111001111011001010101010111011110100101101011011;
#1 $display("%b", po);
# 1  pi=207'b101110010101011011100100011110111010110101010001101101010000010111001001010000110010001001100111001101010000101100011110101111001100000011101101110001011111101101001111000101011001000010011011101100001111110;
#1 $display("%b", po);
# 1  pi=207'b000110110001011110010000011010001011111011111011110010011000100001110000111100000011010001000000110001100000001011000010101001000011010011000001010100011001011101101111111010100110110101111000010110100100111;
#1 $display("%b", po);
# 1  pi=207'b011001011100110101000000000111101111110110100101000111110110001011011111000111011000111111100110101100001111110000001011001100001010100001000011110100000001010110101101011110010001010001111000101100100110101;
#1 $display("%b", po);
# 1  pi=207'b100001111000100110100111110000001111001111101000100110101000101001010110111011100001001101100010010011000011010111001011100110111001100001111100001001111101010111010110101101101101000101011011011010111111001;
#1 $display("%b", po);
# 1  pi=207'b000100010000110101101111010111001001111100010100011111111011101000001111000011111110001100111001001011101011111001011011010101000011010000101100011011001000000101011011111111110011111100100010000011110101100;
#1 $display("%b", po);
# 1  pi=207'b000101010000101111000110101001001110100111110000001111010001010010001010000110000110001011000101110011001001110001000011001011000001011111100101011111011111100010001100100111111001000010001010010000001100110;
#1 $display("%b", po);
# 1  pi=207'b001101000011100001001001010000001011110011011010000010101111011111000110001101001100011000100001010011111000011110011011000101001111100101101110010111111100000100101100001111101111100010111101001111001010111;
#1 $display("%b", po);
# 1  pi=207'b000101001000011000001010100001000010111000000001011001110001111000011101111111010110000010101111100110100001100100000001110111001010111110100111000001110011000101001001010110001100101111101001100001011000110;
#1 $display("%b", po);
# 1  pi=207'b010100000011100001101110101000000001000110110001100110001011001000101100010110001100001011010110011001000001101001010010101011000100100110001011010110011010100000111101111101010000100110010101000100110111010;
#1 $display("%b", po);
# 1  pi=207'b010110000010111110001111000000100101010011110100001111110100101100110100110101110010111110111101001110010000000110000111000011111010100110111110101111000000111100011100100100011001010011000110110100100000001;
#1 $display("%b", po);
# 1  pi=207'b111000000101001110110010010011100000111101110011011111111111110011111111001101010001011100101011110011001100111010110001100101010111000110011011000011101110011101111010110110001001001010100011011001111000111;
#1 $display("%b", po);
# 1  pi=207'b001010100101110111010010100000111111001011111111100010110100110110101111011011011110010001101010111111010000110001111000001001110110100010110000000111101001010001111111110101101010001110111100010110100010001;
#1 $display("%b", po);
# 1  pi=207'b111101010011110101011000010010101100111010010011100010100011010101000000001111101110101111111101000101000100111100011010101100010001100111111010100110001100110101111010111011010011011111010010001001001110010;
#1 $display("%b", po);
# 1  pi=207'b010001011110001011001111111101101000000100111101001101010000000110011101011101010001010000010100111000000000110111000000001011111100011100100110010001000100101110000011000011000000000111100111001010000011101;
#1 $display("%b", po);
# 1  pi=207'b010011111110110000000111111100011000100000100000101111100000110101101111011010000011010101001010111110010110101110010010110000101011100101000100110001010011011010010100110010100100111110001110000000000000000;
#1 $display("%b", po);
# 1  pi=207'b100111101010110000011001111001100111001100111011010111111000000001000010101110011101001101001101011011001110111010110000000100011101111101001110110000001110110111001011010101111100001010011100010000010010010;
#1 $display("%b", po);
# 1  pi=207'b101000001000000110000011001111111100100011110111001011101101011000010100101111110001101010000001000001001111100011000100110101010110101100001010100111001001011011011111100100100000000101010001001100111100110;
#1 $display("%b", po);
# 1  pi=207'b101111101001001110101110011100011100010111000101101101000110100010011111010111010100001101101110010000101100001101110110101110110100100101011001000100010000101010001101010000011000000111010100101111001010010;
#1 $display("%b", po);
# 1  pi=207'b001101110110000110111100011000101101110000101011101111000001101110100000111110110111010111100010100100111000001111100000100101011010101101001000110000010010001101111100100000101000000110000011100101010001010;
#1 $display("%b", po);
# 1  pi=207'b100110110011011010011000101101101001000100011010111000111001111000010001101101001110110110000101101010110110111110101010011101110100111100110001000100010011001111111101001101110011011001001101011101000111010;
#1 $display("%b", po);
# 1  pi=207'b100010110010000101110101101001110010101111110001110100111011100011000111101110001011110111001000111111000101011100011111010010001000000101010111011001011101011100101110111100010000001011111000100100111101011;
#1 $display("%b", po);
# 1  pi=207'b111010111011101011110110100101101101001010011001010100010110110100001100111000110000110011011011100010000001011010111010111111000010001111110010110001101110110101011000011000101100101111010011000000010010011;
#1 $display("%b", po);
# 1  pi=207'b110011011000010001001110011110011101100000001111100000000011100101000010101101001001001100001101110001111010000011101111011101111001011010110001010000010110111011001111100001110100110000001111110101000010110;
#1 $display("%b", po);
# 1  pi=207'b100000011101000110010000100111011010100111001110001110111010001001000010111010110111101010111111111110000111100100010001000110010000010111100000010001100110101000110101111110110101101111011011111000110001111;
#1 $display("%b", po);
# 1  pi=207'b001011111010111010000111101010101111001000110010010100010100111011001010110001001101100101110010100110111100111011011001011001100001011101100001100110101001111000000111000111010000011011100010010010010000111;
#1 $display("%b", po);
# 1  pi=207'b010111101001000100001001001000101010011100001000011010000111011011111010000010010110011111011001001011111110011011101000011001110101011101010010101110100011101100011101111111001000100100110111011010111001100;
#1 $display("%b", po);
# 1  pi=207'b100111011110100100111010111101111011111110001111111100110101110010010011000110110111100000111101000111001101110110100110010000101000010101101000111001110011000100001000011100110100001001000101100100110101100;
#1 $display("%b", po);
# 1  pi=207'b110111101100010100110110101000000101101100001010101001110111011111100101001010111101101010001011010110011111100011000010111011000110011010101000011000111010111111110010010010000101000100100001111010100001001;
#1 $display("%b", po);
# 1  pi=207'b000100111100100011011000000011011100011101000101011001001010010100011001110011111110010110011111100011011101111010101100110110000111101010111101111000110011000010011101001011000100010011110111010100100011101;
#1 $display("%b", po);
# 1  pi=207'b010001000111011010001110111110110011011001100001000100010101101000001010010011110000111111101100011001111001100011010100101001110010101001111111101000100110101001001101110001000000011100101110110011111101111;
#1 $display("%b", po);
# 1  pi=207'b101100000101101001011101111101000000100100110011010101001100010010000010111011110111110010100101010010001000111000101101001011000010011000110111100111111001000101011001111100110100001111111110010110101001110;
#1 $display("%b", po);
# 1  pi=207'b010001101001110111100110001010001011111101001011110011001100110000111000111101010100001100111010101111111111111111011100001010000111101000010010000111010000111101100011100011100101000001100011100001011111010;
#1 $display("%b", po);
# 1  pi=207'b010011111110101100110011011101001110000011111000111000111101010001000011011110000110001110111000011100110111000010000110110101111111000000010111101001000010011110110000101010010100010110001010010110010100101;
#1 $display("%b", po);
# 1  pi=207'b111100111100010010110001111100101100000010111100000011010010001110000010110001011001010110111010000111010110000011011110111011011110111010011011110101110000001100000111000111111000111010010000010110001011011;
#1 $display("%b", po);
# 1  pi=207'b000101110100000100001110110110011111011110100010000100010001011110101101100011001110011000101001111001001001101010001011011000110111001011001100011000010111100111101111110101000000110110000001000011101000110;
#1 $display("%b", po);
# 1  pi=207'b000001100001101010110100001000100001011101100101100101011111100101101010100001000111100011001110011100010010110100101100000111001001011011001000111110111001110110010101100001111100100000110001000111011100010;
#1 $display("%b", po);
# 1  pi=207'b001011101101111100101111000100010000101000011110000010110100000111000001000110010111000010001111000101001110001010111000110111101000010011001111001010111101100010110011100001011100100100001010000101100100101;
#1 $display("%b", po);
# 1  pi=207'b011100010000011011101110010000010110001101100011011011110011111000001000010100110111111011110110000000101110011000100000110000000001101111110111001010010101010000000110110000000101010000100110011101110101010;
#1 $display("%b", po);
# 1  pi=207'b101010101010011110111010101011010010110001000011010110000010011100111010110011101110101001001001111110001110110111010101001101000011110010100101110111011000010010001111011101111010111110111111001001011010110;
#1 $display("%b", po);
# 1  pi=207'b110000101010110011011111111111001010010010010000101010011101100011000100111110011000001011101011001000100100010010011011000011010000010111110101000101011111011011100010100110011001010010111001000111001011111;
#1 $display("%b", po);
# 1  pi=207'b000100011100111100001100111011000011010000111000101001101101010100110010010100111111001100110001100010011010010101101001101111111101000010010001011011110011110000001001010001100110101100111011101000101011101;
#1 $display("%b", po);
# 1  pi=207'b100111000101001101110110011100011100010101111010000010110100100000000101100100101011011101010111000001110001001110100111010001011101110001011011011011101100010011101100011110110100001001100110110000110001111;
#1 $display("%b", po);
# 1  pi=207'b100111101100010100110011111100000111000000001000011110110001001010010100100110010100100101000010101010010010111000100110101010010010100001010100000111111101000010011000010100110111000110100100011011111111001;
#1 $display("%b", po);
# 1  pi=207'b101010100011010000101001011110001001111110001001100101100001010011110010011101000101011001011000111111101011100110011100101011110100101000111111001000100101111111110111011001101001101000011000111000010110000;
#1 $display("%b", po);
# 1  pi=207'b001101111011011101011001111100011010101101011101001110001000111011111011110100000110111110001100011000100000010001100000010111101000101111110110010110001011010010001011101111010111011101000001101000111100101;
#1 $display("%b", po);
# 1  pi=207'b001000111001110000001011001110011001111000001011110001011111001101001011111000101111000111011010011100010111100001100101010001110011110110111101110100011001110011010110101100111100001000101000011011010000101;
#1 $display("%b", po);
# 1  pi=207'b000001110001110001000000001001001001001000100100110000101111111111010110010000100110010110011001110001000010011011000010100001000011101100101011000110010011011000100011100000001010101111110001110110101101001;
#1 $display("%b", po);
# 1  pi=207'b000010111010000111011000101110101111001111010100110101001110100000100001100001011100001010011101100010111100111000010110100111100000010000000111111111101001010011110100110101010101010101111010001010000100000;
#1 $display("%b", po);
# 1  pi=207'b010101100101100000111111001110000111011000101111111010011100110110010111101100001101110101111010100110111110001000110001110101010001101010001010011010111111011000111101011011101000000110111011100100101000101;
#1 $display("%b", po);
# 1  pi=207'b100100101001001000001110001011010011010001101111101010100000100101100110001101110101100001001010001010010111100110010100011000111110010011010100110110100000010100001010010010011110100100101100010110100111011;
#1 $display("%b", po);
# 1  pi=207'b000011111101110011111001111100111010111010010001100101111000111110000010111011100100101000000110101110001000101101011101101010110101111011000101101000101110101101110110011110001011101011111110000101000100011;
#1 $display("%b", po);
# 1  pi=207'b000000000001101011101100101110000010101100111111100101100110100110110100010001001110111010111110100101110000111010111010100010010101111100101001101001010111011110011101000111000111111111100111110101010100110;
#1 $display("%b", po);
# 1  pi=207'b110000111111101110011110010110101011101100110111000100111111100101000000011000101100001011100001100010101001111010110111110100011011101010110000110111000101001101010111110011011000110011110010011101010011100;
#1 $display("%b", po);
# 1  pi=207'b101001011110001100101111000001011010110000101000110010101110000000101001100001101110100000011111111111100011110101010001100010100010011101001010001111001100001011010000100111100011101110001101111011010100000;
#1 $display("%b", po);
# 1  pi=207'b111101010110111110101110010001011110101001100011110001111001011010100101011000111010011001011111100111110010100110100011010011001010010010100010110000101010000000011010001101110001111010110001100011111001101;
#1 $display("%b", po);
# 1  pi=207'b001000001011101011110101110111011011111011100100011110111101011111110110011111110111011010110000111011100101101110010101111001010100101010111100001101111000110100000100000000111100100010101110001100001110001;
#1 $display("%b", po);
# 1  pi=207'b010111101011100110100100111000010100100011111111011100010100110010000001111010000100011100010011100000111110111101101110001100101000111001000011001010010101011010000111010011101010110101011000010010110010101;
#1 $display("%b", po);
# 1  pi=207'b000011001100111000100100010011000011110001100001011000100011100101110011000110011001000000100011100101000100011100110110111101011010011001000110000110101001111110010111100110110110010001111100110000011101111;
#1 $display("%b", po);
# 1  pi=207'b101010010001111000011110010011111101111100010110100100100111011110100001110001101100100000110100101001101010100010101111100011000100000100001111110100100111101011101000110010000111000100101110111110011010111;
#1 $display("%b", po);
# 1  pi=207'b001111110100000101110010011000001001001001110101010110010100000101001101011100100010011001011010110011011000100110010000000000000010001110100010001110111001000111100111011010010101001111111010100111011111000;
#1 $display("%b", po);
# 1  pi=207'b000011110111111111110101011001011100010111010111110111100101010000101111010001000100111111000111111100100111011000010010011010111110011010000011100000010100110101110100000011111111110100101110001010010010010;
#1 $display("%b", po);
# 1  pi=207'b100110101110110111010110010111011001111000110111110001001000101000011111100111001000000110100000001000011010100001010001000111100001000101000101100110100110001110110110110001000000010100101011010011000110011;
#1 $display("%b", po);
# 1  pi=207'b010101111100000101110000110011110000101111001011101010001010101110000010010011010011001111100111101001110101001000001111101000010011110111100001101001110111000010101100101100001010110000101011001000010110111;
#1 $display("%b", po);
# 1  pi=207'b010001000100011111100100110110110110010110011101000111110101000001110110111011101111001000011001110101111010000101001101010010000110010010111000011000110010011111110111001101100011101011110000010001101001100;
#1 $display("%b", po);
# 1  pi=207'b111110100011011101001001001111011010111100011101101100010100010100101011000010101110011100110010101100011110011010001010100001111010000011010000001001100111011011011001110000011100101110101100110001001100000;
#1 $display("%b", po);
# 1  pi=207'b011100110111000110101101001111110011000010001101010001100110011000111000000000011111011010111101001000111110111111011110000000110010001010100010001101011111000000010111110000010101001010111010100100010011110;
#1 $display("%b", po);
# 1  pi=207'b101001010100101101100001011000011111110001010111000001101100010000001101011111111011110001111000111111011101100111010001000011100011001011011100000011001011000111011110010111100100101100000011111011110010111;
#1 $display("%b", po);
# 1  pi=207'b001011100110010010100110000001100001101110010010011100011011101000011100010111010101000111111000010001000010100000000110001100011100000011000101100111110010101001010110101100000111110010000000000100100100010;
#1 $display("%b", po);
# 1  pi=207'b100110011010101100000000001011110011100110001110111001110111111110011111000001011010011010101111000101111011100101111111010100100011100011011001010000000010110110011110000000011110010110001001000010011110101;
#1 $display("%b", po);
# 1  pi=207'b010110110101100001001111100111110110011001011110000110011110011111100000010110101000100010100001001101010100001010101010000111001001000000011010111010001111100010010101010010100000010011100100111101111110001;
#1 $display("%b", po);
# 1  pi=207'b010000111001000110000000100001101011110011001000010001000111110110101011101101000001000000100001101010100011001100001111000010000010010101001011001111110101010011101001011111110000110001011111111101010011110;
#1 $display("%b", po);
# 1  pi=207'b001110011100100100100001101010010000110101111100110000000011000110011001100100100101000100000000001010111111001001011110001010101111111001111110100011110010001101100101101111111010000010110100011010100011100;
#1 $display("%b", po);
# 1  pi=207'b000100011111011000100100101111011001110110111001001001000000001000110101110110101100110000011100010101111000001101101000101000100000100111001100100001010101101100111111011111101100010000111110010010100011011;
#1 $display("%b", po);
# 1  pi=207'b111100111101011100000101011100111110010100100001011100001000001110010010001000111110110100000001101011011110001111101100101101100001100001011010110101000111001110000101110011011000001110110001010011101001101;
#1 $display("%b", po);
# 1  pi=207'b000010001101011100001011100101100100110111010101101110001011010011110111011001000100010001100000011100001111101011000011111001100100111101011101001011000110000000111010101100111110101100011110011111110111100;
#1 $display("%b", po);
# 1  pi=207'b101101100110000101111101011000101111011111100011001111111011000010010010110101001111001000110110000001000101011110010000011101100100110111001011000101110100101110101101001000000010110011101000110000100001010;
#1 $display("%b", po);
# 1  pi=207'b110001001110011110001100001101110110110000111000101111001110101011110100011110101001001110001100011110011000101110100000001000111000000110001000001111110011011001001001000011010110111101110001100011001011001;
#1 $display("%b", po);
# 1  pi=207'b001101011000001101111101010000010001001100101011111001010011000001110010000111110100001100110010001111011000011100000000000100101100111101000101000101101001100000110110100000011001001101100101011110100110111;
#1 $display("%b", po);
# 1  pi=207'b101011101100001111111111100000110011000101110011100000110000111001111100010100100001010000001101100011100011001010001000100101001101111101010000100000011000100000010011101110100111010011000000101010000100001;
#1 $display("%b", po);
# 1  pi=207'b000111000111101001001011110001111111000011110100100011001010110010110001010100000000000011010110100110001000111010001100001111000000111011111100110110100110010100011101010110010111001001111010101101101010110;
#1 $display("%b", po);
# 1  pi=207'b010111001000101011010000110000000100111100100011011101010110010011001101111000100101101101011111101011101100111101000001110001010000100011011011111111100001011101000000010000010000110110001100111110001000111;
#1 $display("%b", po);
# 1  pi=207'b110011101000010111100001100001000111011101111010001111111111011010111111100011110011000010100011101101000101100110101111000001000110101010011101111101011111010111110000110010010101001000001000011001010000100;
#1 $display("%b", po);
# 1  pi=207'b000100001101111000011111101011101100110011011001101110110110111111100111010000011111111011101101100101011011010010100110010011110100111111101110010011010010011001010000000110011000100010100010101100111001110;
#1 $display("%b", po);
# 1  pi=207'b001110101100101001100111110000000100110100101011111100101100011001101010111100010101000111011011100010010011011011001111110110011110101010110100001110100101001111001100001110010110111101010000001100010011110;
#1 $display("%b", po);
# 1  pi=207'b101100011000011100010110010011101111101101100011100010110001101011100010110011100001011000011001111100110010100011101101100000000111101010111011011111110100010010010011101111011001001101111100001100101000101;
#1 $display("%b", po);
# 1  pi=207'b110101011000011110101000100000001100000011111000011100010001011111101100110101100000101011111001111111011011100010101100110111110000001111110100101111111101011111100010101001000000000110101000101000001010110;
#1 $display("%b", po);
# 1  pi=207'b010111101100110010011100011001100000000111110101011100000010100110010011111011001001110101101011001101001110011111011111100010110111100100010111000100000111110011100101110100110000000011111010110011101100010;
#1 $display("%b", po);
# 1  pi=207'b110010100010101011000000011010011111001110101001111000100101111001101110001011001100011110001101001110001011011000011110001110111010010001100101110010000011000000011101100011100111111011101011111010011000001;
#1 $display("%b", po);
# 1  pi=207'b010111001000011010000010001101010100111001010001001011011000100110101000011101001101000111110001001011101111110100010000000101000011111110110100111011001101110110010100100111011100010101000010101100001101100;
#1 $display("%b", po);
# 1  pi=207'b100011010010100101000111101100101001010101001110001100001001011110110100001000010101110100000100110001000010011100010111001010011111100100111010101010001111101010001011100101110000001001100010111001101010011;
#1 $display("%b", po);
# 1  pi=207'b000100001011011101111111101101001110000000011111101010101110011001100101101110101001001110111101000010100000111000111010011000011101000110000110011110110101110111010101011101111111110110110011001100100010111;
#1 $display("%b", po);
# 1  pi=207'b101000111010000100010111111100011011101111010011110111011110101100010111101110010110101000111011100010110101011110010001111010110111010011110111101010011010010100110110110000000000011110010010101100111010001;
#1 $display("%b", po);
# 1  pi=207'b111100000001011101001010100000010100001101000100000000000010000100011101011010101000100101101111000000110000111001110011001000001011000110010010110001110101000001011101010001100110100110010010000101100001101;
#1 $display("%b", po);
# 1  pi=207'b110000100110111110111001001000100000000101000011111101100101100100011000000001100010001111000100100101001100011001000010100001001010100110000111101100010101111101111101011110001010100001000111101010101111110;
#1 $display("%b", po);
# 1  pi=207'b100000111101000111001100011010100010010000001101001110001111010000011000000111111010010100100010101101110011011111110110111010100010001000101100101100010011011010000100001101100101001010010101011100110101000;
#1 $display("%b", po);
# 1  pi=207'b101000011101100010111100011001110010101010000010110000100100000110111001011000011111001000101010101111111011110101011111000011001001011100000010100011011010101111010000001100100011010111101001101000111011110;
#1 $display("%b", po);
# 1  pi=207'b001001101110100010001000110101000101010000110111011111001011000100011111011111010000101001011010100100000001010100011100001011101010010011000001000011011000101011001110001111001010101000011101001101110110010;
#1 $display("%b", po);
# 1  pi=207'b110110101111101111011111100100011111001011010001010111010011110000000100100010010100011000000101011110000000000111110011111101000001100011010100001111001000000000111110011100100001011000111111001111101110100;
#1 $display("%b", po);
# 1  pi=207'b100111011100001100001101001010111000101110111100110001111100011101110000001011000001011111100011111001000011011010111011101101101111110000101001111010111001111011110100000000011010010010111101101001111010001;
#1 $display("%b", po);
# 1  pi=207'b001101011101010101000010100001010011001100000010100011100011011100110001010101110011110101001111101011111111100101011110001011001001101100111001000000110011101011010011100010010111100110110110111010101110011;
#1 $display("%b", po);
# 1  pi=207'b001101101000100011010010000010000001111101110011111111100001110001010111101110011100101110000000100001011100000111111110010100001011101110101110011011011011100111011010101101000011000111111110001000101111011;
#1 $display("%b", po);
# 1  pi=207'b010010111110110011000010100110001001100101001000010000110110101010101101000111001010110100010110001111011110010010110010111110111010101101000000010011010001101010001111101000111011001010111000100001010101101;
#1 $display("%b", po);
# 1  pi=207'b100111101101100011110001000011101100111011011000111010101010001101011101100001110011111000101000110111100010010000001110010010000001010010010010110101110101110110110101011010011010000111010110111011110101011;
#1 $display("%b", po);
# 1  pi=207'b011111111100011010100011101011001010011101111000001101000011011000111011111111010110001111011011100110001111111101101110111110001101100001101000101111000010101011100001110101001011110101000110101110010000010;
#1 $display("%b", po);
# 1  pi=207'b110000010100001100011100100010010001100101011010101101110000110000011011000001111111100101111101101101000101110100110111011101011000011100111011111110010001110001110111010110111010001110000101011011101001101;
#1 $display("%b", po);
# 1  pi=207'b111111100001111101000100101110000111111101000011110011111111110010010011101100111001100111011010101100100010011101111100001001110000001001010011100011111101000111101010000101101101011001011100011110011101101;
#1 $display("%b", po);
# 1  pi=207'b001111001010001110001001000111011010101011111001010111001110111101011000010010000111100110000110111100100101001100011011111111011100011111111101110001110110100001100100001010010110100100101010110110100101100;
#1 $display("%b", po);
# 1  pi=207'b110001110110010101010111000011100110011000110100101001100000111010001100110110101111101000111101000101001010100110010101011100000100111001111111010100001001011111111010101110110000001000011010001010100100000;
#1 $display("%b", po);
# 1  pi=207'b000000011110010000011001001001101000100101001001100100001100101101010101010001101100011011000010001100011000100010100110001001110000100101011010011100111010011100110110100000011000010000000001111000101110101;
#1 $display("%b", po);
# 1  pi=207'b111110110011000000011001011000010001100000011101000101000100010010010010001101111100011000110111110101111111101110001110010001101101011101110101001011111100101010111000001101011000011010110101010110110100000;
#1 $display("%b", po);
# 1  pi=207'b101000110100011101000111001101110101000110111000100101000110011011010100000111010010010100010101101111111000101011110111111010111001101000101010001100100100000101101111000111101011111101010100101110111010111;
#1 $display("%b", po);
# 1  pi=207'b111110000011110010001100110110000001100111011110000001110100011101110110010001110001110010010101101001100111100110001101010000000101110001100010001100000111000001000000110010011101101010001001111101110101110;
#1 $display("%b", po);
# 1  pi=207'b101110111110100110101100111011100010000011100111100010000010101111100000010110001111101100001001110010001010110110010010101010100100111101100010100111000100001000110110001111000000011010011111011010101011010;
#1 $display("%b", po);
# 1  pi=207'b110010110101000111001100101110100011100111010001101101100010111011101100100101011000001001001101111111010101100111000100010011110001000010110111000000101100010110111000001001100111011100110001110111110111010;
#1 $display("%b", po);
# 1  pi=207'b010100110111110110010010110010001000010000110101100100100001111100000100111010011111000101000001011000101101110011010111110010011011011111000111010010000111100111001101110000010100011000000011110000111111010;
#1 $display("%b", po);
# 1  pi=207'b100000010101111000011100111000001000100010111011010110110000001110110010110001100111111101101101011011111101110110010111100010001111100000000101111010000100101110001101010101101000110111010010001111010010011;
#1 $display("%b", po);
# 1  pi=207'b000000011100000100010101101010010100000111100111100010000110011110000110110010011011100110110110101001010010010011000001101111101110010001011001110100001101110111010100001001111101111100010000001111100110010;
#1 $display("%b", po);
# 1  pi=207'b000101010001010101101100111000001000110101110100100101010111011000101001101000110100001110010011001011000010001110110101011101111011100001010001000111111101111111101010000100100010001110111101000101011000011;
#1 $display("%b", po);
# 1  pi=207'b000110100001110011010011001100000001001010000011010011001000001001011111000110110100110011010011101101000100010100110100010000010110000011011110111011001111100001101110000000001010011000010110100100000000001;
#1 $display("%b", po);
# 1  pi=207'b011101101111000111101111010001001010001011000101001100001010100101011010001001000011110001011101101111001001110100011100010101010110001110111010111000001000011101000011011001010010101110110110100000100100011;
#1 $display("%b", po);
# 1  pi=207'b111001011101110010100011100001111001001000000110111010110110011011110000110101000001101000111001110110111100011100111100101000101001000000100110010010011001001101101101000001001101100001111100110010100100111;
#1 $display("%b", po);
# 1  pi=207'b111110010100001101001100000101010011110101111111100001101000010001110100001001011110100011101111010011100000010011101101101010001010000100010000001010001100001011010110111010010101110001001001011110011011000;
#1 $display("%b", po);
# 1  pi=207'b111101011000100111111010101000001001100111011001000001001111010011010111110110010110110001101011101000000101010100110111001110010011001011001001101110111001010110100110100001100000101010010000101110100001011;
#1 $display("%b", po);
# 1  pi=207'b000000110110000110110011100100000000001000101111000000100100000111001001011110000010110111011100000100110010011010000111101101110000101000100010101100000110000011011101111011000110010001001100110111100111110;
#1 $display("%b", po);
# 1  pi=207'b111111010001000101010000001111100100100001001001101100010011110011100010111101110101001101100101010000010110101010010000011110101010010010100010011101110100111011001110011011001110011110011001101011100011010;
#1 $display("%b", po);
# 1  pi=207'b011010101100010010111100110110010001011001010111011010001010011010001101001100001000111000011111011111111011110011110111110010101000011001000110010110101101100110101110011011111010111010110011011101001000010;
#1 $display("%b", po);
# 1  pi=207'b000101001000000111011000110000110000101011101011000011100010010000000101000001000010110011001100001101111110000111100110110010011011101010000110011101101011010000100111010001010110000000111111100111110011100;
#1 $display("%b", po);
# 1  pi=207'b001000011101101110100001111010100011100101100101010010001111010111011100010000001100011100101010000101110100011111110100000010011111001111001110011011110010001010010010001110000110110011000001011100100000110;
#1 $display("%b", po);
# 1  pi=207'b010001100001011111000111110011101111100111010000110101101101111110100101001001111010101010010001001111100101000001011001000101110001001010100000101100111011101000101000101111100111110101010110111010011001100;
#1 $display("%b", po);
# 1  pi=207'b110101010111011111111110101110011100001100011110011100101101001011110001000111000110001110001010010001010111000011001110110001110100110110010010100111110101001000001111101110110100001011010100110001001010001;
#1 $display("%b", po);
# 1  pi=207'b110010110100001010110001100111101000100110000000111101101000001110001010011110101000101001110111111101100100000100000010111111111000110010001001111111011000111101111100100111101101001111111000000110101000111;
#1 $display("%b", po);
# 1  pi=207'b000010010101001011010110100110100101101000110000001010100111100101110110001100101000111110110100001110010000110011110010111000100111010010010001101011011001010101101111101000100001001001110101010000011100111;
#1 $display("%b", po);
# 1  pi=207'b111000100010011000000111000110010100011011010010101011010010100011001100000110001101111110001011010111111000010001110011001100001000100011001000110101010100000101110100011101000101111111110001000011010010001;
#1 $display("%b", po);
# 1  pi=207'b010000111000110011100101101011011011111001100010011110000000010101001010000000101011011000101011100010110011111111010001000111010000010010011011011001100110111000110100001101100000000001110101000110100011110;
#1 $display("%b", po);
# 1  pi=207'b111001011000011110110101111001110010101011011001101100010111100100000100001010110111000011011000001000111000101100110000011100111111110111001101110101110110111001001111111100101101100011110100111010100000000;
#1 $display("%b", po);
# 1  pi=207'b011001010001011010001000110000100110100000100011010011000100000010110000110000100110011101100010100010100101001000101111110110010101011011001001011010101110000011001011000011011001000010011111010010100001001;
#1 $display("%b", po);
# 1  pi=207'b110110111011111110111110010101010110100111110010100011100110000010110110001000001110001001111010111000000001101011010010101100101001000010000000010001001011110110010100111110010011111010001101001001110101011;
#1 $display("%b", po);
# 1  pi=207'b100110101000011111000101001111110111000010001011011010100000010101101100100010111110001111101101101100000101111000101110110110000010010100101000001100010101001010011011010100110000010001111100000011101110100;
#1 $display("%b", po);
# 1  pi=207'b111110001101100010010001011001100000100111100100010111111011100010010000111001011000001011111001000100111001001110110100111011101010011000101010011001101010011111010101100010101111111110011001110100011100110;
#1 $display("%b", po);
# 1  pi=207'b000111101101010111010010011010101000000110100000010011101011111111000110110111111010110111010101011111010011010011110100001000010111001100001011001000001001110001010001111001100001011011101111001111100110010;
#1 $display("%b", po);
# 1  pi=207'b100010000000011000001011110001001111101010100011001011011010000011110110101101101000001110110101010100111110101100101010100001001101110010010000111011010010101000011101011001000111011100011110010110101111100;
#1 $display("%b", po);
# 1  pi=207'b101001110001111110010110001011010110100011001000001101000011111101000000101010010000100011101111100100011010110110000111010101011011010111010101000011011000110101100000100010011111100101000101111110110110010;
#1 $display("%b", po);
# 1  pi=207'b111111101110100100001001011000001110111110100110010100111110100100011101101010100000100001111101010100111001001110010011011001011011110010000111110111111111010001000100010111000101001111101101101101110010001;
#1 $display("%b", po);
# 1  pi=207'b000100011011100000111101110001000011000111001001101001111110010001010001011101001000100111100010101011111100100010011101010110011101100000001111100001010010111010010101011010010010010110110011110010111001001;
#1 $display("%b", po);
# 1  pi=207'b001000111011111111111000000000101110011101101100010110100101011010001000101010010001010110100110001101110101101000001110111011001010100010110010000001011010000011001100010011110010000111010101010010010111001;
#1 $display("%b", po);
# 1  pi=207'b111110011110001110100110100010001001000100111110101011010010011011010011111101000001101111100111000110101011111111011110001101100000000111001000011100101000001001001100100111010100011011100010110000001101000;
#1 $display("%b", po);
# 1  pi=207'b111001111101000101000101001010100010010111010110010110000010110011101100100101000010101100000111110101010010001111001011111001011101111100000101101010100001000011110100000111010001100000110110101011011001010;
#1 $display("%b", po);
# 1  pi=207'b100000001110101100110101111000101111010001001011110001100110000111011110000000110001111011011111001001010010010101111110110110101111010110110011101000101110000011011010000100010000101000101000011111110110101;
#1 $display("%b", po);
# 1  pi=207'b100000101101001001000000111000111100001101001110011010010100000110011001010110110010011101110100001010100011000100110011001101001001010101011000010110111100011100101001010010101010111101000101110101010101111;
#1 $display("%b", po);
# 1  pi=207'b111010101001010101100110000010000100010101000111001000111000001101001001111010100001100111100111000110110000001101110100011000100111000000110101001111100011111011111011001010011101110101111111110100111100000;
#1 $display("%b", po);
# 1  pi=207'b000010100001010110010100110001101010100010011101100111100001100110110001101110000010110111000111001111111000101111111011011100101111010111001001111111001001001000010000111111111101011001000000110100000000111;
#1 $display("%b", po);
# 1  pi=207'b001101011100010111111110100011001110111101011010111011110111001101010000001101000000001101110001100010101000110100100111011111101101001111000001100001000001110010100001101011110100000101101101101001001001110;
#1 $display("%b", po);
# 1  pi=207'b011011100001010011101111001000111100000101010100111100110101111000111000011101011000001100010101100010100110100110010000001101001110100000110101111011111011011111000000010111111110010100010000010010110111101;
#1 $display("%b", po);
# 1  pi=207'b111100011000101111101110001010110111010000101101100010100110111010000110100110111000101110011111010001111111000001100011010001010010110000001001010100011011111110001111001110010101010101111110001111000100010;
#1 $display("%b", po);
# 1  pi=207'b001000100100011101110110110011000000100001101110100101001000111100100110011100011110110011001000110011010001101100001100100010111010010110101101000101101010110010111001100110111111000111101001110101000010001;
#1 $display("%b", po);
# 1  pi=207'b100110111010110101100011000000010000110101011010000010111100101011101000000000001101011011111110101111110111110110001011011001101010011100000101011010111011100000110101000010110000100000101111001001000010110;
#1 $display("%b", po);
# 1  pi=207'b110010000010101111000010111000110011010101001110000111001111101110000111101001000101011010010010010001100101110000100010101101101110110100111111010110000100011011000110110000110011000110101000100101111001011;
#1 $display("%b", po);
# 1  pi=207'b101110000110110001111100011001011110101011101010100000000010010101101001100110001010111011110011100011100111001001111100010110100010100101110011011110000001101110010101001011111010010111100000000001110100011;
#1 $display("%b", po);
# 1  pi=207'b100001001010010000000001001110001100000111000101011001001011000100101101100100011101100010111101000100101101100001101100011011001101100011001001011110111001001100010100110110011101111000001000101111000001111;
#1 $display("%b", po);
# 1  pi=207'b000101010110000110011111110100011010101100001101111001111100011101000101000100011100100111000110100010111010111101000100110110000001000100000000101001000011101101110100110110010110011000011110101111101111001;
#1 $display("%b", po);
# 1  pi=207'b011101101101111110110010110111110010100010000111000110101101111000111011001101110011010100010111000100100010001011100100101011001100101001001001011110101011101111000001011010100011100000000110000011111110100;
#1 $display("%b", po);
# 1  pi=207'b011010100011011100110000010010101011111011110000110111100010001011010101001110110101011000110101011010000100011001011011110011011011001101010011011110111110011011011011100000001111111111010101111001110001011;
#1 $display("%b", po);
# 1  pi=207'b110000101010101100001100001001011000000000110011101101001001110101001110001111000110010100100001000100101101000011010011011011000000110000011001011000100110110100011010010111011100010011011101010010101101110;
#1 $display("%b", po);
# 1  pi=207'b001011101000110100111001001110101011011100011110001110001111111010100101101000101001111100001011110110011011001110011111011100001010110101011010000010001000110010000111000110001110011111010100011111100101110;
#1 $display("%b", po);
# 1  pi=207'b110010001001001101100011111100000001010101011111101101011111100001001000100101000111001110010110101100110001000111001111001111000111010000000001000011100110011010110101110001001100110010001000000111100100111;
#1 $display("%b", po);
# 1  pi=207'b100111101101010100000111111110001001001111011110000010001101000111000010100010110011100000100110111111110110000010011010011111101010110000000101010011100101110011100111000010000000011110110010010000011011010;
#1 $display("%b", po);
# 1  pi=207'b111010111000100100110001110111000110110111010111110000001000010001100111110010101101010011100110111111111010110000110001000100000110000001010000111010101111110000001111111000111110000101011001100101111101110;
#1 $display("%b", po);
# 1  pi=207'b100101010101111110110101010000001010011001101010011011100001110001111011010111101110100101001101110101100001110001000110011011001110011111111110100100000100100010000111010011010011111101111111011001100010110;
#1 $display("%b", po);
# 1  pi=207'b111011010011110100011001000000100010100010011001011001011001110111110000011110001110110011111100011100011110000100100011010101011101110011001001010111011010011001000000111111110000110100001100000111111100111;
#1 $display("%b", po);
# 1  pi=207'b000101110001111110001000011011011101100101111100000001101100110001011100001001101010001110000010011100000000011010110110010110111111110101110111101001000111011111010010001101000001110010111110010111111101100;
#1 $display("%b", po);
# 1  pi=207'b000010101001101011111110000111011011011111101111100000001110011010100101100011101101010110001111110000100111000010111101000101101100110000101000010110100111000101101000110011111111100111001100000010101001100;
#1 $display("%b", po);
# 1  pi=207'b111111011101011111100010010100001111110011000000011010111010110110011100110011000010101010011000111000100011100011100001011000010001000000000110001000010110111100011000001111011000110101011101101100010001101;
#1 $display("%b", po);
# 1  pi=207'b000011100101110101001011110001010110100101111011000100100101100110000000101000000101001100101011010101011110010110110100110110011110011111010001101100100110111101001111111111100010110101100100101101111101000;
#1 $display("%b", po);
# 1  pi=207'b000011110010100011110111100000101010001011100010111110001101011010101011110011110010001101011000011110010110001001100001101111101001101101110101010001010011110011110011111110010100101001001011111101110010111;
#1 $display("%b", po);
# 1  pi=207'b000001111010010111000100001001100110111100100100001110110010010011001011000010010110011011111010110100110011011000110000100000110101111000111111011000101001000011101011110001000110101111100111111111110010011;
#1 $display("%b", po);
# 1  pi=207'b101111001111111110000101101100111010010101011111011000000001001010100001010010101001000000000000010010110010010011000010101010010001011011111000101110110011010011111000101010111101000110110011100110110110100;
#1 $display("%b", po);
# 1  pi=207'b101100111011110011010100111101101010010001010010010110001001011100110000001011111111011110000100010001010011010101000001010000101100111110011100111101001000011010011101000111010110010110011011110111000101100;
#1 $display("%b", po);
# 1  pi=207'b110101010100000000101110011110000011001010100001101000101100110010000010100010011111010010000011110101011101110010011011111101101010011000000001001101100001010110011000110111011111000001011001001101110010110;
#1 $display("%b", po);
# 1  pi=207'b101111100100001011101101000010001000001111111011010100101100110010010111101100110101101011010001010010110011001101001110001001010001111001011100101000011010101101100100001010000110111001111100001011101001101;
#1 $display("%b", po);
# 1  pi=207'b101101111010101001001011100110011101011101010110111011101111010111110111010101011101111001000000110001011101011110010001010000011100111001101001111011010100010010010010000010001010011001011010101111010001101;
#1 $display("%b", po);
# 1  pi=207'b000001110011101100100011000010001000111101110011101010110100101101111101001000011011100111001000101000000110101010000011111000101110101110001001000111100000011101011110110101101110110111010100101001010011000;
#1 $display("%b", po);
# 1  pi=207'b011011111000000101110011011111100111110111001100000011111010000001000001101100010101001000001000101010111000100001000001010110010001110110111100110100101010100110101101110110011100001110101010001001001100111;
#1 $display("%b", po);
# 1  pi=207'b001101010111111001010110010100000011100001100001011000101100010111001101111101011111100110000001011000111000001111001010111000101000110010111011100011100001111110001000111010101111010100010100100100111100011;
#1 $display("%b", po);
# 1  pi=207'b010111011010001010001101010101101110111111101111001011101110111111011000001001000110011001100010110101001001010100101001001011001010000101101010011110011101100100111111101010010001111000111010100001110011101;
#1 $display("%b", po);
# 1  pi=207'b001000000110101000100100010000010001110100100100010111000110011101000111000011011101111110101100011000111100011101110101001000100110111100001100011111111010001110010001000001000111011001000110100111000111111;
#1 $display("%b", po);
# 1  pi=207'b101100011111100101111001010000000001101011100010110011000000011110111010101011100000010111100000001010110000010111001101101000001111000100100101101110011100101000101101001000010111011110000111111100101000101;
#1 $display("%b", po);
# 1  pi=207'b110010110110101100010101001011100010111001001011101111100001001010001110000011001100011010111000111100011000001101100011110011011110001000111110111001110000110000011010001101100100011000111110011101101011000;
#1 $display("%b", po);
# 1  pi=207'b101000100010111110100100111101011101001001001010101100101100011100010011001011010110001000000011010100000001001000100111100101000001010000000110111011001111011000010101011101101010110111100100100001101011101;
#1 $display("%b", po);
# 1  pi=207'b100010110010010100110110011001000111100101111010011001001101111100110000011110010111100000100100111000011000001000111001001110000110110011100001101011000000001100001100110011110011001111110010110001010100010;
#1 $display("%b", po);
# 1  pi=207'b010111111011110010101011010101000100001100011111101110000100111011110101001110110001011011011001101101100000111111111001001110001110101100101100110111111110100101011001101011001110100010111011101010001110000;
#1 $display("%b", po);
# 1  pi=207'b000101100001010000110100110000001010000100110001110101111100001010011110111100101010001001110011010110000101101010000111111010100101110110010101001010010011010110101110111100010011101001010010011101101100011;
#1 $display("%b", po);
# 1  pi=207'b001101101010011011101100100100001101000011010001010101011100011101001001100001010010000001111000001111001011111001100011110100011001011101000111110101110101100000110101111100101001111110110011011101100011000;
#1 $display("%b", po);
# 1  pi=207'b110110111010101111010010101100011000111001110000011010101111110001001010011001011110010000011110000001010010110000001011010000110011111000000100111001010101100100011001100100101110100110011001001110011010110;
#1 $display("%b", po);
# 1  pi=207'b110010100100000010010011011000001100110111100010011011001100110110100000110010101100111100100010001110111010100010001100111011100011111101110110001011011010011010111111110110110101111011010011100000110100110;
#1 $display("%b", po);
# 1  pi=207'b100100011111011110000101010010011101110101100001110101010111001100110000101101001100110010011100000011101001000110101110011001111001101110100010010001111101001101010010110111101101001000110110101111000001110;
#1 $display("%b", po);
# 1  pi=207'b011010110000011010100000100010000110000000110001001000000100100111100100111100110100000111000100111000110000100100010110001110101111101110110001100101111011000100010101100011010101001000110010000001111101011;
#1 $display("%b", po);
# 1  pi=207'b111010011111001101110000000000111001010101101101010001011100011111111010000111001101100111101111110010101101110111010000011101010000101110010010100111101000011001111011110110110101111000000101000101110100111;
#1 $display("%b", po);
# 1  pi=207'b111110111010011010010010010001010110011101111111000000010011101011001111001110000000001010010010010100010010110001100010101111010111110010111101000101101011010111111000110101011110111001011010111100111001100;
#1 $display("%b", po);
# 1  pi=207'b000011000011001001011110100010100101100111100000010011011010101100010011101111001100000101011010111110110100110000011011010101000111011111010101001000101100010101001000000101110100110011111111101111010011100;
#1 $display("%b", po);
# 1  pi=207'b000010110101110010110010101110101101000111001110001001101111000101011000110110110011011111100001100111001100001111001001110110100101000111000011001000010010110110001011101000010000011101011000101010110111110;
#1 $display("%b", po);
# 1  pi=207'b101000100001100101100100111110101111110101101100011101011110111101111110100000100111000000011000100010000111100001100010101111001101001101110101011100001011011110110010000000110011000100011010000000010001101;
#1 $display("%b", po);
# 1  pi=207'b001000010011001000010011100000110011011101010010000001111001101110111001101000000000000001011011000010010100111100100100010110011101001101011110110011001100110001100010100110010101101111100100011000001100101;
#1 $display("%b", po);
# 1  pi=207'b011110010010011111010001010101110100001010010110000100111100110101011111011001001010011001000111100100011110111101110110000000000111000110110100100011011110001111110100011001000000101110010100011101001010111;
#1 $display("%b", po);
# 1  pi=207'b010111011000111100000101110001110001110000110110011010111010100010001110100110111101001100001110000100001110111110001001100110000110111111000101100010111001010000111110110101010011101010101000110001110010000;
#1 $display("%b", po);
# 1  pi=207'b011101010001101110110010001001011110111001010001010111101111000011111010101111011011101011000100000111011111110100011111001011110100101001100000110101100000110010110000010001111000111000100011010110011010100;
#1 $display("%b", po);
# 1  pi=207'b110100110110110010001000001001100101100001100100010111000111001000011010010101101100110000100111111111000111111100011000110001100111100111100100101010010001011101100001110111001100100001000000111100011111100;
#1 $display("%b", po);
# 1  pi=207'b010100001111011110000001110010110000000000001011101100011011010010000110111011001001100101101001001110000011111000111001101100000000000100011110000110011011110101111000011110011111111100010111110011010110110;
#1 $display("%b", po);
# 1  pi=207'b010010101111000111001011001001110110001101110100011101100011101011100110000001100000111110101100000101100011111000001111100001000111010010101000110101101100100111110100111010001100001100000011001110010110101;
#1 $display("%b", po);
# 1  pi=207'b110111000010000100100111000001110001110011001100101001101001000000011010000001100001000001000000010010100001110010101011111101010001011110000111100110111010010110001001101011101101000111001000110001010000111;
#1 $display("%b", po);
# 1  pi=207'b000111011010001101001000100011100000000111001110110000101111110111110010100100000000000010101000010111110111110010110000110101100100101010010100101010111110000010111011101101100101110001010011101001110001101;
#1 $display("%b", po);
# 1  pi=207'b000100100111001010010000101100110111111110000100011010001110010101010101110110110110011011111110101000110001011100001001000101101110010111001001100111110000000111110111111101011000001110000110101110000011000;
#1 $display("%b", po);
# 1  pi=207'b000001011000000011010000101000111100001110000100000110001111111011110110101101010001101010000000100011011110100011000110110101000100011101100010100001001000001001101101101111011100110101110111001001100110111;
#1 $display("%b", po);
# 1  pi=207'b001001010110111000010101100011000010100011111111010101011001001100100011001111001100011011000111101101010100101111001110101101001111100010010101010101000111010101101101000000001111010111000011100000111010111;
#1 $display("%b", po);
# 1  pi=207'b000110001100000001101001001101011100011110110000101000100101111110001011111101000100001111011100110000000001010001110100110111011010110011110101001010000001101100101001111000110011011100101110011011100001000;
#1 $display("%b", po);
# 1  pi=207'b100000100101111011111000001110101111000111011111110100010001000111110010111011101100011011010001011111011011001111000010110001100111111010111101000011011111100101110000101010011100010001111111111111111001101;
#1 $display("%b", po);
# 1  pi=207'b111000101011000100011010111101010010111100000110110101001010111000010011101111011111100010000001100101001110100100111101011001001110011101000000001011001000110111110010011011110111111001001010111110111011011;
#1 $display("%b", po);
# 1  pi=207'b111101011000110001001000010001001000001111111010000011000011110001110001000100000001011011101110011010100100111110111010110000100010100010010101111011111000001111010111011110000111001000100101100100000100011;
#1 $display("%b", po);
# 1  pi=207'b001110100011011000111010011100001010111100111001001101011110001000101101111110001111010001010111010000111011110011110000011010100000000110011111101101000100011100101110111111110000101000101011110100010011011;
#1 $display("%b", po);
# 1  pi=207'b100100100110111110001010011110101111100001110000010110111110110001001010100111101011001000001010100110011011111111000001111001001010001010100011010100100101001110010101010100100111010110010011111101111110001;
#1 $display("%b", po);
# 1  pi=207'b100100010010010010001111010100001100010010001011000111001111000010011110111001011011000110111101000000100100001011110101001000101111011010010100101110010010000101011011001001101111111010001000010000100010100;
#1 $display("%b", po);
# 1  pi=207'b110011000100000011111111001111100110010010101001100000010010110011011000000100101111101001001011110001100111101111110111110101101101101011000100000110111100000111111110100001010001111001100100111001110110000;
#1 $display("%b", po);
# 1  pi=207'b111101111110010011011100100010010100101001100100110100001011101101100100111011110001111010011110000111010000010100000100110011110110100100101010001011011111101001000101011000111000101000110000110110000111110;
#1 $display("%b", po);
# 1  pi=207'b000000011101110110000111100100100011010101010110011100101010101101010001100111101000111001110011010101011001101001101010000001111010011010110010100011010100111000001011101011100101011100001000001010100110111;
#1 $display("%b", po);
# 1  pi=207'b010100110011101111000100100010010010100101110100010010001101000011110011011010011001000001011101011001010111000010111011101101101101110011110011100000010011101110101010010100101011100000100110100111100000011;
#1 $display("%b", po);
# 1  pi=207'b011101001011000010011001111001011011001001110100010100111101111010111111100101110100001011010000011010111000000110011000011000011100000110011110101010111011100001100010110000010001001110110111010011011111100;
#1 $display("%b", po);
# 1  pi=207'b110101001011110010111001111101111100110000011011001010111001001001010010001101110101010101101011011111000001000101000010001110000000011001111111111001100001100101111011101100111101010100111000100101000011011;
#1 $display("%b", po);
# 1  pi=207'b010111001110011110010101100001101010100011011001110010010101101110101111000100001101101111110110101000001001011101011000111000001011111000100011111101111101111001111111111010000110001010110000011000000011101;
#1 $display("%b", po);
# 1  pi=207'b010010101011101011111111000100010011110001000110001010010100001001001010011010001001001111011110011100100001110110010001100000101010000010010001010011001001111110010000101010101111111100100110100100111100100;
#1 $display("%b", po);
# 1  pi=207'b011001001100001110110100110011111110000001100100000101001010110101111001010110101101001101101111010001010110001100010100010110011100110000010110001011110100000011101001110110010100101110001010010001000001000;
#1 $display("%b", po);
# 1  pi=207'b001100101110101101001011100110000101101111010110001110100100110011101000111100000011100001000010111111001111110000000010011001011000110000100101110011011010001110100100010000010110100000100111100010000001010;
#1 $display("%b", po);
# 1  pi=207'b010001100101100010010101100100001011111100001011010000011100001110011011100010111111110100110100011011110100000010100101100111111100100001101011010001000111111011111000100000010100000000010000101011101010110;
#1 $display("%b", po);
# 1  pi=207'b010111000111111100001011101100111000011000001101100100100111100110010011100111101010010100111011111001010101000010010010011101001011011100000000111100000110111011001001000001111011010000001101100100101101011;
#1 $display("%b", po);
# 1  pi=207'b010010011000010101100101110110001000110100000101001010010010110001110101000000110111111110101000110101001110111110010011011011011101111011010110100101011000100011010110101001011001001110010100001001010011011;
#1 $display("%b", po);
# 1  pi=207'b111110000001011100000011100110010101111111011001010001011010011000101001010100000010001101110010001001000101010110001001101111100000010000100000001100011001110000011101100110001100011001010100101110101011100;
#1 $display("%b", po);
# 1  pi=207'b110101010010101000100111111001011001011010111100011001010100000101101100100010101111100110010011101111110010110001001110011110000101110101011101110100101001001011001111011101110010111001001010100001111000100;
#1 $display("%b", po);
# 1  pi=207'b101111101011011000100100010000001100011100010011000100001000011100001101101011100110011011111111000001011000101110111001001011110111001100100100011001100100011111100101000110101001110110001101110011011100110;
#1 $display("%b", po);
# 1  pi=207'b000011111001100101011111110101110110011111100011110100101000000111000100000101001101010100101111001000100111001111100110100100001111000011001010001101001000111100100111101100100111110100000101010010010010100;
#1 $display("%b", po);
# 1  pi=207'b110011001100001001001110010101111011010010101010111100000111011111010010110001001010000101010010011010100100101100011101111111000010100100001110110100101100111011010011111100001011101110010000100001001001100;
#1 $display("%b", po);
# 1  pi=207'b001000011101110101111110101100101011011100111001111100001101000010111101101101101111001110100000001010100100110000100111111001010101101010001010100001000001101111111111000001110111111110110111000001000110000;
#1 $display("%b", po);
# 1  pi=207'b011011011000110010010110100010011101110010000001010000101100001011011100100110001110101011101011100111010111000111010011111000010110000101010001100010101110010010110110010100110100110100110001000011000110010;
#1 $display("%b", po);
# 1  pi=207'b000111000011010101011110001010010100100011011011101011010001100110011110111100011110010011001101110110011010010010110111001010010011001010110110011001001110111000110110011101011001001000111010101011001111100;
#1 $display("%b", po);
# 1  pi=207'b011011011111000110111000001011111001000110100001100100100011001001011010110101100000111010010000001000000110010010111010100101110010001000110000001010010111110111011011101000000011111110010111110100010101000;
#1 $display("%b", po);
# 1  pi=207'b100110011110110101001000000010000000001000001111110000001001101110000111001100001010010111010111001101001011100010110100011010011100011111110001110101101110111110011000111110100001110110110001101000000010110;
#1 $display("%b", po);
# 1  pi=207'b000110111101100100101111110010100001000001000010000100111011000001100000110111011000011100010001000011001111000011000000111100110000110000001100100111101101101011101110001111101011001101011011101011000111000;
#1 $display("%b", po);
# 1  pi=207'b010100111001011100011100010111010000111001100010110100110111011010001001110101010010111000000010010000101011110101001111000100100011001100010000001001101001010001100111101001001110101001000010001110011010111;
#1 $display("%b", po);
# 1  pi=207'b010111000110011010110110011011100110111001001001001100011100011011000011011000111010101011010000011110100010001110000110110001000000101110011111010110001111010111100110101000101001011100100110000000010011101;
#1 $display("%b", po);
# 1  pi=207'b001000000001111011001100101000110111010000100010000110111011101011011010011110101010100101000111111110011010101010100001111010000111011101000001110010000011111101100010110100110010101100100110001100111011000;
#1 $display("%b", po);
# 1  pi=207'b100101101000010010100110101111011010001001100000010011110001000011000001001011000110101000111001111011111111010111010010001001011100001010010100011110001010011100001001011101010101010100110101101001111000000;
#1 $display("%b", po);
# 1  pi=207'b101111010101111111101110100001010011010111010101111011110001011100000011000001110101111010110011000011100000010001100000101110101101100110110110000010001111010000001111001110011101100001100010010011000000001;
#1 $display("%b", po);
# 1  pi=207'b100100001011101010100100111001000101000000101111100101100101111100101010000111001001010100010000101010001100000111001100101111110100001011010011100101111010101110010100100001010101110010110001010011111111011;
#1 $display("%b", po);
# 1  pi=207'b110011101100011111010100011000111100011101111101001010101010100101100011110011100100100101110001010100000101100110100010011000101001010110101000001001001100101000010111011100001011010101011101001010110100100;
#1 $display("%b", po);
# 1  pi=207'b101000111011100011010010101111110101011001001010001100110001000010011101100101101111111100101000011000110000011111100010010101110110000001000101001001100100011101110000101110101000101100001001100011000011001;
#1 $display("%b", po);
# 1  pi=207'b111111001100101100010000111001010011000100100110001101001111000110111110100001011111000010010000100100001110000100110110010000110110110101000001011111000111101011011100101111110000100010010000111110100001100;
#1 $display("%b", po);
# 1  pi=207'b010001110110001101000000001000110010110111010000111001011001101001001000110111011110011001111010011100101000101010110001000100010010110101011101000100111100000000101011110001111010110000000111001011001101011;
#1 $display("%b", po);
# 1  pi=207'b100010001101000101010100111111100010101111101101110001000001111010000100011011001001001001100010000110111000000011111010110010001110000010110111010101100010010110011100011110001101000100000001101100100101000;
#1 $display("%b", po);
# 1  pi=207'b001001110010010011010111010110001111000110010111111101011011010000100000000110101110111001101100100000011110100010100001001110001011010110110100001000001100010011001110001001001000110001111000001101000010001;
#1 $display("%b", po);
# 1  pi=207'b000010110100100001000000010111100000100100011001001000101110101111111011110110000110000011111010010011110111010011101101111000100110101100101010100111001100110101111101100000100001001010110010100100010111000;
#1 $display("%b", po);
# 1  pi=207'b101101010101100000000011000010011000111011101001011100001010011110100011011001100001011111110001101100110010010111111001110011101101011101001001011010000101100001001011111110010110111100100000100001010001001;
#1 $display("%b", po);
# 1  pi=207'b110011001011000011111101011010110000101011010011010110100101110011100000111110011100111000101011000011100110010010101101111101011111100100101100110000110110000110011110000101001110010010100101110100000100010;
#1 $display("%b", po);
# 1  pi=207'b100111111000001001101101110101011000011001101000001100010110111101110000010101000101110000000101100011001000101000001110001000101101110000110000100010101010000011101110111010101111101111101100011011000110000;
#1 $display("%b", po);
# 1  pi=207'b000001100110110111100111001110110100110101001010101101001100111010111011101110000100101100110100110011000111010001000100011001100101111100000110111011111011100110001110110011001011101001001010111001000110010;
#1 $display("%b", po);
# 1  pi=207'b001101111110101101000111001111010100001110110011001101110101100001010010111111000111111011000000000101101011111001001101010100100010000001010001010011000001101110011001000011001100000010100001111001001001011;
#1 $display("%b", po);
# 1  pi=207'b011001001111100110100111110100111101111111011111001001111001000000010010100010001100000011111110111110011110101000101010110111000010101111101000010101010110110000011010111001001000001100011100110111111111110;
#1 $display("%b", po);
# 1  pi=207'b100110010111101101001100001100010011000101010100100110110001101001010111111010100101011110001000011011001111110001101000011111101001100010100101101000101000000110101111011111101000100110101000011000000011100;
#1 $display("%b", po);
# 1  pi=207'b000110010000011001001001011110100110111001110110111101110111101111001101101110100100010101111111011000010011011101111110110101101010101110101111111111001001101001000000110110000110110001100011100100110001101;
#1 $display("%b", po);
# 1  pi=207'b101010101010100001011100000000100000100000010010111000000000111110101001011100000111011101101101111000101001011111001110011111110110011011110000011000100011111110100000000001011001001101001011100101001000100;
#1 $display("%b", po);
# 1  pi=207'b010011011000101011111111010110111111011100011100011111100001010111010011010111100011010110110111110010011011010000011110001001100010111010000110100001101111110111100100000010001111110111110111001100101010001;
#1 $display("%b", po);
# 1  pi=207'b001111000110101100111101101111110001001000000000001101000011000001000100000011111000001011111100110001000001100100011010100101101001000100111000100000101101010111001000001001101111000010111000100000000010101;
#1 $display("%b", po);
# 1  pi=207'b000111010011100110000010010001011001010000100011110101011110100010111101110001100011001000111110000100110010100110001111111100000011001111101110010111110011100011110100101101111100100110001111100010000000000;
#1 $display("%b", po);
# 1  pi=207'b001100100001100101111111011011100101110001001111111100011000011010111100001101100110000010000110111101011011010111000011101011000100000110110010101100110111110101010000101000101111001000100001010011000111100;
#1 $display("%b", po);
# 1  pi=207'b100110000111101001111010000011101111101010111101111100111011001001111110110010101001110111010100011110111110000111000110101001000011100010101001110110100010011101100011110011010110101110101001110111100000111;
#1 $display("%b", po);
# 1  pi=207'b001101100011010001111101110001100000001000011001010101101110010111000000100011111111010111011010010110110011001101100111110100001100101110111000001101001110010101100000101001001101101001110101110111111101111;
#1 $display("%b", po);
# 1  pi=207'b100101001010000010100110010110010011010000101010011111110000110010111110101011111111110010111111010101110010110100101000001111011001101000000000011001111000000110101111000011011010011110110011110000101110111;
#1 $display("%b", po);
# 1  pi=207'b010000010011010111111010101101101010011001011111011100110000100101010011111101010100100101100010000001100110111100111010001000001011010101101111111111100010011101010000001011000101010101101100101011101011110;
#1 $display("%b", po);
# 1  pi=207'b111000010010100000001010100110101010101000110010011000101001000110010100111101001101111000101011011111000000101010010101011101010000001110100000011010100011001001011110101011010010111000100000011000100011101;
#1 $display("%b", po);
# 1  pi=207'b111010100111001110011101101001100101101100010110000000100110110111001000110100111001100011110011111011101000001011011000000100000000001001010111000111101101001110010011100010010100110111111111011100011011001;
#1 $display("%b", po);
# 1  pi=207'b010101110101001100110001111110110101100010011001001100110000100111100110100111101010010100101001011001110110101110110010110110010001111100000011011001100011001110110100000101111101101011111111001100100000110;
#1 $display("%b", po);
# 1  pi=207'b100001011110000101001011000101011100000010011111001110011011100101000110100000111001111100110110000111001111101010011111111011000001000111100110000100001101011100100001101001100100011000101000101000011000001;
#1 $display("%b", po);
# 1  pi=207'b000010010100011100100100110110111000000010110000101000110010100000100001011110001111110011010111110110010000001110010101000100101010000111110100110010111000110010111110001111111110011010101010001010110111011;
#1 $display("%b", po);
# 1  pi=207'b111101111001011000111100000111110011101000011100001111001000110100100111110000010110000110111001100011001000110111001111111100010000100111110000100110010010111110111101101110011011101110110101110000110001001;
#1 $display("%b", po);
# 1  pi=207'b010101010000001111101110000011100111011100110101100110000000101000110111110100011001011101110110000100100101001111110110000011101111100111100011110001001011001101110010000000000101100000100100000101100111101;
#1 $display("%b", po);
# 1  pi=207'b001100000101101011111010110001101000011100100100000111010100101101111011000000010001001111010001100110110011010100101000111101100111101111011001000001100011011000110011001110101100001000100111111000001011111;
#1 $display("%b", po);
# 1  pi=207'b110001110101010100011001010111101111010001101001011000001110101011000001010011011001001110010100000100111000100000010110100111001011011000100111011011000000100110000001100111010101001101000111100011101111011;
#1 $display("%b", po);
# 1  pi=207'b010111000101111010100001111111011110011101001100110000110001111011100111000101111000010010100000100010111000100011011111000110101001111111111000110100010100010111101001001111000001011010100101010011100111100;
#1 $display("%b", po);
# 1  pi=207'b101010100010100101000101111110000100001111011111100011110110110101000010100110100000011111001101100100000101101110001000101000110000111100110101100011001111011010000110101010010111110100110100010111010011110;
#1 $display("%b", po);
# 1  pi=207'b001110100100011100011001011101011100101010011001110111100101100011000111100010011111111100101001110101110100001001110101000000011010110111000110111000101100011001110100000110110001011001111011110111100000010;
#1 $display("%b", po);
# 1  pi=207'b010110001100100010101000100100111000001111011011100000110100101111001111101111101010011011000011110111001101000001000011110011000100110011100010110000001110010100001100010000110111001010100001110010010011110;
#1 $display("%b", po);
# 1  pi=207'b110100000101100011100000111010110101001111101100101110110000110011000011110101011010011100111100100001100100111011101010010101110001011100101101011110001100100010101110010001101011100111010001010111110100000;
#1 $display("%b", po);
# 1  pi=207'b110011101110001010011101001011110111010110100110010011001101111100000001100001000110011110010110101011001101011010011100001000110111011110000000010001100001011110000101000100001110110010110011111011010111110;
#1 $display("%b", po);
# 1  pi=207'b110001010011110111100100011111110010011100001110100000100111101001111010100110100000110100000010110101011010101011101100011001101101001011101000100010101110111011100000111100010111110111111011111010011001000;
#1 $display("%b", po);
# 1  pi=207'b110011011010100011110000011110010010001011011111110011010111011110011001101001111101001010100010101111011000101001111111010000001010101101000110111001001010010101111000001100011010001110000000011010000111001;
#1 $display("%b", po);
# 1  pi=207'b101000001110110111011010101000010111001110001010011101100101010010110001111000101001111000011111110001000111001101101011000100011000000001010001101001101011110100000110101011101110000101111111001111011101111;
#1 $display("%b", po);
# 1  pi=207'b011111011111001110001001010110011100010010010100000000110111110101001001000101101100100011010100011111101001100000111111100110001000000110101001011111110100000010001010111111110111011011111101110111100100001;
#1 $display("%b", po);
# 1  pi=207'b011000100011110111101000010100110111010101110000100110101101100001111110111111000001011110110011110101111010110011101101000101111100101101011111000100010111111100110000000001001111011110000011010110110111001;
#1 $display("%b", po);
# 1  pi=207'b111110111111101010000101111110001001000101111001101011001111011101000101011111110111000010010010011111111100000001010011110010100011010000010011001010111011110111101010111010111000001011001011101000011110100;
#1 $display("%b", po);
# 1  pi=207'b011011101001111001100100110011000010000011000001101000111010100110010001011110100001111111001100100111111111010010100010111111001110000010011011001011011111110001011111010010000001000000111100100010010010000;
#1 $display("%b", po);
# 1  pi=207'b011001000000111101110001100011011110011101010100000111111000111100111000001011000010101001010110111100100100101111110100001111000011100011010011111110111111001111110010111101001100101001110111110001010010100;
#1 $display("%b", po);
# 1  pi=207'b100001000001000110100010111000100000001111010010000000000011100110001111010010000001101100101001100110110010010010100101001100110100111101110000010001101111110000011100010111010010000001100000111011111011000;
#1 $display("%b", po);
# 1  pi=207'b100001111101110010101001001101111001011110001010100011110110011100111100001110101100010111001001111100111101011100110011011001011101100001100011011110011110100000010010001000011101111111100111001110011010011;
#1 $display("%b", po);
# 1  pi=207'b110001001001100000010001110010101010111110111111100010010100010011011000011000101011000110101000011110010011101111100010100101110111011110110101100001101010100111010100001010110011000000111110010110011111110;
#1 $display("%b", po);
# 1  pi=207'b011100111111101100011101010010010000101100100011001101110100011100111111001101000110000001001100100000010100100100101001010000000011100011110111000011111110010101111101100111010111101101001000111001100111101;
#1 $display("%b", po);
# 1  pi=207'b110100100110101111011100110110011111000110111111001111000001011111110110101100010001100000000111101010110000010100100110011110111010110010110000101001000010001010011101110011000011111110100011011000100001010;
#1 $display("%b", po);
# 1  pi=207'b000010111101111010111001100001100101100011011111010010100011011000011001010000000000111000100011101001110001111101100101001111100111010110001100011100010111110110110101100111000000010001111111010101110001110;
#1 $display("%b", po);
# 1  pi=207'b011110110000001100100011011010100100100000110100001000101010001111001111011111001010101111110001110010001100000011101011010111010001000001010001110010111010100100010000111100101100100010101111010001111100111;
#1 $display("%b", po);
# 1  pi=207'b000101111011100101010011000010100000100101111100111001101110100110010100110100011101010110010011100101111110010000010111101010010000001110000101000101111010000011100000000010011011011111001100000001100110001;
#1 $display("%b", po);
# 1  pi=207'b111010010010011100000110000100000101010110101110000101101011100001101101010011110000100000111100010101100101110010111001111101100000100000011010101100111101111010000000100111010100110110000100101110100001011;
#1 $display("%b", po);
# 1  pi=207'b010001101011000110000010011001011100110100000010011101010001100101101001101111110101010111010011111010110001101101111010000110111110000001100100010111111100000110011000101110110110011000111101001100010111011;
#1 $display("%b", po);
# 1  pi=207'b100111110110010110011000111111100111000011111101111000000111011011011000110100011110101000001001101001010011001110010000111110011000101110110110111101011001101111011100001010110111111010110010110000101001010;
#1 $display("%b", po);
# 1  pi=207'b011001111101110001001011100101010000001001110010101101011111111000101101110101011010110001001101000010011010000001110011101100101100101110001010011000100001110101100000010111111010000001101000010101100110100;
#1 $display("%b", po);
# 1  pi=207'b000001011110110101100111000111111000010100000001011000110011010000111010110001101000010010010111100010101110101100011001110010101111111111111100000001101100000000101000000000010011000001100110100101100001011;
#1 $display("%b", po);
# 1  pi=207'b100000001001101011110011100110100110011110001110010011010110011011110100010110001111110010100110000000111111101011000000001001110101101100100000101000100010101001111111110111000010000110011010111111001011001;
#1 $display("%b", po);
# 1  pi=207'b100111000100001010101111101100101001011011000101100010111010101010101101011001001010001001101100100010100101100011000111110110111000010010100101010010111000011100101011101001110010101111110101111101011010101;
#1 $display("%b", po);
# 1  pi=207'b010010111111100011010111110011100101011001100001100010000111001011111010001011001111100010000110010011010011110000100001100010000100001100000111000110000001001010000000101011011111010010100100001111010001000;
#1 $display("%b", po);
# 1  pi=207'b100001000100011110010100111101000000101001001101101000111111011100111110000010001011111101111011100000000101110001001100110100010111011011010001101101010011011011010101101111101111000001100001010100011010111;
#1 $display("%b", po);
# 1  pi=207'b101110000100011110100110111001001001110010111001000101101110101011010010010110011000101011100101111011110101001100001010110011100100001111101110010100100100011101001010110110010110010111001111111100001010111;
#1 $display("%b", po);
# 1  pi=207'b010010101111001110001100101101100001101100110001110100110011010011110110101110001101101101010001101101110010110100001011110110010000111101110000110000101000011001001100001000000111001010100110000010101110110;
#1 $display("%b", po);
# 1  pi=207'b010000111011110100011001011001110000110001001111111110010010101010001010011010010000011010001000101110011010101011110001000010110100110011100011100101011001011011001111010011011100111001101011111001100011110;
#1 $display("%b", po);
# 1  pi=207'b011100101010110100110011110100000110001101111010100011000010011111101011010110110010100000111001101010011111101011010010100100111011010111000011110010100001010101001001010100001110100000001010001001010101010;
#1 $display("%b", po);
# 1  pi=207'b000011111111101110100010100100011100000111010111001110111111111110011011010001111110101111000011111000101110100001110101100111010110001111110000101111111101001111010110111101110000101010100111001111010100001;
#1 $display("%b", po);
# 1  pi=207'b110011000101010011111100110011110010111011110110011110100011011101001010000111110011000100001101001010001101110101011111100011111100010100001100111101011011000000000101100100001000110000110010011100100010010;
#1 $display("%b", po);
# 1  pi=207'b001100111011001001001100110001111000111010101100101011001110101010011010001000101010011010101001001000100110011001100101100111110010010100000011000011111000110011001101110100011000011010100100000100001010001;
#1 $display("%b", po);
# 1  pi=207'b111101100000011001001000010101001101110111100101110010101101110011101111001010110011011011000101111010001110010100011100100111011100000010110011011100100011100000101101000100011111111010000110101010100000111;
#1 $display("%b", po);
# 1  pi=207'b110001010001011111010111001101000111100100001100010001011001110110010010010101000000110111000101011000110111101010111111100101001101000000100000000101011100000101011100010011000010111101110110101000101000100;
#1 $display("%b", po);
# 1  pi=207'b001111100000110011100110111101000111010011000010011110101101010100000010100001100110001010011111100111011110100101100111110111000111001000101101110011001011011001110101101101011011000100111010100101010101110;
#1 $display("%b", po);
# 1  pi=207'b110000001101001001100001011001010111111100011001001110111010001001010101010000000110100111000110100110110000111011001111100000110100001101010100010111000110110110001001101001011100010010010100110111101011100;
#1 $display("%b", po);
# 1  pi=207'b110000110101110010101100111101110100011100111001001010111101100110010011011000111000001010111100000100011111101001100110001110101000100010110010101010110101101111111100010110001101101101010101110110000101110;
#1 $display("%b", po);
# 1  pi=207'b010010101111000111010011101000100110001101011000111110111011000001111111001010111111100111111101111001001111110110100111110000110101000101010101100011000011001000111000100100001000001110010110100110001011010;
#1 $display("%b", po);
# 1  pi=207'b011000010111000000000110111100110100000011000011100000110100110011000001100101111001100001001111111001010110010001000011001100011000100101011011001011101111110111100010011011011001101001000101011010010111001;
#1 $display("%b", po);
# 1  pi=207'b000110110000110111101100011111111010110001001011000111110010010011110111110011110001110100111011100010110110001010000001101011110101011000111010010110000101001011011001110010101111010100000001010101010010110;
#1 $display("%b", po);
# 1  pi=207'b111100001011100101110010100011000001101010110000010011100110100011001111010110011100111100001100000010011001110000001100010111001010000100111011010111111010101110010110001110110010001000110100111000111101010;
#1 $display("%b", po);
# 1  pi=207'b111000000110100100100001100010000111001010101111101101000001101010100001010101001110010100001000001001100110101111111001101100110100100111111010000011101001101010100000100011110011100100000001011000110001011;
#1 $display("%b", po);
# 1  pi=207'b010111011111101101001000011010011101010111011000110100100101000100100100100010101110110010110000011011010100100110011101001001001111001100010101000000010110000001101011000001010111011011101000100011110100011;
#1 $display("%b", po);
# 1  pi=207'b101110110101011100101011011100110100110000110111010001101001100110101000101001110110101100010110110100101000010011001001111100101000000110101100010101011111101011001001011110011101101111000011001111110111100;
#1 $display("%b", po);
# 1  pi=207'b111110001010001111111001001001100100011100001010000001111011001011000001001100101000111001100000101100100111111111101011101010001111001000010000011100111010110100000100100110110001001000011101000010011001001;
#1 $display("%b", po);
# 1  pi=207'b001101101010101100000110111010000110100001010011010110001001111110111101100110011011100101011111001001100111010110010111111011110111000010000001100001001011010001111010111101011110100001000100001100001011011;
#1 $display("%b", po);
# 1  pi=207'b100001000100011011110110101010111011110000100010101111000110110000001100000101001101010001000011001110000001110011000110001101101010010000110010100101101001101011110110011001101000101110111010001010111110100;
#1 $display("%b", po);
# 1  pi=207'b111010111101111010110101101111110001100001101001010111101111100001011001111000010011111110011100101111101101010101101100001101101000000100101101101100101011100000010110100011011111111010101001100100101110010;
#1 $display("%b", po);
# 1  pi=207'b001010010000000001100011011101111101000101111110101010011001011001111010100001100010110010110011000111101010000000100010101111101001010011110000010001001101111100100101011001001001111111011111000100101001101;
#1 $display("%b", po);
# 1  pi=207'b010101100101100001100010000110000000001011000101010001100001100010010110011001110101011010101110001110100001101110011000111110100011000000000111100111110110011001010011000110010000110000101010001110110100011;
#1 $display("%b", po);
# 1  pi=207'b111100010010011100001110001110001111010001101011010001011001110001100100101111001110100010011100111111010111100101110001101111010010011000100101110110010010001011011100100010111001010001011101001000010110100;
#1 $display("%b", po);
# 1  pi=207'b110010100001111101100100010001011001101000010000011001110000000101010000001001101111101000111111110111110110101011100110101001010000100111111011100010110000111010001001111100001011011011100001100000101010111;
#1 $display("%b", po);
# 1  pi=207'b011101001011110101011101011100001101111100100001101000101101110010011010010010101001100010111100011001100101000000101101011010010110001111011001100111001001000011110110000010011110110110011110001111000101110;
#1 $display("%b", po);
# 1  pi=207'b000100000011010111010000100111101001101111111010010101001001111011010110001000001101100100101100011010110010111000101111010110100100100111111101101000100010001111001011000010100010001101110110100001110100011;
#1 $display("%b", po);
# 1  pi=207'b010000110111110101000101010010110001001110001011101100010101010001100101111000010000011101001001101111110100000011000100011000110001011001001101011000001111111011110101111111011110101111010110101010001111100;
#1 $display("%b", po);
# 1  pi=207'b011000010011001011001111001011111110100010001001000100111100001000001110000111011101001111010000101110101000011001100010010111011001010100101101000000010100000011000000000100111011110111010001100100100000010;
#1 $display("%b", po);
# 1  pi=207'b111000010111110000011000111110010000111111100101000010111010101100001000010000111011101100010101011101100111000100110010111100011110110001000100111001110100000110000000000100111110110001100100110111010000101;
#1 $display("%b", po);
# 1  pi=207'b111000100111101100010101100010010011001111000111110101001011011100110101100000010010101101000110001000000001000101011110101101111010011100011010110111010111011101110100110101111100101010010101110111110101101;
#1 $display("%b", po);
# 1  pi=207'b111001001100011111001110110011111111000100011111101111001000011000111010100101101110000100000011101100011111101100010000110001110001011011101010000010110001010011010011011100001010100110110100110110010111111;
#1 $display("%b", po);
# 1  pi=207'b000110100000101000101010101111101010110010010101000010000000111001010100010100000110011010001100010000111110010000111011110001010000100111111011010110101110110110110101011111011100010000010001100001011001001;
#1 $display("%b", po);
# 1  pi=207'b010000000100000000010100111101111010000110000001011001111010010101010101100001110111000001110110110010110000010101101111101001010011111111010111000010010001010100110011101001011000010000001110110110100111011;
#1 $display("%b", po);
# 1  pi=207'b010010011101001111011100111001011100110101001101000110011111000011010101101100001101100000100010111010101001011010110100111010011011001001110001000010101111001011101110101001111111100111111010001000000001010;
#1 $display("%b", po);
# 1  pi=207'b110110011011001001111011000001111011100011010011100011100010000010100000000100100101010001110111011100011100011101011110111100110101111111111101011000000001000101111101101100100010100100001111110000011011111;
#1 $display("%b", po);
# 1  pi=207'b100110001100110100111100101101000011011010111110011001111001100100010101000100101001100000111110110000111010100000111010010101101101100101110110000011000101000101001100000110010011010110110110100011100100111;
#1 $display("%b", po);
# 1  pi=207'b011001110111001011011001011101111011110010000011101011001011001000001001100000101000010100110000101001000000110100001111100010010001000001111100111110011010011011101000001101001010110001110001100011100010101;
#1 $display("%b", po);
# 1  pi=207'b001010110110110111000000101100110110101111100011101101000110110111100000000111011000100111101010110111100010101100010010001011111111101111101110000110101110101101011111000001001000101100100000010000111000000;
#1 $display("%b", po);
# 1  pi=207'b111000000101110100111000010100111010101011100000101000001000000000000111001101001001110111110000111000100110001111001000000011000001010101001000101001011011110111010010011010010011100000101100000101110011001;
#1 $display("%b", po);
# 1  pi=207'b000100001000101101001000010101011001010100000011110101001101000111100000111001101010010110110111110011011100010100000110000011000101110011000110001100010101111110101001100100110100100110100011110000000110010;
#1 $display("%b", po);
# 1  pi=207'b101100100101001000010010110110110011001010101110110001000001001010011011000101010011011000001110100011110111000011100100101110000001001010011011001100110100100001101100010000001100001010011010101100000111000;
#1 $display("%b", po);
# 1  pi=207'b000001000111011110110101111010101001110010110010111101101011000010010110111010111100100010000000011101100100111100101101010100011011100110110010010010101011011100111000001010000110010001101010101111000011111;
#1 $display("%b", po);
# 1  pi=207'b001100111111111011110100011001101111111100000101110000111100011011010101000101000110010100010000000001011110000011011110011100111001100001110001010101010100001100000000010000111011100001100010010110010100000;
#1 $display("%b", po);
# 1  pi=207'b001110001000000001101011011010011011111011000101100010001110111110000110001100110100011010100101110000111011111011000111101011011111001100101100100001001011010100101100110011110101110001110101101101001000011;
#1 $display("%b", po);
# 1  pi=207'b111000111101111101101100110001010011110110011001101011100001110000111000101110010101010110001001011010000000010101111110101011101011001101100110000100001100011001111111100010001100000110000010110010000111100;
#1 $display("%b", po);
# 1  pi=207'b010010101011000000010001001000101101000000000111001001100111111101100101011010111000000110011000001101000110100010011000101001010001011111011011010110011101100000010100010111101111001000101000101110000010010;
#1 $display("%b", po);
# 1  pi=207'b000101111010101111100101010000110001100011101011111100010011001011011111010110110110111011101000100110000001111000011010101001001011101110101100001000111011001010101101100010101001011010010100001000001000101;
#1 $display("%b", po);
# 1  pi=207'b010000000011001001011010111001000110111001100100010111110010100000111010111111100111001110000111101001100100101100011011101100100011110110010010010100111000100101000110110100011101101001110110011000100101101;
#1 $display("%b", po);
# 1  pi=207'b111000101001101100110100001001111010100101110110111001001101000101100001011110011110010110100000100111100100010001011000000000000100001101000000010111100011101111110001110100100101110001000001101110011001001;
#1 $display("%b", po);
# 1  pi=207'b000011111011001001011111110111101010111000101111111100110111010000111000001011111100000010111011010110100110100001011110010010110010101011100111001000010011110000100000100101100000110110111100111011011001011;
#1 $display("%b", po);
# 1  pi=207'b011011111101100111010001010100100111011010110110000101111011101101101100010010000010101110011101010010100100010100011010001111111000100001010101010011110101000111011111001010110111010100101000010010110010101;
#1 $display("%b", po);
# 1  pi=207'b101000011100101011110100100001111011111000001101011111101001011110011000001111110110010001010110101110110110101011111110101001111100011111010110011111111100000100101111100101110011111101100000100001010101010;
#1 $display("%b", po);
# 1  pi=207'b010111000011110110001101110010001000110000000010011110110011101101100000001011110100110000000111000011101000111001101111010001110010101100110111011110010011111111011111111110001100111011110001000010110000101;
#1 $display("%b", po);
# 1  pi=207'b111110011000110110101110010000011100101000011011000111101011010001011100110110100111111000011001001011101100011111001000111111100010101001100000110011101101001000100111100100001100110101000110001001100000111;
#1 $display("%b", po);
# 1  pi=207'b100001111000100110011101000100100101111111011100000011111111111011001010011100001010101000111011000101010010010011011101100011111000101011101000101111000110101000001000000010001110001100000101000101111010110;
#1 $display("%b", po);
# 1  pi=207'b101111111001110110111011101111000001010101111011110001000010011110111011101001110111000101110110000101001100000100010011010100110100011110000001001011110101111110100000001001110001001011100110010010011111010;
#1 $display("%b", po);
# 1  pi=207'b001000010100100110101100111001001001110011000001100101111100110000100010001011011010000110011000101101011100010100010111010100001011010010000100110001100111010000010001101011100000111111100010101000111100001;
#1 $display("%b", po);
# 1  pi=207'b110011001100110110010011110011110101101010110011110011101111011100011101110101011000111011000001010111001001001111000110101010101110010010110000001101110101111000101000010100011011101010111101001110001011011;
#1 $display("%b", po);
# 1  pi=207'b000101100011000011011111111101101011000100111101001100100100111001010110010011111100101011010000011000110001100101010000010010000111000101100000001110000101000100011101110111101011100110001001111101011000101;
#1 $display("%b", po);
# 1  pi=207'b011000010100111010011100000101111001101101101000100000001011000010011010010000010111111111100111101001110100011100010011111111010111000011101010010010000101100010001011001011001110010001011100010011011000010;
#1 $display("%b", po);
# 1  pi=207'b001001010000110101000101000000001111111101000001010000000101001110100010001010100010111110111011101001000111011100111001011100010001100000010001010101010001110111101001111101000101000001100010000000101011110;
#1 $display("%b", po);
# 1  pi=207'b000001000000100101101011000110011011111101110110011110001111101101010010100100000010011010000001111101000100100011010010111001001100001111001001011010111010011001100010101010001010100011100001010100010001111;
#1 $display("%b", po);
# 1  pi=207'b110110000001011011101111100111110000001100110101010000000111100010001101010010100110101110101111011101010010001001000101111001101000110001110100010010101011110111001010100101001011011111011110001010110110110;
#1 $display("%b", po);
# 1  pi=207'b010101111110011010111101001110010101001000010001010110011111011100001100110001111000010001101110111001000100111110101001111011010110010011001000110110100011110010001000000010110010111011101000110100110101001;
#1 $display("%b", po);
# 1  pi=207'b011010100101100011011101111011011011010010000011110000000010010100000100111010000101001010001001001100011000111001011100011011101111001110110011101001010111100011000100111010100010111111101000010111101111000;
#1 $display("%b", po);
# 1  pi=207'b000010100101101011001000110000011100010110000111101000011111001000001011110010101100110110101101111111000000011010100111100000111001001000111011001100000000111110001100111000101101101000011101010111110110100;
#1 $display("%b", po);
# 1  pi=207'b001010001100111101000011101101101001001111001000000110000011011111011111101110101000111110001101110000010011010111110101001010010110000000000000101100101100101100110101000011111011000001000110111111000010010;
#1 $display("%b", po);
# 1  pi=207'b011101000010101001110110101110100101010101000000101001000111110100000100110011111110011000100000110100001111111110000111010000100111001010101010010111001111101100011010001000010111111110000001110000011100010;
#1 $display("%b", po);
# 1  pi=207'b100011110111101011100001010001011010101101000100111110000000010110111111010011001111000001000110111001111100000000000111110010001000101001011101101100011110101010010000010110110100001100000100100100000011101;
#1 $display("%b", po);
# 1  pi=207'b100000011011010000100010010001001101010001010011101000111011010010001111100001001000100110110100101000101111011000011110001111111010011101010111001111111101001001010100100100000101010111010111010111000111000;
#1 $display("%b", po);
# 1  pi=207'b011100011000110011101110001101101100100100110011001101111100010110000110101100001010000110110101010101101011110000000001010000100010101000100011111100111001100001001000100010010000100111000110010110010011110;
#1 $display("%b", po);
# 1  pi=207'b010011011011010011100110000100000101111011110010000101001100000010010010011101100110001010010111110111001100000000011111111001101100011101100100110011101011011110001000000100111000011110010100010110001001011;
#1 $display("%b", po);
# 1  pi=207'b101010001111001100011011011011100100010011001001011000001010010001010011000000011001001001110101101100110010001110110010101111100010111110111110101110000101110100011110010000001100010000000001100111000011001;
#1 $display("%b", po);
# 1  pi=207'b000110111000010011100101010010010011000010000000000111001000101000011001110100110101000101100001010000011011011111101011111011010100001010100010011011010011101111111101101100011110110111000111100010010101010;
#1 $display("%b", po);
# 1  pi=207'b100011101110001111010110111111001100011001100111001010111101111111001111000000010111101101101010001001110101010000110001000001110001011001111001100011100001011100000000010010011000011010100001000100111101011;
#1 $display("%b", po);
# 1  pi=207'b110101110100101011101000000101101101011100000100111011000111100100101111011000101101001111101011000101000111010110001100010000011110001110011101001000100010111011011011010010101000101010011101011101010001001;
#1 $display("%b", po);
# 1  pi=207'b111011110101001100100111000000110111111101001001011101010000001010100111000111101000110010111101011101000011100111101000001000101010110010101110010010100010111110101000101001001110000000100000011001100011111;
#1 $display("%b", po);
# 1  pi=207'b001011010001011101011101000000001000010010111010110000110100110000110100011101000011011010101101100000001100101000110101101001101011000110000010000011101111110111011011010111100110101011110111111110110101110;
#1 $display("%b", po);
# 1  pi=207'b010111011111011010101010100001001111000100001010011010001111001010100010111001001101101000001000011001011000010010010011111111010010000001110010011001110111011110000001111010100000010001010111000100011100011;
#1 $display("%b", po);
# 1  pi=207'b010001011010010000100000001011011100011100100100011101100110110101000110100100100011100111011000111111111001001111100110001101001010000000100001101010110011000010000011000010011001100101100001110000000000000;
#1 $display("%b", po);
# 1  pi=207'b000000100110011000011011011100000001111011011011110110110100000110010111101110101001111001101010011101001000100100010101001010001000000100011001111111110011001010001101111110100111010101001011001101000001000;
#1 $display("%b", po);
# 1  pi=207'b101111101110110011001101101000001101011111010011011000100011110101101001100010100010000011100011111101010010111100001010111000011001101100100111001000110100001001111100010101111101100110000000011010010010010;
#1 $display("%b", po);
# 1  pi=207'b000110111011010100111101101110110011001110100111010100111101111000111001010111101100010110000011010011100100010101000001110010101111101100011111101111000101001110010111010110101001101011001011011110011101110;
#1 $display("%b", po);
# 1  pi=207'b011010101100110100111101110101011001101010001010100101110000010110100001111110101101011010001110101101101111100000010010010110011001100001110100010110001001100111100011101001010100010111000101100110100001101;
#1 $display("%b", po);
# 1  pi=207'b100001010010101000100101110100111000010110100100010100001000111110110001001000011010001100110100011100010000100001100101001010110000111010111111010101001010011000010000001101011001000011110011010101100010010;
#1 $display("%b", po);
# 1  pi=207'b000111101100110111100101101001011010101010100110101100100111111010111001000001100010000010000100001000000000111010100101001111011110110100011101001101101001011101010011111000100110010101111010000001001010010;
#1 $display("%b", po);
# 1  pi=207'b001101010110100010000111101111100100100110010001010010111100100001010011101100110010001011111011000010111001011101110001000111000101100110010011010011111110001110010000111000000101100111101111100000001000101;
#1 $display("%b", po);
# 1  pi=207'b001000110000111011010110100010011101111101000001110000000110101000110111101011000011100010100010000101100000000010010110000101111111110111000000111010101001010100110101001000001001000001110100101110101001010;
#1 $display("%b", po);
# 1  pi=207'b000011111001110100111110001001101000111100001000011101100011100011010000101101100101110001011001101010111110110000000101011000010110111010111111101010101001000001100101000001011101110110001101110001100101001;
#1 $display("%b", po);
# 1  pi=207'b001011010100010111000100011010010010000111011100101101110010111011000010100101110100110000001010000100011001010110010111010110100100011110011111011011010110111001001011011100010100111110011010010000111010011;
#1 $display("%b", po);
# 1  pi=207'b001101111001101101000001001101011010000111100001111001100100100101010101100001000000001000111100101110100110010001100001100000101000001000101101101011111110110101110011110110000111000001000110010100111000001;
#1 $display("%b", po);
# 1  pi=207'b010001100000011001000110111111100111111100001001110000011110101100110000011101010011100111111001001111000001100011100000111000111000001001011101011000000000101001101010000000000011101100010111100101010100101;
#1 $display("%b", po);
# 1  pi=207'b111000101000010010001010111110100000010101100001001011111001110010011001101100001110010000011101101110101011010100100000011001001111101000100111110001011011110100001001011110110110000011010101000101000101101;
#1 $display("%b", po);
# 1  pi=207'b110110100011010111100010101001001111011001011000001100000000101000111101001100111110000110010110110110010100111000101010001101111011111011001110110011000110110100101101110011100011101011010001010111010001001;
#1 $display("%b", po);
# 1  pi=207'b101111011001000010001110010001010110010101010101010110101011000001111001101010100010110001101100100101101110001100000110000110110100001000010010101000101011100101011000101100110101101101010010101100011011100;
#1 $display("%b", po);
# 1  pi=207'b100010011101011100101000011110111101000010000001101101001111110110000100001111000101101001011101011101111101010000000001011101101100110111100000010011101001010110111110110010110011011101111001010000101011111;
#1 $display("%b", po);
# 1  pi=207'b011101011110100011001000001110011000100110100111111101001010001100111011101100101000010010100011001000111000111110100100010111100110111101110101100010010010001011010001111011000010000110010011111111100000111;
#1 $display("%b", po);
# 1  pi=207'b100001001101100110110101110001110111010010100011000111111100111101001110110010010010100110111110111110101110101001110110101111110101010100010110001101100111011100110011110111110101111111011000000100001101001;
#1 $display("%b", po);
# 1  pi=207'b001111100101111000001001111001001010001010001011111011010101001111101010100110011100001011111001100101011000110001000100100000100000111111001010001011010110000011000010001010011000100110011101100010001101101;
#1 $display("%b", po);
# 1  pi=207'b011101111100011011111101010101011110100010111100000001001110000111011100001011000110010001011011010000101101000001100010101011001110011001101111111011010010100111101010001100111111110111010100011101001010001;
#1 $display("%b", po);
# 1  pi=207'b100000101011000110001001000001011110101001100000010111101100000101001010000111001000101111110010100101101000001110010000010101000101101111010010001011100110110101001111000110110010010111010011110001111111000;
#1 $display("%b", po);
# 1  pi=207'b000111111000010011001101111000101110001010101101010000000011101001000111110000011111101001111110100000100101101010110100011011101101100111001111111011111111011001011110000101011111010011101100010010101100101;
#1 $display("%b", po);
# 1  pi=207'b011010101111101111000111101101101010011101000100111011110110100000111010101010111111111011100111001111111001110111001101010110011110100101101011110000000111101111110011111011001110001000111001100101101001111;
#1 $display("%b", po);
# 1  pi=207'b000110100000111100111001101011010100011100010000110110101111101110100010001111101101011010111110010111110100010111000110110010001101100000000000111111111110001000111000001010001001010010101011110010000010101;
#1 $display("%b", po);
# 1  pi=207'b111011011110011010010101001000000101110100111010001010110101001011101111001001010011110111011111010101101010101010110011010111010100011011101110000011111110101011100001011111011100101111000010011010010000101;
#1 $display("%b", po);
# 1  pi=207'b001000010001100010110001110101011111000100111011111111010101100111100100100100100101101100010100101101010011100011100111101000111100010011101111101000010000010111011011001100011100000101100101001001000001000;
#1 $display("%b", po);
# 1  pi=207'b001011011001010000000000010100100100000100101011010100111010001100110011101010000100000000100001100010110011110001000101110100100000101110101011000100101101011100000000110011011111001100000100101001011000010;
#1 $display("%b", po);
# 1  pi=207'b001000100101011101001010101111110000111000101100010111110010011101001110010000100110011111000101110011110111111101001111101011101111001001100101101110011000111110000000101101101001111001111010011111100010011;
#1 $display("%b", po);
# 1  pi=207'b111000010000001000010010110000001010010000111000101011010011000001010100111101111010011011101101110101100101110011111100110011100010001010001011111111101100110001000100011100101000001111110110110101001010011;
#1 $display("%b", po);
# 1  pi=207'b101110100110111000011000110101011001110100100011000011000000000110010100001001000111011100000110011010001011001001111001111101010010000111110111111010011001000000111110111010111010111010111011100100110011100;
#1 $display("%b", po);
# 1  pi=207'b100011001000111010011101111000100101010100000110011101111000011100011101010011010111100011110010011010011001110101010000001110111110101010001011000101011110010001110100111000001110110111011001001001000100001;
#1 $display("%b", po);
# 1  pi=207'b111100110100110001001000001011101011001100000001111000101011100110000000010000110101010010101000101000001100111011101001001000110010110011010001100000101011000010011010000010011100101100101010001100000010101;
#1 $display("%b", po);
# 1  pi=207'b110011100111101000100000111010101001101110011010011101000101111010000011010101111011011111000110011110011101101110000011000010110010111111010001010011111010001000000000001000110010011001011101100010111001100;
#1 $display("%b", po);
# 1  pi=207'b101011111000001111111101010001111101001110110000011100001110101101011101001111101101111001110011000100110100110000010001011101101101101111001110001011111001100110010111100010010100111010100010001010111010001;
#1 $display("%b", po);
# 1  pi=207'b110111100100010101010011100110010011010001000011010000101001001001100010000001001111111101101001101000101000000111111000001101001101110100110100000011101100010000011001100000110111010011110010100001111000101;
#1 $display("%b", po);
# 1  pi=207'b101001010101011110110110100101110100010011010010110100110000011000011101100010001010001100001010110011001001010100010011100001010001000010100100110111100111001011100100101101101101100000001000100110011111101;
#1 $display("%b", po);
# 1  pi=207'b001001001010100010001011000111110111011000010101111010100110110100100100100010011000101110100100011101010101001010111000010011101110011001011001000110110111101110000101001111110001000101011011110101010000110;
#1 $display("%b", po);
# 1  pi=207'b111000001100110010111011000001001000100110011111110000101000010101100100010111010101101010101111010111100100000011000001111001001010011001011100000010001100111011110101100011101010001100001100001111100111010;
#1 $display("%b", po);
# 1  pi=207'b111110101110001001111011110000010001000010000000110111100001011111111111000001101110000100011010110101110110100100110111000100000100100011110011101001101111000101100011001100000100100001101101111001101101101;
#1 $display("%b", po);
# 1  pi=207'b011001111000000110011101100010001100010001110110001011000111011101000110101001010010111110011000111000101100110011010000011101000100110010011101111001100111100100101111000110110111110001001100110010111111001;
#1 $display("%b", po);
# 1  pi=207'b111011001000011000101100000011100100100101100001010100100011011101010111100001000000110010111100010101000101001000110110100100010110110010110000110110100010010011011110001011011000110101010111010110000111110;
#1 $display("%b", po);
# 1  pi=207'b110100010011010001110110001101101001101111101010000111000000111111010101011101000110011011010001111110011111000001111001000101110101101100111110111010001101010000001101101011011111100111101011010101011010110;
#1 $display("%b", po);
# 1  pi=207'b010001101000101010110111110011111010101111011101111000111111100001011011000010000010111100100000111000111111110011100100110100000011001101010101001111011011010001010100101100100110100010001110010010001111011;
#1 $display("%b", po);
# 1  pi=207'b010110100110111000001111000000001100001100011100000010011111000010001000110000111111000011010101011110011011000110010110101100110100110000110001011111100100000011110001110001010001111110110100010100111111001;
#1 $display("%b", po);
# 1  pi=207'b111111011111101111011001010111101001110110000101101101001011001111011010001010111001101011001010111011001010000010101111101010011111110000101001101110011111011100011110001011000111000010101111101001101111101;
#1 $display("%b", po);
# 1  pi=207'b111000011000011110111101001111010011111001110100101111100111100111100101000110110010010111111001110111010010110001110001111111100110011111000101100101000110101010001001110010101100000010000110111101100000100;
#1 $display("%b", po);
# 1  pi=207'b000100101010101011100110111101100000110001001010000101010010011110100101010111010011100010010111110100001110011100000100000000010000010110010111111110010110101010001110111100100001100101111001110000001000100;
#1 $display("%b", po);
# 1  pi=207'b101001111011001010000101110000000110111111001100110110010000011010000010110011110100000011011111100010101101110101010000001001100001110011000101100000010111010011001111101101111100110010111100011011110111111;
#1 $display("%b", po);
# 1  pi=207'b000011010001001101111000000100010111100011111001111110010011001010011110110111011001100111111111110011110011000001010001110010011101001101101100110100011011111001000111110110001010011110101101010001101111011;
#1 $display("%b", po);
# 1  pi=207'b010001110000001000110100111011010001001100000011100000011010111011000101000000010010110010010011000100100101111100111101111011110011110000001111010111100010100101111010010111110101001110100100110110010000001;
#1 $display("%b", po);
# 1  pi=207'b000100111100110010111110110000110101000001010101000011000100001011010010110100110100110000111101011011101111001110001011001011101111011111010110111000101100111010011100100011111100010010001101100110101101010;
#1 $display("%b", po);
# 1  pi=207'b011101010001011110111110010111011011000100010101011010110010110001101010100000010011010011001011110010100000000010100010101011010111011001111001101011000010111011101000110000010110100001100111110010111101011;
#1 $display("%b", po);
# 1  pi=207'b000101110001011110010111010000100000101100000100000110001111010111011011101011001010010111010000010110110011111110101110001111110100001111011100111011111100111011011110010010111011101111000010001111001100000;
#1 $display("%b", po);
# 1  pi=207'b111100010011001101100100011001010000000111000111000000101111011111101001011000000111011111110010011010000101111100001011110001101011001001001111011101011000111100000010001111101101101010100101110100110000011;
#1 $display("%b", po);
# 1  pi=207'b111011100000111101001110101001111100100101010100110011000010010010111001011101000001010111111110010011110001000000011111000010101000011001110110011000000000001001010100100000101001010101000010101111010100011;
#1 $display("%b", po);
# 1  pi=207'b101001010000001101111101110001111011100100001100100100100011100100110000111011010010101001001011110100001111110101000111101010101010011011111110000100111100110010100000111010000001111011011110011011011101000;
#1 $display("%b", po);
# 1  pi=207'b111110010000100110101011011100001111001001011110110110010010110100000010101100011010110110111011111010100001001010000111110101010001110111010111111010010001000111111010000010110110100110001110110111000110101;
#1 $display("%b", po);
# 1  pi=207'b000010111000010110000101110100101001101110111000011100011010100010001100001011111101101111101110100011001111000010011011101011001110000000100111000011000011101010010101000001010000001100011111110101110010111;
#1 $display("%b", po);
# 1  pi=207'b100101110101101110011110101111001111101011111010100111010000011101100011000100111100001011000111010001011111101110100010011111110011000110101000111011100100111110001101111111001011011011110111011010011011110;
#1 $display("%b", po);
# 1  pi=207'b010000100000010111001101101011010100110101111101000110010101111101000011110100010100011110001001111011011110010111011101001011110110010100111001101100111110000110001000111010000011010110010011100100001110011;
#1 $display("%b", po);
# 1  pi=207'b101001010110000000100101011100111010010101011101011100011000011110110010000101101001111110110000110101010000100111011101000111010010001000100110001001010001001000111100100110100100010001110110000001100100111;
#1 $display("%b", po);
# 1  pi=207'b101001010111001100000000001101011001000100101111111100000010001111110000111001111101011001110001110111110000100010011011101010011101110111101000000111010001101011000101000010100111010100111000000111100110110;
#1 $display("%b", po);
# 1  pi=207'b111011010111101010000000000111100100110111101110111101100001000011011101010101101110110010011101010100100001001111100101000000100010111011111101000011110111010110001100110011111100100100011110000100001011000;
#1 $display("%b", po);
# 1  pi=207'b000110111100001001001111000101001010010101011100111111100000111111000101100001111000010011101100110101110010101010110000101101011010011001101100100000100010001011000110110110111011101101110111100100001110011;
#1 $display("%b", po);
# 1  pi=207'b001111010110101010100110001110111111100111110101000010111001010110101111001000111001110100001111111010011001001001010010110100010111111101111000101101001001011101111000000000111100010010111000111010001111001;
#1 $display("%b", po);
# 1  pi=207'b000000001010101110011101000001001010010101000100000110101101100101000110100111110011111111001000101100101000010011011000111100011100000111110010100011101001101110101101001010100111101100101001011101001111110;
#1 $display("%b", po);
# 1  pi=207'b001001111100000100011001011101000100001110111011010101011101000001111001000101011011110011100000001101010001010110101111100101001111000001101100001111000000101011100100110010000000000100000111100010010011101;
#1 $display("%b", po);
# 1  pi=207'b111110110111000000100111100101110001001011111001110010010110011101111011111100101011011010100011010110011111000100011000001110111111100000001000110010100000000011111011011110111010001010100000111100101100100;
#1 $display("%b", po);
# 1  pi=207'b100010100000010000100110101001001111001101001110011001110100001011101101000100111111101110010010111111001001000001000010101110001110000000010011111001011000001101110110010100000010010111010001010001110011100;
#1 $display("%b", po);
# 1  pi=207'b010001000110010010111010111111111100110010011010000100111011001110110010111101000000111111110010010110110001100010110010000100100100101000011111000010101111000110010000101001000101011011000000011111101110101;
#1 $display("%b", po);
# 1  pi=207'b011110010100010100111100111011001011111111010011100111001100011001110011000000101000110110100101010000000011000111011110011111100111011111101100111010110101100101011010000011011111010110100110010000001000011;
#1 $display("%b", po);
# 1  pi=207'b000100001100101111001101000101000011000100010011100000000111001100100010001000110011000100011110101001100011110011100101110011100001110100101010100011011001010010000101000011111100100000010001110100010010011;
#1 $display("%b", po);
# 1  pi=207'b110110010000000000101110000101100110000000001011010011111111010110001101011011111001111100100010100111000110001101010011111011011000100010000111001001011010011101010000010101010001001010101000100110101100100;
#1 $display("%b", po);
# 1  pi=207'b000011010000111001110101111111111100000000110110100110011001111100101111101011011101010000110011001100001101010001101001100100111001000110011110100000001000000011011001001110000100000100000000010000110011110;
#1 $display("%b", po);
# 1  pi=207'b010001010101100100010100111000001010111000010111101100101011000010111000110111001111100111000110110101011000110100000010001000000001010011111111110010010100110001011101100011001001011000001001111011111010001;
#1 $display("%b", po);
# 1  pi=207'b101101011111000001000001001111010110000110100000001100110000000010011101000100101101000101101010111010010101100100011110101111011100010011000100000011101011010001001110110110100001111011000011001110111111000;
#1 $display("%b", po);
# 1  pi=207'b110111110100110000100001101111000111011001111010111001110010011101011011100011100111011010011001011001111010010001101010110000110110110011101000110011011111100011101000101010000101111010010111011000111101100;
#1 $display("%b", po);
# 1  pi=207'b001011101100001010010001101000011101100111111011111001011011001111001111001001011001111000110001011011100100011111000010010110001110100100011010110000001001011111110000101001011101111101110100100010110110111;
#1 $display("%b", po);
# 1  pi=207'b111100101101111000011001101100100111101100010110110100000011001001011101110010010000011100001111011111011001100011010000000110101111010010011110011010101011101010111101111110000110010111110001110010101011110;
#1 $display("%b", po);
# 1  pi=207'b100111101001001111001100001010100101000101011110011101001001011101101011101111110101001011110001011011001001011001011010110100111111001100101011010001100000010011010110010101101101000110000000110001101000100;
#1 $display("%b", po);
# 1  pi=207'b011001100100101000011111110111111001110101010000110000111000000010001000011010100001001100011100000010100000000111011010001010000110010101000110000100001101001101100001100010100010010010000011000011000001010;
#1 $display("%b", po);
# 1  pi=207'b010111101011011001101000100110010011100001100000000001110111011111000100111111101000101111101110001010111101111101010110111001101001000110001001101011111101101110100100010011010111010000110110011000011000000;
#1 $display("%b", po);
# 1  pi=207'b111010000110011101010000011111010001000011001001100011110010100100000111110000111111000100011010011001100011100110101101100010101110101001000011011111010111001111101100101101000011000011010011101001100000000;
#1 $display("%b", po);
# 1  pi=207'b000100001000011000110110011000111101101000010010101110101110000000011000111010110100101011110010110100111110101111101010110100000100000010111000000010100100001011011100111001010010011111100100101101001001101;
#1 $display("%b", po);
# 1  pi=207'b000000001001000011100110100001001111010110111111001010001011111010110000011011001010000110010001001011100000101110011110001100100100010101101101010110110001000110000100010011101010111101001010011010101100110;
#1 $display("%b", po);
# 1  pi=207'b011011010001111000101101001101001110100111000000110011110010110010000101000111111110000111101010011001110101000110100101111001001100010110010100100000110100000110111101001100110101000111100111100110001101010;
#1 $display("%b", po);
# 1  pi=207'b001101001010000101110110001100111111101000111000011111010100100001101101010000100101110010000001010100111110010111011101001000111101100011101101111110011100110101001111001110000110011110101011110000010111110;
#1 $display("%b", po);
# 1  pi=207'b101001000001110000100101001001011001010110001111011100100110110010111101011101111000111011000100000101000001010001011010111100011010001000100000100000000000011000111011010100111000111100100000101110000110100;
#1 $display("%b", po);
# 1  pi=207'b010001010010110110100000111100101101011110111100111110010001111100010111101011100101110111100111101110101011100011011010111001110100010101110010110110111001000100101110110000000000011110110000001010101011001;
#1 $display("%b", po);
# 1  pi=207'b001110001001011010010100001010010010100010011001101001100110001111010110000110000100000100101110100010100001010000001001110001101000101010110010010000001000011100100101010011100100011010111100101011100110101;
#1 $display("%b", po);
# 1  pi=207'b010010000010110000010010001100100010001110000011111011000010100011011000001011010111100111011100111111001100110001010010111011111101000000010101101101000101111111001000110011011101001111000001110010011101110;
#1 $display("%b", po);
# 1  pi=207'b110001011101010001000011110100000010110000010101010011110001001101110111011011111011000100011001001100101101110000011111001111101110001111011011011110011110100110100101110001000000001011000010111111111111111;
#1 $display("%b", po);
# 1  pi=207'b100011111100111100110000001011000111101110100110001101101000010010010010111101110001101000101010100100000101010001000001011000001000000011100001101001111111000000111111000101011001100001000100010000101001100;
#1 $display("%b", po);
# 1  pi=207'b111100100000110000101010000011100010101001100110110000010111110111111001101000100011101110010010110111011101010111111110111100110000011110011101110011011010100101100010111010100000011111011010101010100011110;
#1 $display("%b", po);
# 1  pi=207'b101001010111110110001110001111100101001011111101000010001011111100110101100110001101110110110011011101101110001000101101110011100000100111000100100111010100110011101111011101100000111011001011001001110110101;
#1 $display("%b", po);
# 1  pi=207'b110010101101010010000110000010000011001001100100011111111110000010111110110100101101110001010000111111101000100001110111001011010001111000001000100001001000100010011110110110000110111000001011101001101110001;
#1 $display("%b", po);
# 1  pi=207'b101000110010000001011000001100001101101110010111011111100011111111011011100001101011011110111010111011001010100100111011001101001010101101000111011001001100101011001010011011001000100000010001010010100100000;
#1 $display("%b", po);
# 1  pi=207'b010111011101000001100100000110000001101001010010000010100101000010000001010110010001010011010010001000111011011001001001000011111101110011011000110001101111101001111101111001011111010111111111011101101000100;
#1 $display("%b", po);
# 1  pi=207'b101101110111001110010100010001000011111011111101100100100010100111100110100001100010010010101011111111100110111101100100011011111000010011000101100111001111100111110100000100110110011000111100110101100101011;
#1 $display("%b", po);
# 1  pi=207'b111110110000000011001101000000100100000001110100111101101000101110100111110011110011000110010110010000010010100101000110111011101100001000101111010101011010001100000111111100100111101001101001011001110111010;
#1 $display("%b", po);
# 1  pi=207'b000111110001100000110000001110011010111011100110110011111001111001011000001001011011001011000000010011101010101101101000110100110000000011000011001000111011101110110101011000110001100001011011101011100001000;
#1 $display("%b", po);
# 1  pi=207'b000101111101101011001010011110111000011001001000010010010101100110101000010100011101001110100111110001100111001101111011100101100111101101101100010001101101100100000101010011111011010110111011011110010111110;
#1 $display("%b", po);
# 1  pi=207'b110111110100100001001101110111010111011001100000111000010001110110010010000111011101011010000101100101110100100010101001110111101000011111001010100001000001010000111001000010111000111010100001000111100110100;
#1 $display("%b", po);
# 1  pi=207'b111110001010111000011110001000100110001100011000110000001100010010000011111110010001111000011111111000110101110000000110010010101101001101001111101011001001011110011101101001001110010010001011101110001000110;
#1 $display("%b", po);
# 1  pi=207'b011011001111111110101101011100100111011110001101010111010010011110000001101101010001110000001110111011101100001000101010100011010000010100110011100101001100100110100101000110110000100110111111100111000000000;
#1 $display("%b", po);
# 1  pi=207'b111011001011010000101001000000010001110011010110101100110000101001101110010000100000100101000011101101100100110101110001010010010100000100000011111110010101111111110011100000011011000100011010001100011000100;
#1 $display("%b", po);
# 1  pi=207'b001110100001100111100100000111001110010111110111001101111100111110001010100111111111010110100110111111011000000100110110101000111010100000110011100110000110011000101100101010000110011110011101100010110010101;
#1 $display("%b", po);
# 1  pi=207'b101000101011000011101100100100001001101100110010111000111101011001111101010110011111011001111011101010011101010101110010000000111001011101111100000000100001001100011111010100010110101100100111011100110111100;
#1 $display("%b", po);
# 1  pi=207'b100011111111111001111110010111011100101000000101011011101001111011000001101011111100111001011011010000010001110110101111000111110011000010011010100110001001100010110001100011111001000100100101111100010010111;
#1 $display("%b", po);
# 1  pi=207'b011000100011111111010000000011111000010111010110001111010111000110101011111001010010001010111110011100011111011011010010111101100000100100010110010010100111010111101000000110100001100011111111010100110111101;
#1 $display("%b", po);
# 1  pi=207'b010100100010100001010100010100010010011010010100000010001110101100010011101111100110011000011101111001011101010111011011011111010110001011010010100111011000001111101101001110111110011111000010010101001001001;
#1 $display("%b", po);
# 1  pi=207'b011000010111010101100001100101110100001001111100110101100110100110010011110101110010101110000111100011111111111111010111010011111111101000011101000101110101110001100010110101010101110110000111110100111000010;
#1 $display("%b", po);
# 1  pi=207'b011111000010111011101010110101101011011011100010010101110111100011000011111000000110100011010110100000001110010000011100100100000001110100000011010011110101111111001110011100101110011101010100111101111010010;
#1 $display("%b", po);
# 1  pi=207'b000000000010010111001001010001000000110001100100010011001011101110100001010100010010001011001001110111100110110110111001101001011011100100001001100111100111011000000100000011100001100011100001001110011011010;
#1 $display("%b", po);
# 1  pi=207'b001101010111100001000010111010000011010010100111001000001110111111001101001100101101010100101001111001011111010110111100100011100000111001100110001010000011011100101100000011000000110000101010001101111110000;
#1 $display("%b", po);
# 1  pi=207'b110110000101100100011011011111001011010101000010000001000101110101010010001100101101010011000010110101111110100110010001001110111010101110100001100100111111010011101110110111000100111111110010101000101100001;
#1 $display("%b", po);
# 1  pi=207'b010010000110010000100111101011010110100001000010101100001100110101111101011001101001111011110000110110000011111101000011011110011000001111110111100101011101110000100110110110000011011000100011011011000111110;
#1 $display("%b", po);
# 1  pi=207'b110101110111000110010011011000111011010010010111011000110101011111111111000111001111001011011110110110101100100001011110111011101101101001001001001111110100100111101100000100000100100001010001100011101010001;
#1 $display("%b", po);
# 1  pi=207'b101100111001011111010000000111110111011011011001000100000100111000101000001011010100010111001011000000000000001100100110001001001011111101010010000110111100000001010101011110000010010100010100100000111010010;
#1 $display("%b", po);
# 1  pi=207'b100001011011001110111100110010001000101011100110000110101100010101001001101000111001101011111100111000101100010111101110110000010011101010010110110000101010111011001011101000011010110111110111010011100100011;
#1 $display("%b", po);
# 1  pi=207'b000111111101100011100011000001001111101001001010110011000100010000011111010101111001100010100100100010110010000100010010000100001011010110110001101010111101000010000011110001001110011111101111000001100100110;
#1 $display("%b", po);
# 1  pi=207'b110001000111010000000110001110000011000110010111010001010110000100011101101010011110100111010111001000101110111010001000001011111011101000100100011101001010101111100101100111101100001011001000010100000100011;
#1 $display("%b", po);
# 1  pi=207'b101111100111001111100010111011110111101110101001110100010001111101101101111000111011111000110111000100001110000100011001010011100000101110100010100101101000000110000000111001101101011010111101011011101001110;
#1 $display("%b", po);
# 1  pi=207'b111011111110110011010000100101110011001000011100011110101000011101000000010101100010000011000100010100111011101011111010111010100101111011011010111011010110101100110011010110000101110010011000110110001111110;
#1 $display("%b", po);
# 1  pi=207'b000010100100001000101110100100101001000111011000111101111000111010001011101001001110101101000111000010100010001010100011010101111111100101010111000110000000001011100111011010101000001100011000011000000100010;
#1 $display("%b", po);
# 1  pi=207'b111110001111110110111010110110010110000010010010111001111101010010000001111010001100010010000100101110111100000000100101001101011011111111111101001110011111010101011100000001011011111011111100010110111001000;
#1 $display("%b", po);
# 1  pi=207'b011101011010111000011010001110011010000111110110011010010101101010101100110001000010100110010001010101000101101010100011111110001101001101010001110110001000101001111100110001110010110001001100011010010111010;
#1 $display("%b", po);
# 1  pi=207'b100011010110011000011100110101011110011010000000100001100011100010110111101100110010101101010100000010010000100011011011000010011001101111101001101111010110001011110100011010000100111011101101001000111011011;
#1 $display("%b", po);
# 1  pi=207'b111111011010111001010100001110010111011011100100111000010101100100000111011111000111001010000011011100110100000101111110010000011001010111010000010010101000111101100101010000001010000011100100110010111001100;
#1 $display("%b", po);
# 1  pi=207'b011111110101101010100110101100001001000111111000001010101101111110001111001010000101001101110010000010010110000100010111011111010101001111001000100100101111011001011100000011010001110111001100100110110001010;
#1 $display("%b", po);
# 1  pi=207'b000011010111101000110110001000011000010000100111001100000010011000010101110010101011000001110001101111100100000100100110001000011000111010010100111011011110011000001100101011001000000001101101010010001100000;
#1 $display("%b", po);
# 1  pi=207'b111010011100101111011010100010110011110101101101001111111000000000100100100101011101000101111100111110000100010001111101110001010101101000001001000010110001011000001001110000011111101100110000011001011011100;
#1 $display("%b", po);
# 1  pi=207'b111100100110010010101010101110100100100100110001000100001011101111100001111011111101111011101010110111110101010011011101110000010000010011100110100110001111010111000100101110101001110010110000101000100010001;
#1 $display("%b", po);
# 1  pi=207'b110000001110011010111110001110010011110111101101101110110000011001101000101010000101000001000100111001100010100100110111010001111011000011000011010110010001000110111111111110001101111100001110110101111101000;
#1 $display("%b", po);
# 1  pi=207'b100110111011001010100110110100100001010011011011000000010111000110111101110010110111011011001111010000000111011101100010101100001000010110111000100011101000010010111100111100000110011100011011001010000111111;
#1 $display("%b", po);
# 1  pi=207'b110101101110001011000010100001101011011101000010110100010010111011100011000110111011001111110001000000000001111101110011100111110000010111110010110001010100001011000011101000101111110010010110110010111111011;
#1 $display("%b", po);
# 1  pi=207'b101000000111111110001000111001010001100101111011100101101101101100001100101110011111111111110001010001110110110001011001101110001100000000101010101111011100110000111010101011010001000010011010000111011000000;
#1 $display("%b", po);
# 1  pi=207'b001101001100101111101000111001111100100010010000011110100110001110000010100111111010100010001010011001011010010101011111101001010110010110010110101000010001110110000011011100011001001001011000010101100100100;
#1 $display("%b", po);
# 1  pi=207'b011000000111111011001000101100110011111011011110101111001011000101111011011001000100101110101110101000010011110110001000010000111000110001111000001100011010110001111000111101011001110110111011111000101011011;
#1 $display("%b", po);
# 1  pi=207'b010110111010000100010010001011000111001000000100110111001010001100110001101101111000111000100000001011111010100001001110000000011111010100011110001101001100011010101100000110100010001101000011011110100110101;
#1 $display("%b", po);
# 1  pi=207'b010010001000001101000001101101011111011000001000010011110011011110110001110111111001101111111111100100000011001010000010111111100011100010111110001010111110111100001101011110101001000100100000111110101000011;
#1 $display("%b", po);
# 1  pi=207'b101000111010001001100100011000000101100001011110111100010101010010110000111001100111000110111101111111111011111011101010111101001000000100111101111011011011101001011100001101111000100111100001011010010101011;
#1 $display("%b", po);
# 1  pi=207'b001101010010011100000000011011011001110110010110011011000101101001000000000010111100011000010100100000000000101010011001000111100111100000010111001001111010110000000110011010011100000011111010111011011000011;
#1 $display("%b", po);
# 1  pi=207'b101000101110010111011000110010010101001100011001010011111001001100001010111100011011111101001011101011111010000111000110111100111001001101010000011010101010100011101110111011001110011000111110100000110011001;
#1 $display("%b", po);
# 1  pi=207'b000001111011010110001010001001010101110110100111111001010010011111111011111110110100001101101101010110000001110000100010101101001001100010011111111011010110011101010100001000000111011010100011110010010100010;
#1 $display("%b", po);
# 1  pi=207'b010101000000001101111101101101001011110110110111111110000100101010100001001101111010010101101100101110100110100010000100101101000011101011010000111011001000011101001111000111111101011110101011111100100100011;
#1 $display("%b", po);
# 1  pi=207'b000101001101110000101001010010010100111010001010111010000001110001111010100100011010101000111001010110010110110010011111110011000111101000100100111101111100011111001000110101001010000101111011100010001101100;
#1 $display("%b", po);
# 1  pi=207'b001000111100101100001000100010010101100011110010101011100110000111111110010111110111111000000011101001010010100111100111111110110011000101001100100000011101101111100111100101000011000101011000000001010010010;
#1 $display("%b", po);
# 1  pi=207'b000110110001111001101100000000110001110110000110111111101011110111110110000110110101110011000111000110000111110100111011111111101101111011010001101101100000001001101011101110110010111000100110011001111110101;
#1 $display("%b", po);
# 1  pi=207'b100111110011011100000001111011100000000101010110000001100010110011100011111000101011100100110111111010000001111110011101100101111011100110010001000111001111111100101111110010011101101000100101111010110100110;
#1 $display("%b", po);
# 1  pi=207'b000000000010100011101110111110000001110100001100110111011111101011001001100000100001100101010110101001011011100001000010100000111000101001000111011100100010000100001101001001100100100001101000111011010010001;
#1 $display("%b", po);
# 1  pi=207'b010101100001010111001111000101110001001110111010011011100010001001001110101010111010001010011011000110011010100110101101100010010011001011001110000101111011111010111100010100100101011110101110001100110011101;
#1 $display("%b", po);
# 1  pi=207'b010010011010110111010001110110110101100111111101010100110100101100000100011101011111111001011001001010100001000111001000110111001010001110010100011010001001000100111011110010111001010010000110110100111011110;
#1 $display("%b", po);
# 1  pi=207'b011111001011100000001101111011110110000101011010100001001110001000000111100011101111101111101011100010101100011011100011110110001000110001111011010000100110110000100111100111010001110010100001100010100100100;
#1 $display("%b", po);
# 1  pi=207'b100011010000101101101110001111010011010001010101011001010000001001101010111111101101001000100011100111011011010010100100110010000111110100101101101111110110110001010100100001111100100110100101001101100001001;
#1 $display("%b", po);
# 1  pi=207'b001100011011101010000001010001101010001110001000000100011110001000110001000000111110110001001010110101110101100111101110111101000100100101101011010101011110110011010000010110100100101011101101010001111001101;
#1 $display("%b", po);
# 1  pi=207'b011100000001101111010000100111111111101001011000111010100101011111010011000100001110010000110001010100000000010000110100000101111000000011000000111101100100001101010001001110000101101010001101110110010110110;
#1 $display("%b", po);
# 1  pi=207'b111010000101110111010110111101100010111101110010010010000110010000100010100011101110001001001101001101101110011001101010011111110011110111011101110001001100010011111010011100010011010100101111010100110011001;
#1 $display("%b", po);
# 1  pi=207'b011100110101110011010001010001001001101001111110011101000111111001110111110111111011101000111111101001001101000001000000000100010000101000101000111001101010100110011110010100100110100010110001011010001101110;
#1 $display("%b", po);
# 1  pi=207'b111011010100011001001010010110011100110001101100001101010011000100011111001100100110100111111001100111011110010001001001111110110111110110000111101010001011001011101011001011001111111001101111101010110000111;
#1 $display("%b", po);
# 1  pi=207'b000101111100101110000100011000100111101100110010001011100001001010100101011001011010110010101100000000100000000111000011000101111001110010100010011011110110011010110010100110101100111001000111011010001011110;
#1 $display("%b", po);
# 1  pi=207'b011000011000110001010001000110000110111001000001001100101100110100010100001010101011001010101101101101011000010100100101001100000100010000001111000010100111100110010101010101101010011011011010111100110000001;
#1 $display("%b", po);
# 1  pi=207'b100100000100110110101100101001101100111011100001101111101100011111001010001100101010011110000011000100100000111110100100011000111011111111000100111111011110101000101100110000000100010000101111011000111010011;
#1 $display("%b", po);
# 1  pi=207'b100010110001010101101010011001001101110100010111100010011101000100010101001100011010010101100001111000010111000100111100100100101110010000100011100000110011111110111010011011100100111110111111011001110101011;
#1 $display("%b", po);
# 1  pi=207'b010010100110010000010001000011010101111000010111001001001011011110100000100110001001101000100100001000101101111100000111101001010011110010100000111000101000010010100101110111001100011101101111100111011000010;
#1 $display("%b", po);
# 1  pi=207'b111111010110000101101100010111111111100111110011001010010100011010110100110111101011110110011101011011011100111011001010100010111001111011010011100000111101010100100000111110100101010001111110011111111101110;
#1 $display("%b", po);
# 1  pi=207'b111111011101101101100010100010011000011000010101110101110111010110000011010001010100111100010001010011010011010111110011011111001110010111001100000001101011001001111111101010011101100000100100010001000011110;
#1 $display("%b", po);
# 1  pi=207'b010011000010101101100100100110110110001110001111111010011100111010010000000110100100010110101001111001010111001110010011100100000000010000010010100101100101000010001111111010100111101001011110010110001100010;
#1 $display("%b", po);
# 1  pi=207'b100001111010011100100100111100101000001000001111011101010001110010110010011010100101101111000110111101001000011111011101111110000101011111100010001100011101111010101101001101100000101111010111101001111110010;
#1 $display("%b", po);
# 1  pi=207'b111100110101011101011110000001000110101000110111110101101001010001001101010011100000110110001011010001010101000100111001101000010000100010001011011101001011000110000111111010111100111011010001000000101010100;
#1 $display("%b", po);
# 1  pi=207'b010100011111100101011110011111010111100110011010101101011111111101110000100010111111000000011010111110011011001110010111001011011000011111111010010100110100011111110001001000001011100100100001101011110010110;
#1 $display("%b", po);
# 1  pi=207'b100100000100010101010011100011111101011000001000010100110000111110101111101111000000000110000100011001111110111010110100000010010110010101100100010111010001110001100101011011010111111010001110100000001000110;
#1 $display("%b", po);
# 1  pi=207'b110010100000111110101111101110110111111011101110100001111001011101111111101101101101000000111010011111001110000001101110100011110110101100011110010001000100000011000110000110110000001001011001011010101100000;
#1 $display("%b", po);
# 1  pi=207'b101111000110111111100001101100100110010011101010010101010011111111110010011000010110011101001000001001001100111011100110111101001111101110011011001001100100110010100110101101011110110101110001100001011101101;
#1 $display("%b", po);
# 1  pi=207'b001100100110011100010111101001010111110011111000110101011010111011100100000011001100010101110000100101001010111111011111101101000001101000110110001001010000101001010001110010110001100110001001011001001100100;
#1 $display("%b", po);
# 1  pi=207'b101101000000100101000000001000001100101101001100000001110101000111001101001000000001011110001001111011111011010000101110101011000001001011100000101111100110010101001110000100101010010100000010001101111000001;
#1 $display("%b", po);
# 1  pi=207'b110010011101000000000001101000101110100101111010101111010101101001100101011000011110111011010010010011100110111011100111111011010101110110110000000110110110111001011011100000001000000011101000001110001011110;
#1 $display("%b", po);
# 1  pi=207'b000101111100110101110010010000010001000110011010001010001101101110001011000111011010110000001000001100111101001111101110110011011100001010100111110001010010110101101000111100001001010101000011100110100110111;
#1 $display("%b", po);
# 1  pi=207'b001001010111001000000011001011001001010000010001101110001000001010010010111011010000100101000101111111100101100100110001001000111100010100011111001110110000101101100000100110011000001100000101001010111110101;
#1 $display("%b", po);
# 1  pi=207'b101111110001100111011010001010111101100001111000000100110011000001011110100111001100011111000110101110101010101001110110000000010111001000111101111010111010110100110011001010111100111101100110111101111000111;
#1 $display("%b", po);
# 1  pi=207'b011100100000111011101111100010001001000111010111001101110011111010010000011101001101111111111001011101101011001101010100001000011101111001010111001011111111111110100100111001110001110111011101110011010101101;
#1 $display("%b", po);
# 1  pi=207'b010101111110000001100101111010101010100000100101000011100100101100011110000100110001011000100111001100010101001010001100001011011010111110111010001100011100100100011011100001100011100101011000000110101110111;
#1 $display("%b", po);
# 1  pi=207'b010101110011101001111010111111010101010100100101011110111000110111000010100001001111001011001111000111101111011010001000111000111001111110100101011001010011101010111101001110010100010100001001101100111001101;
#1 $display("%b", po);
# 1  pi=207'b011110101101000110000010001111100000011110010010000001101101111001110100001000110010011010101000110010011001010001111101000001100000001001110111111101010000110100001010000001111000000010010000110110001000101;
#1 $display("%b", po);
# 1  pi=207'b001110101100001111101000110111001111010101101000110100101110000101011111110010111100001101110111010000011011100000010110101010001011101011001111000001001001001111100101010111001110110110101101110001000000101;
#1 $display("%b", po);
# 1  pi=207'b010010100100101110011000000001011101100000110000000001000111000111010111000100010111010110010000110001100010110111101100100010000000010101111011001000010111101100000010011101001010011111001010000001010011101;
#1 $display("%b", po);
# 1  pi=207'b111010010110110011101110111000110101010101011111111000011010110011110111101000000111010100011111100010011110001110101000100101101011100110010111100101110101101000110011000111111000001010001011110011111100111;
#1 $display("%b", po);
# 1  pi=207'b011110011111010000000010000010110111100011110000111100111111110000110001001111000100110010011111100111110110111000110101011110100100010100011000111100110111001001111001001011111001100110001101110011011001010;
#1 $display("%b", po);
# 1  pi=207'b111001111000101110110111011001110101111010010110101100010111011000100010001001001100011001000101010100010100110000101011111000110001001011011001000111010000011000111100111101110101010000100010010111010011110;
#1 $display("%b", po);
# 1  pi=207'b110111100001111011111001100011110001100100101100100001000100000001011010010100010011110111110110010000111010001100010110011101100001111101011011010101111000010110110011011000111010101011011001110010001110001;
#1 $display("%b", po);
# 1  pi=207'b010001001110011111001000111010000100100111101011000110011101111011110101100001001110110000101110011001110010101110101110000000101011110011001100001011011111000111100001110101010011010010010010001101011000101;
#1 $display("%b", po);
# 1  pi=207'b101011110111000111101011010110111100001001010111110111000100011011100101010101000000101111001010000110000000010011001101111010111111110000101101011011101100001100010001110011101001110110001101110100100110100;
#1 $display("%b", po);
# 1  pi=207'b111000010101101111110100011101101001011111110100010010010110100011010001011110111010111100010101000000011110011101101110011101010000111111111100011111000100001001100110010010110011101110101111000000111101110;
#1 $display("%b", po);
# 1  pi=207'b110010111111000010110000010001001110100110111101010110110010101011000110010110101101010001101001000111010111011001010011100010001100011000011101011011011000101111110011111110000111010111100110010101011111001;
#1 $display("%b", po);
# 1  pi=207'b111101000110100111101110011001111110010100111100000000000010010000111111100000011010110110101001101111010110101000011110011101100010110010110111111111111101110111010000101101111100011011011001110100110110011;
#1 $display("%b", po);
# 1  pi=207'b100001011011111101100100100110101011001000110101101001101011010001011111000111101100001101000111110100101010011100010000011111010000110011110100011001011110001100101001100110110000110010100101101110110111101;
#1 $display("%b", po);
# 1  pi=207'b001100100010101101111010101110110110110011011000011111010101010101010111111101001100001000110110011011001001000100111100110011101011100101011010111010111100100110100100111110010101101110010100111001001010011;
#1 $display("%b", po);
# 1  pi=207'b011111110101000100110011110101011101100010100110011010010101011101011001011011001110001111100111010100011111100010000100111111101111001001011110011111001110001011011110110000010100100101100111101101000000111;
#1 $display("%b", po);
# 1  pi=207'b110111110001011000101101111110010010100001101101000110001001010001010010010000011110001101110011111010011000100000000011001101100100101011010110101001001100011100100110110111000100011101001111010100111000110;
#1 $display("%b", po);
# 1  pi=207'b101111110000001101110011111110011001000011001101011010001110110000000011111101101100000000000101110100001000100000110101100011111110010000011111110001010010010000110111001110111111010001111001010011001111000;
#1 $display("%b", po);
# 1  pi=207'b111110010111101010001110101011110011001110010010110001010001000001011011110000010001010101110010111010110000101101000110111111100011011110000001110011001000110010111111001000111111110100100111000000010010100;
#1 $display("%b", po);
# 1  pi=207'b011100011101100100111101000101011000100100011011111010001100001100101011001100101000001000100101101001001100110000101111010111001101100011101101000111101011000101101010110101101010001111000110010111010010010;
#1 $display("%b", po);
# 1  pi=207'b001001001001110001010110001100110010011011011111011100011011110001100011111101101101000111001011101111111110010111011001110111010100010111100101011111110000100110100010000100111011010001111001111011000011000;
#1 $display("%b", po);
# 1  pi=207'b001111001010110110110100010100001000000001011001110111001011000110101101111110001101100010110101000111001100010011001000011101111010000100011101011000100001011010111100000110010111011110111011110010100101100;
#1 $display("%b", po);
# 1  pi=207'b110000100010000000001000001011111010001011101000000100011010011001111000000001011011101011001010001100001100111011110011010101001111110010100001000100011110111111111000101011000011100101100110101101101111101;
#1 $display("%b", po);
# 1  pi=207'b011101000110010010111011011010101111011100111001001101100000110000001000100101111010101101111001111011101101011001000011000011111110111100011000011010001100011010011111001101011111111100010001010101000111110;
#1 $display("%b", po);
# 1  pi=207'b100011100000000111101111101111010001001111001110100100000111111001001011001001010000000001001110111110111010011000001100011111010111011011010011111010011110101001100000111110110001011011000110100100110111011;
#1 $display("%b", po);
# 1  pi=207'b010100110100001111100101001000111100111111101110010011011111011000001111001111000111110111001011110011100111101111110101011101110011001000110100011000000100011100101001101110101000110001001111011111111101111;
#1 $display("%b", po);
# 1  pi=207'b100101011001110011111011000010001010110000100011110000110111111000010011010100011111001010011000000010011101011111101101000111100011110111001100100010110111101100110000110000110000110111111101111100111000001;
#1 $display("%b", po);
# 1  pi=207'b111010001100011011101010001010001001111001010010001101010101100011110100100110110000101110111000111110100001111000000100110100110100011001011101011101011100011011100101111101101000111001010110111000111011010;
#1 $display("%b", po);
# 1  pi=207'b110100000010100110001101111011110110001100011011000001001000101101001001001101111010110110101010011101110010000001010011000000001001011010000100110000010011011010110111001010111111000100111010001010010110000;
#1 $display("%b", po);
# 1  pi=207'b000001110010111001101001111000000111010110001110011011001011000110000111101001101110011101010101100011111110101101001101001100010001011001011001100011111101100101011101110010001101011010101100111011111110011;
#1 $display("%b", po);
# 1  pi=207'b100101101010100011010110111111010010001111100011110000101000001010000010000000010101000111010100001111001011101011001011001111101111101101000101011000001011010001110010010011010001110010100111010010001111011;
#1 $display("%b", po);
# 1  pi=207'b000010011100100110110111000100101010111100000111111101000001010111010010100110011011100110111010000100011100000100111111111110101010100010110011101010100110100001011010100111000101000100001001100011110011011;
#1 $display("%b", po);
# 1  pi=207'b111011001010100000101101111101000111110010110100110111111010011011001111111001110111110011001001011100101100101111010011111010101001101010001110000000010111011010111000110111011111011000010011001000010101010;
#1 $display("%b", po);
# 1  pi=207'b100011011011000101111111110001010101011011101100010001110001101001010001001100001110111111000100111101101001111101000010001010011101000011001000000010110010001010101111110100011100010011100111001111011000101;
#1 $display("%b", po);
# 1  pi=207'b011001101111101111111100101010010111100111011001011010001000100010111010110010101101011011010001100100100111100110100101100001101011101100100110001100111100100011011010110000100111111000100110110000100001110;
#1 $display("%b", po);
# 1  pi=207'b010101010011010111110101001100110011001100110111100000110101100101100001110100101000111111001100100111000010011101100101100010000110000010111001101110011011010011010010001001101001100001010100001100010000100;
#1 $display("%b", po);
# 1  pi=207'b100000100111011111011111101101100111010111000000101111011011000101100111000000000001100010101010000010010001011001101111100100111110011100001110111011010111101011011001111010000111100011101101000101000000000;
#1 $display("%b", po);
# 1  pi=207'b100100111010100011010110000011111000101101011011110010001011000100101100101101111101010100011111100100011110110010000110111010010111011110010001100000110110010101110110111011110100000000100000001100001011111;
#1 $display("%b", po);
# 1  pi=207'b001010100001100111001100000100000101110010001110100110010110111110100000101101110110010010011011011000101100110010001100010010001010011100001101010111111010001110111011001001010000001100101010110011110100110;
#1 $display("%b", po);
# 1  pi=207'b111111011110100000011101100011111100111101111100100011110110101110000011101000001010000101010011111100001100011010101111010110111111110001101111001110000111101010001111100000100010110000110111100000001100001;
#1 $display("%b", po);
# 1  pi=207'b001001101001011000000101110110010000100101001010101001100111100111110000110111110010000111010101100100010010100000010000011100111011100111110110110110110010001111101001101000101010111001010111011001111110101;
#1 $display("%b", po);
# 1  pi=207'b011010001011101101111100101001101101101010111111110100010101101010000000011100100011101100111110111001001110100011100101000101101110110111001110010110100001110110010011111011000000111101000111001111001100010;
#1 $display("%b", po);
# 1  pi=207'b100111010011010001100101010100101111100010010100000100100001111111001100001110100010100011010001100101001101001111010011111010101011010000111001001011001001110111001111101110000010101101101001010011100100011;
#1 $display("%b", po);
# 1  pi=207'b010011100110010110111111011101101110110101101000110111110100011110111011101110011001011111000101000111111011110111100000000101100010110100010110001111001011001101100011010101010000010011111111101001110000010;
#1 $display("%b", po);
# 1  pi=207'b011100001000100101111100111000011010010001100010000110110000101100101001110000110111001110000001000010100110010101001001111110001110011000011010010001000111010110100101111110111000010111001101101100011101101;
#1 $display("%b", po);
# 1  pi=207'b101111101010100010101100111010100001100101011011001101111000101000000010000111100101010001001011001000101001001101100101101000100010111110101111000011110111100000111010101111001010010010101001001110100011011;
#1 $display("%b", po);
# 1  pi=207'b101110010111000010110011100010100110100001011100000100000001011100111100110011001111000101011100001011011110101011011001011000111010000100011100111011101011110000100110111011011101001010110100000110000001001;
#1 $display("%b", po);
# 1  pi=207'b011000111110110111100101010111101010000000000001111100010010010000111110011100001101110001100110111001010111110101000111000000111111001101000001010100100101110011011010010110101011100010010100100100110000010;
#1 $display("%b", po);
# 1  pi=207'b101110111100101101001101010101011001111101000011111001011010111100101100000111001011110010000101100010111111001011010110000000110010101111001111010111011001100101101001101011010001110101000000111100011000100;
#1 $display("%b", po);
# 1  pi=207'b110100110000110110111011001001100001001000001101011010000010111111011010001010101010110100010010110101000001100001100000011100000001111011100010011100001100001001110001100000100011000000000110010000000110011;
#1 $display("%b", po);
# 1  pi=207'b000001000011110011010100110101011010111010010000001001111011011110011100111111101111101000100101011010000001100110000110000011000110000000011110011101010010000101111011101111101011010011100100001000001100110;
#1 $display("%b", po);
# 1  pi=207'b111010100100111001110101010110000010101000100110100111010111010010101100100010001010101111000001010011110110101100010001110100101011000110101101111111000110001100010000001001100100011111111101100001110100011;
#1 $display("%b", po);
# 1  pi=207'b101000100000001111110010110110011110100001000001000000111101010011010101111001010101010001010011111010111011111001000100101100100010101011101001011100001001000100101101010001000000101001010110111111111010011;
#1 $display("%b", po);
# 1  pi=207'b000111111010111100011110011101111010101111011101111101100111000001110011001100110110010111011101111000000111111011000111000000101101110001011101110011010001001110001101111011110010111110101001010011001011000;
#1 $display("%b", po);
# 1  pi=207'b010100001111001000100010010011010111000101110011000101010101001111010100010101001110110111100101001000110100110010001000110111001100011111011101111100110110011010001010111000111001000011001100010010110110011;
#1 $display("%b", po);
# 1  pi=207'b110001011001010011010100100010011011001110111001100101000101110110000011010111011010000001010000101100010001001101011000010111101100101000010001000011100010010111110010011000001010101010011000011001111111010;
#1 $display("%b", po);
# 1  pi=207'b101000111000110101000001111100110111101100100100110111111000101011000110001101011110111011011110010111001011101010100100010011011001111100010111110111010010000100010100110101011010011101110100111011010011011;
#1 $display("%b", po);
# 1  pi=207'b000111011100110000101110101001011101011011111001001011000001110001110110001010000100010110100001011011001101010000001000000110010101100001100100000001101110100100101101111101000101110011111000011010000101100;
#1 $display("%b", po);
# 1  pi=207'b110011100011001010011111010101011001001110010100010101111010001110101110100010010100000001110010000100011000000000000111001010000100100110000100011000101100010110001100000001001110100100010001100100101001110;
#1 $display("%b", po);
# 1  pi=207'b100110001111010001001111110101101110011011110010100011101100101010001110011001101011001001011110101010100011000010011101011100000011111111001101001111000010000010101001111011011000101111101110111110110000111;
#1 $display("%b", po);
# 1  pi=207'b001100001010101110101101111001001101000100101111101000011100111010100000000000000000011001110010000000011111111110100010101110111010111101111010111000100111010100010001110100101001100000000000110010100101111;
#1 $display("%b", po);
# 1  pi=207'b101000010000001110111101010100000101011101110010001100011111000001011000100110110101011000100000011000111010100111110100010101000001011001101011111010101111010010101001111110110010101110001110110010100100100;
#1 $display("%b", po);
# 1  pi=207'b111111101011010001011110010010011000001011010001001101000100000100001000000011111000111010011001100101010110000011110110000001001101011101001101000100000001011001111010000101110110010010100111101101000110010;
#1 $display("%b", po);
# 1  pi=207'b001110011110001111111101010010001011111000010000001010100011011110001011101010011110011111100100000000000011111011001111011010110110100111101110001101000010111111101011010110111001011110001000100101111011101;
#1 $display("%b", po);
# 1  pi=207'b001101011110010111001001110101110001010000000000010011010111000000010001001111000110111010101110011001110010011110000011001101101100010011011110111000010111110110001001111110111001101101101100100100100111011;
#1 $display("%b", po);
# 1  pi=207'b000101000100011110111110011010110000111001011101110111111011001011111000000111111101100011011111100000010101010010001100010111011100100111111011110010111110101000111000110011111000110100000101101001011011011;
#1 $display("%b", po);
# 1  pi=207'b010010100000000100001100000010100011101000100101001011111110001100110010110101110101011010111001110101101001101110001110100011100111010110011100000001101101111010101101001100101100111000011001110111101110110;
#1 $display("%b", po);
# 1  pi=207'b001000011011111000010110110100010001110010010110011101001100111001010001010100100100110111111011110000111101110000010011001111010100000101111001111100011010011111000110000011110110100001100001011110101000011;
#1 $display("%b", po);
# 1  pi=207'b110111100011100111100110011000001100011110110100110011010111111101110001101001000001001010011100001111100011011110101100001011010000011101110111010011010111000011111001100010000000001000100110100000001000000;
#1 $display("%b", po);
# 1  pi=207'b010001100100101010101101111100001100111011100100001010101001001111100110110011111011001011110010000100010111110010010100010110111001001111000100010101001010001100101001001000011011111011100011001011001011111;
#1 $display("%b", po);
# 1  pi=207'b010000110100111001001001101011101111111101010000111010001000110100010110011001010000101101100110000001000001111100011001110101011110000100101100001100110001010100101111101111111100000100011101010001101110101;
#1 $display("%b", po);
# 1  pi=207'b101001011100011100010100111011110000111110110111010100111111001100110101011100000111111111001010001001110010100101111110011000111110010100100010000101101001000110100101111000101010000101000101010001010001100;
#1 $display("%b", po);
# 1  pi=207'b011001001000100101011111011011001101010101000100110001010111011000011001001111100110011111011001111100011010000100001010101100111010001000010111111100001000001010001100010110110011100011101000100001101000010;
#1 $display("%b", po);
# 1  pi=207'b011101110100010001100101100101000000100100110100101000111110000001001000110001101100001111100001101100001100100100111011100011111110011110101100011010110110011001101011010111100010001010110001010110011010010;
#1 $display("%b", po);
# 1  pi=207'b010111010100110110100000110101000010001000111110111001000110001011100011111001111010111010000011011110110111110110001000000100111100001001010101101011111000111001110110011101011010011001101100100100110110001;
#1 $display("%b", po);
# 1  pi=207'b111100110000000111000100110001000010001100001000010100110011001101100000111111100010001110101000000111011010110100011110000011011000100111101100010010000101111100010011001010101011010010110100011101000001010;
#1 $display("%b", po);
# 1  pi=207'b010011010101110000010011000110001001101110011010110111110110100001000000100101000100111100100001000111111000000010011000000101101110000101010100100000000011001101000000101001010001110001111010100010010000000;
#1 $display("%b", po);
# 1  pi=207'b000100011101011110001000001001011001000001001110001011001000101001001111110010110000010011000110000001110010001000111011011101010001001111000011111100011000001111010010101010010001001101100000010001011011011;
#1 $display("%b", po);
# 1  pi=207'b100010100010110001100110000110011111110001000110000010110110000011101000011000010011010111100000111011010011110110101000000101111110010110110111010010001100100100110100011110110100001010001111000001111000111;
#1 $display("%b", po);
# 1  pi=207'b001111110111111001101101000100100110101011110001100001001110010011001101011101010101010011110000101000101000001001100101010100011111001100110001101110110101010111000110001100010001101000001010001001001101101;
#1 $display("%b", po);
# 1  pi=207'b110110011001101010001011010111101101101111111000010001001000111001011010010001110010010010100010101001110010111000001110101010000000100101000011010001100011111011101101010110110100101001111110000101111100000;
#1 $display("%b", po);
# 1  pi=207'b001101111111111011101010111110001010001110010010110101110010111100111100101010100000000101110000000111001111011001001001110100100110111111001111011001000101011111010001110111101001101000100010010100000110001;
#1 $display("%b", po);
# 1  pi=207'b101000111000101000001100100100100101110111110010100111010101100100111101110100110101111111000100010000100111111110001000110100111110001010100000001111001101110000011111011001100011101001011010111111011100000;
#1 $display("%b", po);
# 1  pi=207'b001110000001001001110010100010111111000000100001110000001100100011011111001111001100101001110101010010011110010010110000011010110011010111011011001111110000000000111011100001101000101011100000110001100111010;
#1 $display("%b", po);
# 1  pi=207'b010000011010001101100111011010100010011001010101110111010000110111011111111011001110011110111011110100101001000000101100101000011011001001110000001101111111111101111010010111010010011110111010010110010000101;
#1 $display("%b", po);
# 1  pi=207'b101110110111100001111000110110010011011110111100110010110010111100011100000111001010001010100011001101010101001011001111101000101101011101101110010000110100101000000010101011111111000101111010000100111100000;
#1 $display("%b", po);
# 1  pi=207'b010000101111010001011110110101000110010101001000100110000010101100000110111101011011001111011001111100000101010010101000010010010011000010000011110100001010010011000001000000100110101100110001001100100001001;
#1 $display("%b", po);
# 1  pi=207'b110110010001000111110001010011110001000010111010000011111110011100011110010110101100010011101111001010101111011001000101110110010011000000100011100011011101100000010000101100100011011000000101101010001110011;
#1 $display("%b", po);
# 1  pi=207'b101010011101010111010110010110001001110101001101100100101000010101111110011001100011011110101001011111111111010100110111110111010001001011010101100111101111100110010000011001010110100101110100100101110110110;
#1 $display("%b", po);
# 1  pi=207'b101011101101001000111000100010110000100110011001010011100011010011111100110100110010101000100111010100100011111000111111111100110000100000000101000101110001000000010101010100110011110011100101011010100100100;
#1 $display("%b", po);
# 1  pi=207'b101000111001101011100011101111010110100110001010011000011000001011001001100001101111001010011010111010010111111000110010010110101110011110011111001100001010101001100011100010100010011001000111000011110100110;
#1 $display("%b", po);
# 1  pi=207'b100001011000111100011100010011101000110000001100110100011110101100111110111101110010000110000000000100110100110001011110100100001011101011011111011001000111000110011101010011000101000111010000111111111111110;
#1 $display("%b", po);
# 1  pi=207'b111101010011001010100011011010001100010111100001000001011100001011100111010001110111101000110001110011100111000010110101010010010001000010110001100111001110111011010110111100110101011000011100101010000111110;
#1 $display("%b", po);
# 1  pi=207'b111111100101001010010000101011100011110110000101110110010100111100011110110001011101001111001001110101001001001011011001101111001110001000011001000001011001000001001100100100001001101101110110001001100111001;
#1 $display("%b", po);
# 1  pi=207'b011011011101010100001110110110110101011111010110000011100101001001100010100001111111100001011011101111000110101001111111111011000101101000010100101101011111000011100100010101011111011000110101111110011001100;
#1 $display("%b", po);
# 1  pi=207'b100000110010000011001111110110101101110000010000101001100001011010010110011010010010010000000010110011111010011010100001101111110000101001111101010011101001100101100110000110010001110000011000101100001010011;
#1 $display("%b", po);
# 1  pi=207'b101111011000101101000101100110100101010100001001011000101001001000010110111011111111101000010101100110001111011000011011111110101001001011011011101011000111100111000000100101001101010111010100101101011100111;
#1 $display("%b", po);
# 1  pi=207'b001101000101011011001111001011110010001011010100101010000100101010000001100111110111001100010111001111111000000100101101001101111110111110100010000000000001011111111101100111000001110101001111100101001101010;
#1 $display("%b", po);
# 1  pi=207'b010110111011000100111000110000010000101110101101100010001001101111100111101100111101110100101000101100011101011100101100101001110100111010010110100100010101000000001011101000000001110110111111011000010101011;
#1 $display("%b", po);
# 1  pi=207'b101010000101100001010110110100010100000101001100001111000111010100000111010000011010011011101101101000000011010100100001110101110011100100011110111011111010001100001101000011100011101000011111010101110110011;
#1 $display("%b", po);
# 1  pi=207'b110001111110101101111010011001010111011011111110111010100111010011111001101101000110110100100101111000010110011101001111000011000001011001101011010000011101011001000101001001011011011001011110100100000110110;
#1 $display("%b", po);
# 1  pi=207'b101110110001110011111110111001000100010100010000101110011001110100011110000111101000100011110000100111001010100001000000000101101111110110000101110101111111111111110111110001101000001100011101001101001011011;
#1 $display("%b", po);
# 1  pi=207'b001101110101101111001110111111110110010010001010011011001011110101100111111111100001110001100010011101110110110000100010010111010010000001001111011000011010111010100011010101001001010101100101001011100000110;
#1 $display("%b", po);
# 1  pi=207'b100100111000110101110111111001110100010101000010000001111100111101111111101111111111010110100010110011000011000001100001011010110000011101111100010001011100110010100011011110000100111001110000011010000010110;
#1 $display("%b", po);
# 1  pi=207'b000100100011001000010111101100110011100110011110101110100011001010010000011000111000000000101000111011011110011100110101001111101101011111100001101010101110011001011111111101111100000100110010101101001110110;
#1 $display("%b", po);
# 1  pi=207'b110001000111110011001011010110000001000010100100001010110111100010001001000111010011101111100001111101001011100010000100011100110011001001000001011101100011000010111011111110011101110101100111110011110110011;
#1 $display("%b", po);
# 1  pi=207'b011001101101001110010111001010001011100100000110110001111111111000101111011100010101001010100110010100001000010011000011001101110101110001100011111100000100001011011011001001011101000010011100110101011001101;
#1 $display("%b", po);
# 1  pi=207'b110000101001101010101011110011100001011100010010000000011110111000111100101101110000110111010010100100110011010010011000110110111000000100011101110000000011010100000000101111101111101000111001101010101010010;
#1 $display("%b", po);
# 1  pi=207'b101001001111100000110100000101011111010110011011110011100101000101001111010000100000101110100101100100111001010111011001111000101111101001101000011001010000011011010100001000101101100000011111000010110101111;
#1 $display("%b", po);
# 1  pi=207'b111111011000011101000011100011111111000011010011111000010100100001100111100100001110010110100010100001000111011111111100101101011010010010100101100110011010010111110111011101110111001101111111101010010110000;
#1 $display("%b", po);
# 1  pi=207'b111000100011011001100111001011010011110100000011101010100101001001011111100001000000010101100000000000101110101011101101011101111010111101100100011000101011001101000101110100100010110110001010111101010001110;
#1 $display("%b", po);
# 1  pi=207'b001010110010110001100011001010001100010001101111111101110100001101101101010101001110100101110100001110011001110001100100011010010010010011011000010100100110101100110110111001100001001111111000001111001111001;
#1 $display("%b", po);
# 1  pi=207'b010101000000010101100111011100110110010000101011111101001110100100101000010101001000001110100101101000111100000100111111000000110110010001001101111010011100010000001101000011110100000110111111011110100101010;
#1 $display("%b", po);
# 1  pi=207'b100101010001011110100011001000001110011010111110010000011110100011001101111011001111100101100000101001001100101100011111011110101100110100100001100101100010100010000100111010100000110111001001010111000101100;
#1 $display("%b", po);
# 1  pi=207'b110010001000010011110111011001010111100111100001011010001001100010010100100101110111101111100010111111011110011110000100110110101011010011110100010110110101111000111110001000101010100111111100110100110111100;
#1 $display("%b", po);
# 1  pi=207'b110111111110001011100001010001010111101110010011001110010001101010111001101001011001000010100100101111010000011101000000011100100111101110000001101100111010001011001100100100111101100111011100000010001101010;
#1 $display("%b", po);
# 1  pi=207'b010101101011101011101000010110011001001001001010001010100010110100110100100000001110111001111111110001111001110100111000000101010011010101001000000100110101011000010110100111110010111010101101111000011011100;
#1 $display("%b", po);
# 1  pi=207'b100101101001111111000010100001011101101111111000010111010000101000101110111101001101001101111010001001100100010111111111011001110110010011111010010111011110001001110110110001010101001011100111101000110111110;
#1 $display("%b", po);
# 1  pi=207'b111010110111011000111111000000001100011101000000001100101110111110101101100010011100001110001110100010001001101010000011100111000111101011000111101011010000100101001000101111010010100101000000010111001011100;
#1 $display("%b", po);
# 1  pi=207'b111000110110100100110011110000110001101110011111111011011001111001101011101100110000111110001010001000011001000001110011101011011111001101110100000101110011110110011101001011100101010000100011000100111110001;
#1 $display("%b", po);
# 1  pi=207'b001011100110010001011100001010000101101100100010010111100101011101011111001100101101100000000000111001111010000011001110101111111000010111011000001001101010110011001011101110001010100100000110001101010011010;
#1 $display("%b", po);
# 1  pi=207'b110010100001000011101100110111001100100110101101011111010001100001110000111111001001010010011111111001000101100110111000010000111111000011101110010111101010011000100011001011010000001110101000110000100110001;
#1 $display("%b", po);
# 1  pi=207'b110111000110001100101110110111100000010011111100001000010001011010011100110011010011011101110000010011110110010100101001110011000100110101110000011100111101100111011011111010111110000100110011010000100111001;
#1 $display("%b", po);
# 1  pi=207'b111100110000010010101110111111110010000011001101011010101110000010100111100111011010101111100000101001000111010010011001011001001101001101001100111110011011011110110111110000011011010011001011101110000111101;
#1 $display("%b", po);
# 1  pi=207'b100010010110001100110001010001001100011010110011110110000011110111100100101101111011101011100100100001000001010010001001100111010010010011001010101001011001111000011100101000010101011110000101000000001111110;
#1 $display("%b", po);
# 1  pi=207'b000111011111010111000010011000001111001010101001000110011001010001101000101101010101011010011111000011101011000000100000001011110101100011000100110100010001110111101100101000101010011100001011011101101011110;
#1 $display("%b", po);
# 1  pi=207'b011010110111110101101011010111011001110101000000111011001011000110011000111111001011010001000001011110010111010000010010100101101011110010001011101011110110000001000000011000001100011000011011101000101011110;
#1 $display("%b", po);
# 1  pi=207'b101011101101000011110111110101111010000100001111011011110100000110011100011101011011011111011110110110000011010011110110111110011101011001001010111100100010011110111101011010100010111111111110001111011111001;
#1 $display("%b", po);
# 1  pi=207'b100010101011000100010111111111110010010000110101110011101000101011001011100111010001010111011111100110001110100111000101101011111101110111000010100000101011110100001100101011001101010100000011111111001000101;
#1 $display("%b", po);
# 1  pi=207'b101000110111000001100101110101100000110011101010001011110101010110011110101010101100111111001001111001011100110011110100011101011001001111111111010100110101100100110100100001000110100100100101110010011001111;
#1 $display("%b", po);
# 1  pi=207'b100001001000111000110100001100010001101100000101110100000000001100001010010110001100100011010010110100001100001101011001001001001001101011010000110100111110011101001110111011101101110011001100100000111111101;
#1 $display("%b", po);
# 1  pi=207'b110010111110100011011000111100100100000001111011101101100101101001101101010000011110010011001111101101111110001110011111010100011001110000000101110010010011110010011110101110011110111010110111010111011001000;
#1 $display("%b", po);
# 1  pi=207'b111000010001110011011001111101000110111101111001011000010101101000100111001001110101000000100111010011110011101100110100000000000100111110010100001100010111010010101100001000010011001000111001010111011111101;
#1 $display("%b", po);
# 1  pi=207'b010000110011110011000101011001010010100100110110110000111010101111000110000101000011101111111110100101000101001011100001101010010101010000100111001111111101001001111010111110011101101100100100011001010011010;
#1 $display("%b", po);
# 1  pi=207'b100111101100011011001111011001011101000101111101011100000101100011010110001101110111100111010000011101100011001011110011010010100001100111010111011010100100000110111011001111000101010100111100000100011010010;
#1 $display("%b", po);
# 1  pi=207'b000100010011101101000000000100001000100111010110001001011110101010110101001001110001001000000101000001011100001110100011111110001100110001101100100110101110011000111110101000011001100010001000011101111111001;
#1 $display("%b", po);
# 1  pi=207'b101101001111011111000001110000010010010001011101101110101110001100100010110110001010000001011000110111010111101100101111000000100010101011111001110000011011111100111011011111101000001000011010001011001010011;
#1 $display("%b", po);
# 1  pi=207'b011011101011111001000111001000111100011001111100110110001101110100010010111011111100111110000010011011010001010100110011010011101101110011110101001101001001110001111100011011000100101100101011001100111100101;
#1 $display("%b", po);
# 1  pi=207'b010101001010011000001010100100001100110010100000110101001111000010110011000100001100111100101101000110111000110100011010011010100000010010011111001110000001110110000000000111100100011111110010011011110000101;
#1 $display("%b", po);
# 1  pi=207'b001010011110101110101110100001000011100001101101100111011110110111010011011000010001100000010000001101110100111001010110101001111100100110100000011010111010100101111101010111101000000101110010111011000000000;
#1 $display("%b", po);
# 1  pi=207'b100101100001000100001000100010001010111111001111001010101000100101000001010101001110110110111111010011111111101000111111001010001100000000111010000101110100011011111101001100010011011111100000010000100110101;
#1 $display("%b", po);
# 1  pi=207'b011101011101001011100100110110000010101000110000101100001001001010101110110100110000010100111011101010100101101011100110100111101100101100010011101111001110011101110110011100111001000101010000110010111111001;
#1 $display("%b", po);
# 1  pi=207'b111101001111101010010101000001000110010011011100010010111010111111000101001101101000110101001100001010011101111000110111011011000101110001111100000100110101101111001110011011001010000001011000011100101011010;
#1 $display("%b", po);
# 1  pi=207'b110110001001010011001100111110011010101011011011010101100000001111001000000000011000011100000001101001010101010111000001001110111000010000000101000101101111001010010101111111101110111110000100010101001100011;
#1 $display("%b", po);
# 1  pi=207'b101010010101010001111111101011101001011111100000010111110100001111110001011100000001100000110000000011011100000001100001000011011110111100001110101001000111110011110101111110100101110110011000010010011111100;
#1 $display("%b", po);
# 1  pi=207'b011110011011100001111101100111110010101000010011110111110011010101000100110001000001101101111111101011011011010001000011001111110011100101110011111000001011100101100101011010010111101000011011100001011001101;
#1 $display("%b", po);
# 1  pi=207'b001001111001111000101101110000111001001111101100000000011110101011100101110110010001101010000111101110100100001001000100000010110110001011001011010100110111101111100100110011011110000110000011000010011000100;
#1 $display("%b", po);
# 1  pi=207'b111010000110010110101001001111001100010100011000110000100010100000111000011010101010011110111010100010101110000110000000010101011011001000100011111010010010100110001011110010110000110010101110101001011010010;
#1 $display("%b", po);
# 1  pi=207'b000101101100110111111111101010000111110011011011001110100110101110100000010011011100110110111010001000001101001101001101000101101111001101011111100111101111111111010001111000100000001001001100100011110110001;
#1 $display("%b", po);
# 1  pi=207'b001011111010111010011110111000110011000001001111000100111110010000110011101000011110110010110011110101010111110111010001111100011110101100111101011101010111111011101000100101001100100001111100111101100100101;
#1 $display("%b", po);
# 1  pi=207'b100111000010100001011010011010001000110010110100000010011101110010000101110000101011000111010011011111010110110100101101010000100110110011110011001101011110111110011100110101010011011000100000010001111110100;
#1 $display("%b", po);
# 1  pi=207'b010110101011110101100110000110111011100110001111110101011101000101001110111110000011110000100101001011110110001000100011101110011100101111001101111110000000001011101110100110010110101001000011000010111011111;
#1 $display("%b", po);
# 1  pi=207'b110010111010000010011100010110111001101101001110101011110101101001001000011100110010001001101001110000111000110101111111010001011110100001010100110111111000111000100000011111011111111101111000100111110001000;
#1 $display("%b", po);
# 1  pi=207'b001011110000110111100000101010010111001000001001101010110111101111010101101101000010010001100111011101011110000100001100110010110000110101010011101101110011010001010000111000101011111010000101111000101111000;
#1 $display("%b", po);
# 1  pi=207'b101000100100110000000100101101010101111000101010110100111010110010101000010111000111111011010110101010000100111000100000011011011111011110101011110011010111011100011010001010000000001001011010101010001011100;
#1 $display("%b", po);
# 1  pi=207'b101110010110111110111000001111010110111110111101111011001111010100000100111000011111011101000000111000101011011010100101111000001000110010010000101100110101111000001000101111100100111000101011010001110000101;
#1 $display("%b", po);
# 1  pi=207'b010011001000111000000001100111111110111010000001011011011101101101101111110100111011000101010101010010011011111111010001011010111100010111011000000110111111111101111001011100100010110001001111011111110110010;
#1 $display("%b", po);
# 1  pi=207'b001100000001100011001111100111011000100101111010000011101011011000111100001101000011110000101010000101100010111010011101011110101101111000010110001111011000000000010101010101100101001001011111001011000111101;
#1 $display("%b", po);
# 1  pi=207'b011011001011101001110001011100011100101011110101010111001111001101011001101010111010111001001000100100001011000001010100011000000001100111011111011101011010010101011011011111001001111111000100100011110111111;
#1 $display("%b", po);
# 1  pi=207'b010000110101100010100111011101100010011000100010110010111011100101100111111000000110101111100010001100101101100111000011111110000000010011011010001111010010010011101101111011010010001000000001001010010111100;
#1 $display("%b", po);
# 1  pi=207'b111110111110100101011100011011011110001000010011011011100001110011101110110100011101101011101110010111101001000111011001001000001101010000001101011000011110110110100011011110010100010100100111010000111011110;
#1 $display("%b", po);
# 1  pi=207'b011101100000110110101110011010101010100001010001000001001100000101000000111101011100011101100010001000100001110011101100110101010001001011010001000110100100011111011011100000110100001011110001000111000110010;
#1 $display("%b", po);
# 1  pi=207'b011100001001011000010010001000000011000110101101111010001110011001000010001010100101100111100011001101110110011111011101110110001011011000100001001011011011000101000101000111001010110011001100100110101111110;
#1 $display("%b", po);
# 1  pi=207'b100011011101010011011010100111011100110110011001101011101011001001001000000001000011100101110010111000001000111111111001010111011101100100011011000000101111001110100111101011111000110011101011111000000011010;
#1 $display("%b", po);
# 1  pi=207'b011110000001101010111001111100000100001000011011011001111111100000101111110101011111111000111000101010001100101101011000001101110111000011111110010011100111100011000010011110100001110101000010110110101001001;
#1 $display("%b", po);
# 1  pi=207'b101110101000000110000110001001110001010101101100000000111101010010101101100100010010000101111010110100101000110001100101001101000001000011000101110101001011010000000101001100000010100100110001001111000100000;
#1 $display("%b", po);
# 1  pi=207'b110100101011001000110110001110001010000100100100001110010100001011100000000011101000101100010000001000111011000100101100011100010001011000101000110001101101111111010101100110101001110010011110110010001110010;
#1 $display("%b", po);
# 1  pi=207'b101101001011010010011100101100010101010100001011000111000101111101000100101010011010001101111000100010101111001011011101101001111100111110001010010110011111001001101001000100000010010010010101011111010101010;
#1 $display("%b", po);
# 1  pi=207'b010010110001000111001111000110001110011001111010000010000111100111100110100010000111101011101100011100110001110000001100100111011110100100011000111001100001010111101011011010101110111011010000100000010101101;
#1 $display("%b", po);
# 1  pi=207'b001011011100001010101010110010110001011111011001111111011010010111011101110111011001000011011101101110100010010111011110101001011001101110100000011011101110100011110111111101101101111011110010001000000010110;
#1 $display("%b", po);
# 1  pi=207'b001101101010011000010100101100011000000100110010010011010110011010011001101110111011001011100001011110011100000011101001101011010010000101100011000000010011011100101000110111001111011010000110000000001111001;
#1 $display("%b", po);
# 1  pi=207'b110111101010100111100110111000111000101100101000010000001100000011000110101111010100100110111000011011000100110100110011011101110100111011000011111101010111101000111001111011011100111001001011111101001100010;
#1 $display("%b", po);
# 1  pi=207'b111000011001010111100011011000000101101101000111100011000000000001000000011001101110010100010001011010110001011011001111101010010010100100100011111101000111010111101000000000010101010011011011101110111100111;
#1 $display("%b", po);
# 1  pi=207'b010110100110101111110011101010101001010111000101011001001011110100000000000011011111001001111001100100111000110100000000110011001110000101011100101000100101111001010101110110011010100001010011010110110000011;
#1 $display("%b", po);
# 1  pi=207'b001110011010000011000101010010010110001011011000001100111110100011100101101100011010111010100111001001111110001001011100110110111010001101001110010100100111010001111101100011000001110101011111010011100000010;
#1 $display("%b", po);
# 1  pi=207'b001110100001110010011100010110000101011001001001010100100100000100000011000111110100001001110011001111111001101111000011110001000110101111100010100010100110011100010000110010010001010010001010100100111000101;
#1 $display("%b", po);
# 1  pi=207'b000111100001011000001100001110000001001110000101010101110001001010110010101110010011111011101110011001000001001111101011011010001001001001110011000001001101111110000000010011000100100111101100010011011001011;
#1 $display("%b", po);
# 1  pi=207'b111111011011010100110000010100010001110011100000110111000011101001010000111010000010110110010101011001100110100011011000010011110100001101011101101111100000000010101100011001111010100110110110110101011100110;
#1 $display("%b", po);
# 1  pi=207'b100011001111100111000110100001010010110100110001010111011011000110100001101110011001001000011001010011111100010010001010011111101100010011111101000000100001111010110001001000010110101111010111011101001101010;
#1 $display("%b", po);
# 1  pi=207'b000000100110110101011100010010100100101000110001000000110001001010100110101101111110010101000101001101000000011000001010011000100011111010011100111101111100010010110001101000001011000000110011111001100010000;
#1 $display("%b", po);
# 1  pi=207'b010110000011000011110101101101110111111011010001010000001010000110011000110010110000001001010110011011101110110110100010010001110010110011110001111101110100000000001111101101100001001001011100011010111101110;
#1 $display("%b", po);
# 1  pi=207'b011111101101111000100111111101100110001010101011000001111011110110000111001011000010001101001101101001100001010001101100110010001010011011001110010010100000101100111001101001001111001000000011100110111111111;
#1 $display("%b", po);
# 1  pi=207'b001010011110101000110101110000101011101101100100000110011001000100100010000011110010011000110110000110100110001001011010111011001110100101000001000100100101010111001101001110001110110110011100101000111110111;
#1 $display("%b", po);
# 1  pi=207'b100011010100000010000100100110111011001010010100010100100111000110100111011101010010110100011100110100111001111000111111100011110101000010101101000011011000111111010111011100110101011001110100110110110101000;
#1 $display("%b", po);
# 1  pi=207'b110101111001100011000111011000110000000100100010001011101111100101001111100001011011100001000101011110111101001100011110011100001100110101010110011001111010100010111010110100100111111010100001010001101001111;
#1 $display("%b", po);
# 1  pi=207'b000000101010010110100101110101001100111011000101101101100111001101110011101110000101111111001110000101010100110101110000010100001101100100010111100100000111101011101110001101111101010010000111010011100101100;
#1 $display("%b", po);
# 1  pi=207'b010101111110001010100010101010010001001101101010011000010001011011110011111010101010111101110001001011001100001001000001011001000100101100111010111100111110111011011001111101011000000110000101010111111010000;
#1 $display("%b", po);
# 1  pi=207'b010100111000001000001011111101001001011001000001101001011101101110000001010100100010010011010011001001011010000001100111011110001011001011000011001110000001001001100110010111101110010101010110011101101101001;
#1 $display("%b", po);
# 1  pi=207'b111111100110011100101001100110111101111101010101111100000011110000001111001010011011011001010010111010000100101011101011100011000100100100110111100100011011111110011110001100001100100110001110010100010011111;
#1 $display("%b", po);
# 1  pi=207'b010100000010001110110011101000110111111011011100100011111101101100110000000100111111110111100101010100111000000111110000110011001101000101111100101110001111010001000110110011100100010100101010101101011011100;
#1 $display("%b", po);
# 1  pi=207'b001011000011001101110001101111100010110110100000010011011010011000100111000001100001101000000010111011110100000101000011010101000101110011111000000010101101011111011111010001011011100101100101110011000000010;
#1 $display("%b", po);
# 1  pi=207'b101100011101011010101000000111100000010010000000101111000100111000100011100000110100111011010001000011010000010000101010011001001100010111001010110110001100111101011101101110101111011101110110001001110111010;
#1 $display("%b", po);
# 1  pi=207'b010011100111010110101011010001111000110101011110100101010001010111101010000101110010111101110101000110111011000010000010010110010011110111010111011000000001100100111111011111100101010011000000011110101001011;
#1 $display("%b", po);
# 1  pi=207'b110101110011001010100111111010101101011100100110110111110011101101110111001101000110001011011111111000010010111110010101100111010000011101011100100000100100111010000010110010111001100101111001010000010101110;
#1 $display("%b", po);
# 1  pi=207'b111011011000010110011110000000101111110101000000111001000000110011001111100011101010101001010101111100010101011111110101011011000010111101111110010100010010111101110100100011101100111110111101101110011110101;
#1 $display("%b", po);
# 1  pi=207'b010110100111010100111111110010000100101011101101101100100001101101111111011110100111101101001111001101101010011100010011111010100101100011011010111101100110011011110011011111001001101101000001001100010001111;
#1 $display("%b", po);
# 1  pi=207'b001010011010010011110101100111001011101010010001010111100111011100001111111001000101110100110110101011100110100000000011011010100011101101011110111001000000000011010101111001000001100000110001000111001001111;
#1 $display("%b", po);
# 1  pi=207'b100001000110100110011011011000010101011100101101001000100001010111010101001111010110011011000000000100100100000111010110110000001011100000010011011011110101110111001001101101111111100001110111101001000011011;
#1 $display("%b", po);
# 1  pi=207'b001011100010010010110010000110111001011111100010101111101000001110111010110010101100000111001011111011001111111011110010111100011100001010111110101011111011111100100000010111100111000111001011100001100111101;
#1 $display("%b", po);
# 1  pi=207'b001001001000101111100001101010110111100110111110010000111101110000111010010111111000011010110111001010101001001011010111001110101101001110001000010010000100100001101100001100001010101000000011101010110100111;
#1 $display("%b", po);
# 1  pi=207'b100100100101100001100011011000110100011101001110111010000011011111110011001001101111111110011111000110101100100010000010010111101011110010101101011101110100010100000100100110010011001011000101111101010101101;
#1 $display("%b", po);
# 1  pi=207'b010101101110111100110001111001010000011110010010111110010011000001010010011011000010000010100001110101100101000111101000111000101001000010011100011111100100000010001000100011111111000111001111000011010101111;
#1 $display("%b", po);
# 1  pi=207'b011011001000010101111100000000001100000010100111011001100100101101010101011111101000101100000001010001001100111100001101000110010100011111101001011011001111101111001110001101100110111000001110101100001111100;
#1 $display("%b", po);
# 1  pi=207'b100100111000001101100011110101111010100101101000001000110111011101111111111001101000000111001111110100001010111000001001000100000010001001110001111000011101011000111111000011101010100011101011110000101000101;
#1 $display("%b", po);
# 1  pi=207'b101110111101110101001110111011110111010010001001110010110100000010011000011001000110100000110011011111011111111110011000001000000101010110001000000111100011000000011010101000010011010001001111110111110000000;
#1 $display("%b", po);
# 1  pi=207'b100001001110010110101001111010100100101010011100100011000010110001100001001111100010111010001110010010100111000000011100111110101010110110010100000100010100100100101010110110001101111100100000010000101101000;
#1 $display("%b", po);
# 1  pi=207'b011000011010010111101110000110101001010110011010011111000001111000111101101111001000000010010000000011011010001101010010011110010101101110010001101100001100111001111111111000010101000111010000000101101111011;
#1 $display("%b", po);
# 1  pi=207'b001000101101000111101110111001111100100010101101101101010011100101101110001001110100110111000101010111001110100110100101001000110111100111001100010101011000001100011000110111011000101011111111010011000011111;
#1 $display("%b", po);
# 1  pi=207'b011100011001011010010111010100110100110000101000010000100000010110100111111100101110011101011110101100100010001110000010110000101001010000100001100110101101000110010010011100100000111000110100101101000100101;
#1 $display("%b", po);
# 1  pi=207'b000110001010000011001010101010100111010010110010101100010110011000111001001001011111000001100010001100010000001111010001101110111010111100010110010011010111000011010010000110001011010001000111000000100001101;
#1 $display("%b", po);
# 1  pi=207'b101101011000010111101001111111000100111111000110101101110011000010100110111010011010110000100101101111100100000101101111000001110111100000100101100001011010000011011010100011010000100111111001111001111000011;
#1 $display("%b", po);
# 1  pi=207'b101001111011111111010000111011010010001101011011000100010010111001011111011001001110111100001010001100110100000010101000010101011111011011011101011110011101000001100010011101100000000000000101100000100011010;
#1 $display("%b", po);
# 1  pi=207'b100111111101011000100000111000101011011111010101001101001101001011100100110000111000000111101111010010110111011100100100110000001001100110110110101111101111010011011011011001011000110110111011010011100000011;
#1 $display("%b", po);
# 1  pi=207'b011101000011011010111111111010111000001010001110010111101010010110101010110011000101000001010010011110011010100100110100010100010011011101010111001011111110000001000011101111001111010011011100011101110011111;
#1 $display("%b", po);
# 1  pi=207'b111101010110111011011011110011010011100001100100000101000101110010101110011010110001011110011001010010100110101010000010000000011111100111100010010101010001101000011110001100010111111011010000001001101010101;
#1 $display("%b", po);
# 1  pi=207'b001110111010110011111000110110000100111011000101100101010101111000100001000010110010111100000111001100011110111010001010010110100100011010101100100011001010001110111010100101000111100011000111010011110111010;
#1 $display("%b", po);
# 1  pi=207'b110001101001001110110011101110110011110010101100100100010111011111011010101110111110110011010010100010000011100010110111010110001101101011100010010101001101100001100110111110011101110110111000110101000011000;
#1 $display("%b", po);
# 1  pi=207'b000001000001111111010011100101100001001100111111011010100100000011010001000011110000100101100010010101001001110111011011111110000110001100011111100110111111110100000000110000100100100011011011000001111000000;
#1 $display("%b", po);
# 1  pi=207'b101110100011111110001010101011101110111001111001001110110111100110101001110110001011110100000100011000001000101010110000100101001000110110010011111100110001000100100000011101111001111000100000101000111111100;
#1 $display("%b", po);
# 1  pi=207'b101001111110110011001111100011011000101101110100011101000000111111100001101100010000101100000101000111110111011111010000011011111111010110010111000000101101101000111011000010000101110001010001101010111000101;
#1 $display("%b", po);
# 1  pi=207'b011111101010111010000110100011101000101011001010101011011101110010011000010111110111111100001011100001000110110101111001101101101010100100011010100110011100010011010100101000101100000111001011100000010011101;
#1 $display("%b", po);
# 1  pi=207'b100000110111101111100111011101101111100110111010100101101011110010111010010010111011000111101110111000000111101010000110111100011111100011010100000111110110101000101100100010111010010001000010010011001011111;
#1 $display("%b", po);
# 1  pi=207'b101000000001010001100001110101100010000011011110001000000111000010010100101111010101011101011011010100011100010011110010101100111110011001101010011001100001101010000110001010001001111111011011111110111101010;
#1 $display("%b", po);
# 1  pi=207'b110001011010100001111000010111101111101000100110001111011001100101010110000100000010001100111010010100011100111011000001001100110100001100001000111110001111100010100111010000111001111000001001000100101000101;
#1 $display("%b", po);
# 1  pi=207'b010111000001011110010000101110100001000001111110000100111111101001111111000101011011110010011011010100000001111000100010100000110111110111100110000100010000000100101111011111011010001101010011100111011100100;
#1 $display("%b", po);
# 1  pi=207'b111111111101000101111001001011101000011111110001011100101101011111110100010001100101010001100000000000010101001111000001100011011101001101101001011000101010110000100010011001000011100100001001111010111111001;
#1 $display("%b", po);
# 1  pi=207'b101111100000111101101101001100111000101100001000001101101011111110011101001111111100111101001001101100000010001101101101110000000100001110101110010011011111011101111101100010000100100110000011100100001110001;
#1 $display("%b", po);
# 1  pi=207'b100110110010110110110010110100101101000000001001110011100111101110111011111101101111000100111010010110000001010100010110100000000000000000000011000010111101101010001000010110110010000011110001001111110001101;
#1 $display("%b", po);
# 1  pi=207'b001100011001010101011111100111101011110010000110001111101011101001001111100000111000101000000110111001001100011110100111010000010100000110110100001010011100111001011110111010001111101001001100001101111000011;
#1 $display("%b", po);
# 1  pi=207'b100000100101010100000101110001011011110010110001110000101011001011000010110010000100010100010011011000010011000100110111100001101000111100001001100111111011001001011011000011000001000011000001010100011100010;
#1 $display("%b", po);
# 1  pi=207'b010110111100011111010111111110000000010100001111111010111001010100111001110001101100011010100111111010100101100110011001100110110001100110000101011110000010101011010011100001101000010100010101000111100001111;
#1 $display("%b", po);
# 1  pi=207'b100001100110010100100110100000111001110010011010000110010110110010101111011010110010101000110110100111100100100010100101101101000101000001100111111100111100100011000111110001111100100011010011100100100001000;
#1 $display("%b", po);
# 1  pi=207'b110111011000011101001011101101011011010110011001110000001101011101000101011111001011011000011001110101000101101001100110011111101111110101101111010010001101111000100110100011111111011001101011000101111100111;
#1 $display("%b", po);
# 1  pi=207'b010010001000001001110110101110001100010100001111010110000100000110000011000000100101100101001101111110011111101100110000110000101000000011001101010101100011100100111111101011111100000011101011111001011010010;
#1 $display("%b", po);
# 1  pi=207'b010000011001101111101111100111110010011100011100000101101111010101110001100001111110101001000101111110011100101000101001110110110101011010011110001010100010110100010110000001000110011100110001100101100001000;
#1 $display("%b", po);
# 1  pi=207'b000010001101000000010000111100000100100111001011001110011111001101100010010111101101100111101001000001110100000001111110111100110011110010100110110000010101011010011001011001001101110000111011000110010100111;
#1 $display("%b", po);
# 1  pi=207'b111011011100011101010001100100111001100001100101101001000010100010100101110000011111000000010010101000001010100010101100010011011101011011000010000101000110110100000011100000011110100110010011010010101001111;
#1 $display("%b", po);
# 1  pi=207'b010110110010011000000111101001111111110011000001001000101001000000011000100001100000101010010110000010000011010001110100110101010011100001111110111001101011001011001011101111011010001100011111101001000100100;
#1 $display("%b", po);
# 1  pi=207'b010100010000000011001010101011101000111001001010000000110100000000000000110101110010000010111010010010000100010010100100000010001001001100101100110011000010011001101100100111110001011111001101011000111010010;
#1 $display("%b", po);
# 1  pi=207'b111001010100100111010110110100011011001111111001100011111101011100010000101100000111001100110000000111000111011011001110111111011100010101101011101110001111110111001110110101000010000001000001110010011101001;
#1 $display("%b", po);
# 1  pi=207'b010110011100000000101000111111011101111101101111011001011110101100111000100110111111101111010001000100110110011010010100111000001100100111100001101110111000111001010000110011001010000111000001001101101111110;
#1 $display("%b", po);
# 1  pi=207'b111101011000010101110010101001101111100110100010001100100000011110111110100000111110111001111011010001010111001100011111100100011111000101000011011101110000100011111101100001010111101111100001100011100001101;
#1 $display("%b", po);
# 1  pi=207'b010111010001010100001101011011001110010000010010000010111100011111001001011011000100010011111001101001000111110001100101101000010101110000000010100000100011000100100001101010011011000110000000010100011001110;
#1 $display("%b", po);
# 1  pi=207'b011111000100000101001110000010001000010001110110111011010001000111110011100011000010110000010101010100001010110001110001010111100010111111001001010100100010001011100011100010000111111101001011011100001100101;
#1 $display("%b", po);
# 1  pi=207'b011100000010100001001011000101000010001111110011000110101000101001111111010010110101100101111010110100110100100010010001101011110101110110000011010010001110010010110010111010011011110010000000101111011100010;
#1 $display("%b", po);
# 1  pi=207'b111101111011100101011110111010011010110010101110001010001101011001110101001101000011110111001110110111000100111101111011011011011101000000110110111010000111000110011001000011001011011010001001000110011100000;
#1 $display("%b", po);
# 1  pi=207'b001011000100100011110101010000101000111000110011111100000000101010000110111100000111001100111000000010100000001011010001111011101100101011101101110110111011111110110100111010110111100101101101100011111000110;
#1 $display("%b", po);
# 1  pi=207'b010111111000000110101000001101010110000001001011011110010100000110011010101111111001010101000111001000100110111010000001000111111010100010101110010001000110111110100011110101010110011001001010001111111101111;
#1 $display("%b", po);
# 1  pi=207'b001001011101100000000100100000110111100101101011100110101100000011101000010101011101110011011000011011011111001111000110011110100111000001110111111011101010001100101011101110110101110000100000001111000100011;
#1 $display("%b", po);
# 1  pi=207'b110111011001000011100001000001010000101010110000111101000100101100000001101011010000010100011001000000010011110110010000011110010010010010010010100000001101101001011000101001100101110101110001101110110100101;
#1 $display("%b", po);
# 1  pi=207'b000011001011000000001001110110110001000011001000110000001000001100001011000101011011101101101110110111000111000000010010001010010110001100101100011111111101010001101111000101001111101110110000111101100011010;
#1 $display("%b", po);
# 1  pi=207'b001011010000110000110001000011101110110101100010000011111010000101000110111011010101101011010011101100100010010111101110111111101100110100111101101100100100101111010001101000100100011011101000111010010110011;
#1 $display("%b", po);
# 1  pi=207'b111010011011010110011001101000011000111001110011100111001111101110111110010011101000000101010101000111101111100100111100101100010111111110001110000000111101011000001111101001111110000010001000000010001000100;
#1 $display("%b", po);
# 1  pi=207'b110100011011010011010100011111011110001001010101001100000001110011001111011011011100100100000100101111100101011000100000100010100000110001011010000000101001101111100100011110110110100011100000010110010000101;
#1 $display("%b", po);
# 1  pi=207'b010000011010101000101010011011110111001010011111101000101010101011011110011001100010010011100100111011101101010000000110100001000100101010001101010011010010010111000101000100000000100011100010100010101011000;
#1 $display("%b", po);
# 1  pi=207'b010011101011001000101110010001111001000010011001001100001011010001011010001111000100101010001110110001011010011110111110011110010000100101011101101111000111111111011001101101111001111100101001100100101100011;
#1 $display("%b", po);
# 1  pi=207'b100100010111111101111001110111011001110010111001111100001110000011001001110111111000100111000011111111000110111110001101110110110111110100010101011100101101011100011101101111110111011101110100101101110111101;
#1 $display("%b", po);
# 1  pi=207'b001111000100100100011010101010000101010101011010000110101000011110101111010000001100001001100110001011010111101001000101000010100110111100000010101001101010101010010111100011001010111000110011100100101010000;
#1 $display("%b", po);
# 1  pi=207'b010000011110111001000011111000100011011001100100110110111101101111011010110111101011101100110001110001010101011111001001001010010110000011001100001111000000100100000111111001010010001000001111111000010101101;
#1 $display("%b", po);
# 1  pi=207'b010110011110011101101100101110000001110010000111010001001110001010110011010101011101100011011011100110111110101000010111011110111010011000001111001101011110101011110011000100001000101000000111011111011011110;
#1 $display("%b", po);
# 1  pi=207'b101101101111111001110010000100001100011111011111000001100110011011111101101000000100010001111100001001011110010010010101110101110101111000011000111010011111101101110001010110101110110111100110000001100111110;
#1 $display("%b", po);
# 1  pi=207'b011010011011100010010011001100000100011111011011101101000010001101111011100001101010100110001100000011000101101000101010011001101110010111011100001000111001100001000000110111100001011110111111110010000101101;
#1 $display("%b", po);
# 1  pi=207'b010011101110101101111110010100001100011110111011100101001010010011110100100000101101000011000011010011110001000001111100010001100001111000011100100100001001011000000111111010111101111001001110100001001010100;
#1 $display("%b", po);
# 1  pi=207'b100111011100011001011001110101100100100001110111101110010111011010010110101101000110100001101111101010010000101000111001100111011000001101011110011100111110010000101011101111001000000101100010000111001111110;
#1 $display("%b", po);
# 1  pi=207'b110000000111000001100111010111111101000110101111010111010110000011101101111100000011110101101010110111111000100110010000000110000010110110000101000001000000001110100111100000010110110010110010110100101001000;
#1 $display("%b", po);
# 1  pi=207'b000000111000100110001100010100001100110100010010111010011111101001101101001001000100001110101010001010100101111110011011110000001011000111100101000001111100010011010001010000000011001100001010010010011101010;
#1 $display("%b", po);
# 1  pi=207'b011101000000001000000011101001001100001101011010010000110001110101100100000101011110000000010011011001011010010001100101011010110111110111110001001000110011111000010100011110111000110111100101110100110110000;
#1 $display("%b", po);
# 1  pi=207'b111001111111111000101111110110010100010000001011100011110101101101010111110000010011011001000111111100001001110110110100010111100111011110010000011000010000101001100001000011010001100010110000010110100010000;
#1 $display("%b", po);
# 1  pi=207'b000110100101110010111111110001011001010111000101001110100010010001010111110011001101000010000111100001111000111110011011011010100001110100001111001001001001111100011011101100001101110011111010000010111011110;
#1 $display("%b", po);
# 1  pi=207'b010001001101001100010001000000101011111100101111101010010100111000110101010010001111001011100001111000110100000010000100111111001111001010001010101100110010111000100000101010100011000101111100010001000101110;
#1 $display("%b", po);
# 1  pi=207'b010010101110101100000110000011111100111011111101010111100001111111001110101000010011110001100011101001000000100001111011000100101000011110111000110101011100001011000000010000111001110010100011011001101110001;
#1 $display("%b", po);
# 1  pi=207'b011101000101001011010001111010110101011001100100000101111110001011111110011010110110110000110001101000011010100101000100101001110101011011101011110110110000010101111110000100111011000010001111111011000100111;
#1 $display("%b", po);
# 1  pi=207'b101111010110010100011001001000010111110011101010100011010001110010000010101101111101010110000001101101011010111001011111011001000110011100001000010011011111000110010110011100101001110111101000001101111110000;
#1 $display("%b", po);
# 1  pi=207'b010000111111111010010000000110000100000000111001001011011100111000000110010100000001011100101110100111010011101100010101001000110100000111110000011000101110001101100010011011000000001010010011010001100011101;
#1 $display("%b", po);
# 1  pi=207'b000000101101001010001101011000101101101110000111010011000100111101100001100001110111000101010111001110001001000101011011100101000011000011111100000011011011001011110110100000110111101000000111010101100101000;
#1 $display("%b", po);
# 1  pi=207'b100111000010110011101111110011110110010001001000110010000001001000011010011011011011101100100010011010110010010001011011010100100000011101000000001011011010001100001110011111011001110101100101000001111101101;
#1 $display("%b", po);
# 1  pi=207'b101010110000100110101111101000000000000101100000111100001101110111000010000101011011010101111100111101101000001010111010100001111010111011010011001110101001001011111101111100011110010110011000110101100001000;
#1 $display("%b", po);
# 1  pi=207'b100111100010101101110010110010101000000100100001110011000111000001111011100110100100011101001100001111011100100100111100101111101000000001010111010100110111011011010111000111010011110011101110011010110110010;
#1 $display("%b", po);
# 1  pi=207'b010010010101000010010111111111110100110111010101000010110111000000110101011011010010100110111111000101011110011010000000110101011001111010000010010111110111011001111001111111001100001011110111100101000111000;
#1 $display("%b", po);
# 1  pi=207'b101001110000010000110000011111111001101111100110111110111001101111001110010100000011110001111010001010000111101000011000010101100011001001000110010100100101100111110011110101001001000110000011010010100010011;
#1 $display("%b", po);
# 1  pi=207'b011110101111110010100000010101110111100100011100001000001000010001001011100100000111000000111000101000111111110111110010101001011100110111011010110101000000010001000001001011101001110100010010110001010010101;
#1 $display("%b", po);
# 1  pi=207'b101110010010111010110100101100100010010100111101101101100111010001000110000001000010001001111111111101001110011101011010000111110011010010111110010000011111111001110010000010000001100011011111110011011111011;
#1 $display("%b", po);
# 1  pi=207'b010011111000101111110010010011011101001111010000010010111010010110000001110111110010011011101100110101100110100101111010000100010100100111001010000000010111000110000001101100000101110110100110100000101011100;
#1 $display("%b", po);
# 1  pi=207'b011110100011000111000001010000100011100110011011010000010010111010010100000100011001101010001110101111011000100100110010010010000011011000010011100011101001001001100011010011110010001100101111001011111010000;
#1 $display("%b", po);
# 1  pi=207'b101110010110001010011010010011111001001001011000101011000011100000111100001010000101111101011011001000110100100010100111011100111010011101001001100011101011001000010111001101001100110010101010010110100010101;
#1 $display("%b", po);
# 1  pi=207'b111000100101101101010011100000010110010011010100001111000011100000010100011000000100101011111101000100101101011100001010111100011001111001001101111100100000010111011011101100100110110111001010111001111001000;
#1 $display("%b", po);
# 1  pi=207'b010100011111001000000001000001001101110110101110011001001000000111011101011001011101011011101110010101001011101111101000111010001101001000000000011001000001000001000110101110011011100001100001011111101010010;
#1 $display("%b", po);
# 1  pi=207'b101111011100110100110000000111000011111001001001101010110010011010010110111101100010111101000000010000101000111111110010000010110110010100010001001101011101100101010011101111010111000100000011010001010100110;
#1 $display("%b", po);
# 1  pi=207'b111011010100011010000111001110110001000110001100001011000010100111111101110001100010001111001110001101110110100001011100110001011010011011010100010100110111111010110111111000100001000001100010000111000101100;
#1 $display("%b", po);
# 1  pi=207'b101000001110011010101100111111000010111111111001010011011011100000010010001111010100000101001011011101110111110101011100001000101111010101000001111010101011110001101000001111001100111100000111010010100101011;
#1 $display("%b", po);
# 1  pi=207'b110111100110100000110001011010001000111011111110110001101101010101111011110010101011001101100101001101100011110011111110111011100111111101101101001101011001000111000010001101011110001100101111110000011100110;
#1 $display("%b", po);
# 1  pi=207'b111111100110110011110010100101111100001110000000101100001010110100010101101011110010000011111010011010010000111001010101101101011001100000101001110000010011110100011111011111111101001001010001010011000101111;
#1 $display("%b", po);
# 1  pi=207'b111100001011000011011111010010100011000110001100111010000111111011110000010001100111101101011001110101110111110101111110110110110001111101100110001010101100111011101011100000111010010100110110100000010000000;
#1 $display("%b", po);
# 1  pi=207'b000110110000101001011000000001110001000111110000011010100010010010111010000001110011001101010111011101111010000101110110000110010101100100110110001101011101010001110010110101111010110111101111101000111100010;
#1 $display("%b", po);
# 1  pi=207'b100110110100000000111010111100101110100010100000110010100001110100100110100111101011001100000000111000110101001010010111000010010000001100001001101000110011110001100011101100010000010001010011011100101110101;
#1 $display("%b", po);
# 1  pi=207'b101011101110101011001000001111001011110010111111100010100011011011000010101100010011100001001100100111110100000100000111001101101101010011001000110010011000000010101001010101111000011000010101000101000010000;
#1 $display("%b", po);
# 1  pi=207'b101111100110011001001111110010100010011011100011111001101010111000000001011001100001101000101010111001111101010100001101100010000110011010011000000000111111111101000111000100110100000010111100111110100111100;
#1 $display("%b", po);
# 1  pi=207'b100110100010100100001000101101010011000001010110110100010010010110000101011111111000010001111010101110010101100010001011110100110110000011011110001111110110011100110101100010011000110010000000111011010011010;
#1 $display("%b", po);
# 1  pi=207'b010010010010001100000110011011010100101101100011011011100010000010000100010111100111000110010100011011000110001110000101001000111000010000110000100011101011100100100000010010001000110001101100001010100010101;
#1 $display("%b", po);
# 1  pi=207'b001101011110100111001000111011111100011000011010011001101101000110101000010000100001001001110100100001001100101111010101010100010011011010100010111111001001000000011010011001101101001100100111000010101001010;
#1 $display("%b", po);
# 1  pi=207'b001101001101011010111101101111101011000010101110110001011101000011000111011001000101110100001011111100000010101111111110011001010000111000010000111001111101100010110011110011101101100001011010001110010011111;
#1 $display("%b", po);
# 1  pi=207'b010111110001000000011000001010011011101100111100000010000101011010101101101111100010000001010001011110000010010111001111000011100011001100010011001110001100100100101101001011101101000100101111111101010100001;
#1 $display("%b", po);
# 1  pi=207'b110001011010101000110010001000111110000110100011111111101100100000011101001000010011011101100110110101001011010110110001001000000111010111011010001101010111111101111101100001100100010100001001011011100001101;
#1 $display("%b", po);
# 1  pi=207'b000100000111111110001101010110110001100011010000000001110010000001000001100100111011011111100001011011011001000101100101100101101011110101100101111001001010111110011111000110111111010000111100010110101000001;
#1 $display("%b", po);
# 1  pi=207'b101100110010100100010010010100001100010111100100010001010000100100100001011111000011001110001110001010101000011010110011111101110101011111001111000100000111001010011000101101100010010110011001110101110110001;
#1 $display("%b", po);
# 1  pi=207'b001010011010000111000010010111001000010000101100100010011110010001110100000110101111001101011001101111110000011001101011100110110100110011011100011110001000000100110001110010110111011101001000011100000110000;
#1 $display("%b", po);
# 1  pi=207'b000001100000010011000001101110011110010010011100000010001000011101101110111011110110100001111111011010000011110001100100111000000111001001010111000111010101110100011010001111000010011101101111011111000111000;
#1 $display("%b", po);
# 1  pi=207'b101001011011011101101000101000011101010001010111010000100011111110100101100111100000010101110101100100110011000001011001110000100110011010101110110111110111110110011001101011011001011100001000011001010111111;
#1 $display("%b", po);
# 1  pi=207'b110101111000010100100001001101110100001011000111100100110110111100100000111011000100001101000100010000010100001000011001111011001011100000110100111101011000000111110101100111000010101111100000101110011100110;
#1 $display("%b", po);
# 1  pi=207'b010010000110100100111101001000010001111010010110010010110001111100001111010111000011111101101000000111110010011011010111011011101101101100111111011000100011010010000001111111100111101101001100000110110100100;
#1 $display("%b", po);
# 1  pi=207'b100100110111101011011100111001100001011001010110111001101100101100110010011101111010010100100000000100101001000011111011000111011111000100010001111111011110011101001110101111111011110111100001101010010101011;
#1 $display("%b", po);
# 1  pi=207'b011111110111010001101100011000110100110000111010011100110001001010001111010101110011011011111011010111101011100101010000110110110010000000011001011101010000001100110100010000110010101010101111001110000110110;
#1 $display("%b", po);
# 1  pi=207'b000110111000100100011010010000011111011001001101010100101000100011000001011000101101111000000011111001110011011001111000100000100001111101010001011011110110111101101111001110101110010001111111110100110010011;
#1 $display("%b", po);
# 1  pi=207'b011001110011001001100101111110110111011001011000100111010101011000100100001000011000011110010000011100100101101100011001110010111100001110111001011101111001111010011101100111000100110110111101100110100001010;
#1 $display("%b", po);
# 1  pi=207'b111011111100100100101000110011110001011010110000100111010100011110110000011001010111000001010010011100001010000100100010000100110100010010110001001101000101111100100000010111111011111000101111010111000011011;
#1 $display("%b", po);
# 1  pi=207'b111000110110001011011000010011001111100001111000101011001011100100011111110000101010101011100010000111001010001111110110010011110011001100110100100110000011110110001100110000111001011100001111101011110011101;
#1 $display("%b", po);
# 1  pi=207'b000000110001000001100111000001010000000101100110000010111100110110100001011111010101111111000111110000101110101001010001000010000100110011111001011100011011001101001110111000011011100111100100101010111100000;
#1 $display("%b", po);
# 1  pi=207'b101000110001101100010011001110011010000111001100010011010001101010100111001110001010111010100001111011001000101110111000111000000101010010110001011111100100001101000111111110110101001001111100000101101000100;
#1 $display("%b", po);
# 1  pi=207'b010101101110111110011001100000110101111101001001111010010010101011111011100111010010001011001111111111110100101011111001000110010010000101110001001011110100100111100001000010010111011100000000000111101011100;
#1 $display("%b", po);
# 1  pi=207'b010110101000010000011000110110001000011101110011010100111011100001111101010001111010100011000100100001110001010010010101110001101100101111110000100000110101100010101001111000010101100111111011101010001101000;
#1 $display("%b", po);
# 1  pi=207'b011010110000000010100110001000010101011000000100101100010101111001100001011010111100001111010011110100111010101110110100100011011101011100011000100100110000100110101001111000111010010010001101101110101010011;
#1 $display("%b", po);
# 1  pi=207'b000101111000001110010111110110111000000110010111000110101011101000111000111000011011101010000101000011110110011010101101001101011000000101010011101101000110101011101111110101000101100011000110110110101010011;
#1 $display("%b", po);
# 1  pi=207'b111010101101101101010010010110101001000000001000001100000111001000011010000110000010001011100100100100110001010011110010011000011000100011110001000110011000100010011101011000101100101010011000001011011110110;
#1 $display("%b", po);
# 1  pi=207'b111101111101110000110110001110011011101000000101000101110100010010101000001001110101011010000001110110010110000110001001011111111001110110011011111001110100011001111101001111001010101100000101101101110101111;
#1 $display("%b", po);
# 1  pi=207'b111110101110001000101011111010001010100101011110100101110000011100001100010010001100010110101010011100110100000000101101010111011001101100101100011011100001010010011110101010001011001001111111011011110100001;
#1 $display("%b", po);
# 1  pi=207'b000001110010001101011101001110001111011010111110100100010011001100001111100100110011101101000000110101110111010101111000010010000010101111000101110011110100110010010100001110100000110011111010101011011011101;
#1 $display("%b", po);
# 1  pi=207'b110011000011111100101011111101001110011100111011111100101010001100110110110101001000000010010110001000100010001001001011000011110101001100101110010111110101001100101100101000001001101001100101000101100101110;
#1 $display("%b", po);
# 1  pi=207'b000011111110011001001100000110101110000000110101111011011110000000011110011100000111010110011000010100000100011001011010110010010001001110100000111001010011010101100001001111110001000110011010001110001100111;
#1 $display("%b", po);
# 1  pi=207'b110000000101110011101010111100100111000010101011011001011101110000010000001011111100100001001100001100110110010111110001000001010101000101100110110001011101010111000100111001100101010111100101111011000001111;
#1 $display("%b", po);
# 1  pi=207'b000010111000111010101110110110010111000010101011110101111000101110100001011110111010000010011011000110010010000000011010001001001011010101111011010011010011001111000011111101001100011110010110100100101100100;
#1 $display("%b", po);
# 1  pi=207'b101011101111000101111100100011110001001110111101100011110100000000110001100011001011001100010001001111011001001000111101001000000100000101110011110010111101001100111001100010011001110001111000101110101010111;
#1 $display("%b", po);
# 1  pi=207'b000101100001001000001011110100110011110010010100000111000001100000110110110011001110101100011100110110010110010100100011111011101100100100100101100000001000000000101101100100110110111010010011101010001000111;
#1 $display("%b", po);
# 1  pi=207'b101111111111101101011100000101100111001110000010011101111110010111011100010110101111001100100101010100111100111110110001100110110010010101101011000000010010011101001100011000010111100110010011010011110111110;
#1 $display("%b", po);
# 1  pi=207'b001010101111011111110110001111011000111101010000110011111100100011000100110010000110110011010010101110111010101101100011011010010101010101110111001111101010000111101111011100101000001010110111011000011101011;
#1 $display("%b", po);
# 1  pi=207'b001011010011001000001000001100110110010100101110100001101100101000110011011001110011010100101110110111111110010000011100011110110000101010111101010010101000000100101011110100101101100011110101000000011100011;
#1 $display("%b", po);
# 1  pi=207'b111001000100011100100101000010100100100100100010110001101110100100001110111110100100100101000000101000010110000100100111111100011111101001101100010001010011000110110100100100111001110001111011110111100011001;
#1 $display("%b", po);
# 1  pi=207'b101100110110000111111011101110101011111111000101111101010101000111111110100100101000100100010110111011110101011011111111000001010001011000101001000001110010100100010110001001100111100000110010100011100100101;
#1 $display("%b", po);
# 1  pi=207'b111001011011001110010111011101101110110010011011011001101001001011101011110101000010110111010011101000101100010100001011110101001110111001110110111010000111010010011101111110011000110000100000100100000101100;
#1 $display("%b", po);
# 1  pi=207'b000100001110100101111001101111100011000010100010011011111011010000010110001110101101011010100111011111001000101100100100001110001010111100001100001100010001011000001010100101000101000001001010000110001100100;
#1 $display("%b", po);
# 1  pi=207'b100100110100110110000100110011000100011011010000100000100111010100001010001111000011011101001011110001111100011101011000101111101100000111011111101111001010100001110111110100001011101001001101101010101100001;
#1 $display("%b", po);
# 1  pi=207'b001000110101001100000110001110110010001010110000110101010101100101001101111001101101010101001000000010110100011011000111000011001101010010011000000000011011010111011011101010110010101110011110100001100100001;
#1 $display("%b", po);
# 1  pi=207'b100100001000010000100101010001010000000101110011000111001110011111011001001000101011000101001101111010111010011110010011001010001000100011110011101101000001100010010111000110101010100011011000000000110001001;
#1 $display("%b", po);
# 1  pi=207'b101010100100101111101101001101001000100011011110011110100011111000000110001111110101101111101001111110001000101101010110100101000010010001010110001010110001110010100110011011111100111100110010001110000111010;
#1 $display("%b", po);
# 1  pi=207'b000010100111100010010110110101110111011001010010110011101100110110011001011001101110001111011100010101100101111100110100101111110000100100011011110000111010011010110101111110001110100100100110011001101101110;
#1 $display("%b", po);
# 1  pi=207'b101000001101101001000000011111011100010111010100110101100010010000011110010101000000000010101101111111000000001111111111100000111110110101000011110111000110010010010100011101010101110100111101010111011011101;
#1 $display("%b", po);
# 1  pi=207'b100010101011001110101101111010111010110110100010001110111011110100111110100010001010101011000000010011110000110001000001010010000011000110111000001110100101011101111010101000111010011001010111000110010111111;
#1 $display("%b", po);
# 1  pi=207'b110100000110010001000100011000000111100000010010001011011001100111000110111011001011101010011101010010000000001110011110001111101011000110001000101110111100000000000010000110111000000010101001011101100010101;
#1 $display("%b", po);
# 1  pi=207'b011011101101000001010111110000011110011000000111111001111001111001011010101010000000010011000111001110100101101101011010001010000111001110010001001010101000110110100011100111000000101101000010000100101001111;
#1 $display("%b", po);
# 1  pi=207'b000101010111110001101101101101100000110011001111001110010111011100000000001111001001001100001000111000011100001001010000111111110100110000111101110101100100001010011001000011101100100101100011000100010111111;
#1 $display("%b", po);
# 1  pi=207'b011010111010101010010101001000010010101100111000010000000101010010000001000101011000100010000011011101010011000110011010011110010100011111100011110110110010110000110101110000000111101011000100000110110101000;
#1 $display("%b", po);
# 1  pi=207'b011110001001011101111000010000000010010111011010000100111101100000111011010010101000011101010000010000111011011010001011010110100101110100011010001010001111101000010011010101011001111101100111110100111001100;
#1 $display("%b", po);
# 1  pi=207'b001101000110110001100111011111110101001111110001011111101010110111100101110000000001011110000100111001111111010000111011110100110101010010011001001111111001100111011100000101110001001101010101100010100101010;
#1 $display("%b", po);
# 1  pi=207'b010101010100010101111010011101011000100001011001111110111111001001010011111101010011110001101111100101001010110101101101010001101100111001111100101010010000000101011110011011011110110011101000111110100010010;
#1 $display("%b", po);
# 1  pi=207'b100111110111110100001101000000011001111010110011111111010100111001000000010100001100101101000101010110000010000110010001101100010010001110100101111011011111010111011001111001010011010101100101101111110010101;
#1 $display("%b", po);
# 1  pi=207'b101101100111010100011100011110000010101100100011000011000111000001110010111001010000011000011101011010110101100001111000011110001110111110001100011010101101111001111100000110100111101010101011011110111111001;
#1 $display("%b", po);
# 1  pi=207'b010111100010100111110011101000011101110001111000111110111100100010011001011000100101000101011011101011110111011001001000101111111101111100100100000010001011101001001011111000001010011111011000010010100111011;
#1 $display("%b", po);
# 1  pi=207'b010111000011100011011000001110000010101101100100101010111100100101101010110001001101110000110110011000100001011111101000101000011101001111011101100011011111001010110100011101100111111111101101110101101100100;
#1 $display("%b", po);
# 1  pi=207'b100101111001100000010000011010001000010101100101100111110010111100101000111000111000100100111111100001110100001000011000101101000000000011111110001010101110010110101110100000110111100010110110001000111001111;
#1 $display("%b", po);
# 1  pi=207'b001100100100011010010111101101110000111001001100000001010100011100000111010100011000000010010000010011001011001110111110101000100111100101110000100100101101110101100010100011110010011010010011001010010011000;
#1 $display("%b", po);
# 1  pi=207'b001000010010101000100001110001001010100101110110011010110001001101000010111110001011110111011111100100010110100000000010101111100101111111100001101101000100000010111000001010111101011101001111010100001001100;
#1 $display("%b", po);
# 1  pi=207'b000001000110010000010111111101101000101110010111101001000011000010111100011001111101110111100010011001111111100100100111001110001100000101111110101000011010000111010001110101010011101010110011110000011001011;
#1 $display("%b", po);
# 1  pi=207'b100011101101011110010000001111101100000010001110111000010000100101101010100000001001111011010011110010010101011101001011110001011011110010110110001110011010110110101110100101010011011101000110111000000001110;
#1 $display("%b", po);
# 1  pi=207'b100111110101100001110000010110001001100010101000111100000100101000011011101010100000100010010111111111101011001101000110110101111001010000010010100111111010011010100010101110100000010011110000000111000100100;
#1 $display("%b", po);
# 1  pi=207'b001000001010101100101010011110000111111100010100000000001111011101000111100100001000011010010101011101011011001111111010110011011000000100010000001000001101111011100000110010000010110101001011011001101001111;
#1 $display("%b", po);
# 1  pi=207'b101011001110111101010010111011000111011100110100100100010000110001001110001110100111110011000001001011011101110100101101011100100000110111001001000001010001101111111101110100111010001001110010011010011101011;
#1 $display("%b", po);
# 1  pi=207'b010111011010000001100011001000110001100000000101101001111111000101111111111100001000111100000110011101110011010101010110100001001101100011000010010001000101111001010111100000011010100101100010110111101101001;
#1 $display("%b", po);
# 1  pi=207'b110010000101011011010011101100111110001101011111110110000100010001110101010101000110011101111011111001100101001000010110101110011000100100010100110000111101011111010010000010011111011111101000000000100000111;
#1 $display("%b", po);
# 1  pi=207'b010100101110101111000101001010110100011101101111110011110001011000110110111001110101100000110001000000011000010100010010001010001011101100111110001011100001010101010101110110000001111101110001011010110111110;
#1 $display("%b", po);
# 1  pi=207'b100111011001011010110001101111011010001011000101001000111011111100101001011111010000010110011011100100000111001111111111010110000011000110110001010011001001001000000010100111001111110010111100100110011101011;
#1 $display("%b", po);
# 1  pi=207'b001011010010110011100110111000011001101001011111110010111001100001111111011000000110001001011010110110001000000001001010101110111001101011101010110011100111010011111111110111000110011100000110101111011110101;
#1 $display("%b", po);
# 1  pi=207'b001110000001101010010100011010010010000010100001111101100010101001010000101100110001110001000010000001011011001100110010100111100111001011010011000010011100001001011000010011100100111100111011100001111001100;
#1 $display("%b", po);
# 1  pi=207'b001110101010110000000111001001011110001011000001001111111111100010100101011111000101011100001011000111000011100110101101011101100001010000011011000111000111001000011100010010101100101100110011111110001110101;
#1 $display("%b", po);
# 1  pi=207'b100001101011110110000001101000110101000011110000010101001100000000111110100101101011011100001100011100110110111101010011001100011101110111110000111111000001011110001110000111110100001111010001100100101110101;
#1 $display("%b", po);
# 1  pi=207'b000001101000111001100000011111110111110011111010010101100010111111101000110100000001101101010101100001001010000011001100111001011011101010011100000100100111010000000010000111000001001000011000111110101000111;
#1 $display("%b", po);
# 1  pi=207'b111001001001101111110011011100011011000010110011100010110101110101000111101000000010110001011010110110001000011001011101110111111110101111100110000111001000001001101010001010001001110011100001010110101000000;
#1 $display("%b", po);
# 1  pi=207'b110110100100011110100101110001011111000101011100110101001100000111100101000110101100001111110101011010001110110100001011100101000111100000010111000010110110011000101010011110111010011110010110010110101110010;
#1 $display("%b", po);
# 1  pi=207'b100000100000111011010110011000100010111100101010000100011111001001000100001010010101011100110111101000001110010111001001101101101110101101110011100110011110100010000001110101101101111101000011001011011101011;
#1 $display("%b", po);
# 1  pi=207'b110011001111001101111111000100100010110001111111101100110101000011111000111000011100010011100111011000011011101001101101101101001110011110110111000000001100110010101000000101100001011110101110001101001001001;
#1 $display("%b", po);
# 1  pi=207'b001000101101000010010001100000011100001100101110011101101101011000011010010011101110110000001011010011000011101100111011010111111111111101100101100011100110101110111111110001000000000010001001011111110011001;
#1 $display("%b", po);
# 1  pi=207'b100010100101010011010111010101100100011101010011010010110001001000001110100000110110111001010110110111110000000000111111010010111101100000111001010100100010111010100011101011100101100101011101001010011000011;
#1 $display("%b", po);
# 1  pi=207'b100110100100001001101111000011010100111101001100001011110010111000101011000100100101111000100101011010001001110111010101101011000111001001010001000011000101001110110011100111100000111110000100100110001111110;
#1 $display("%b", po);
# 1  pi=207'b110110011110101001101010101011010100110110001111111111010110001111010001011111100111100010001100101011101101100010100010011001100000100111000111111001101110000000011111100110011010010010110010111011000111000;
#1 $display("%b", po);
# 1  pi=207'b001100111100100111100101110101100110001101101101010011000011111001001000101110000000001010011011010100100001001100011100111001111101000001011101111110101110011111011000000111110010001110010010100011110101100;
#1 $display("%b", po);
# 1  pi=207'b001110000101010001001010000100011101110100010011010001110111101111110001011011000110111110000001111111110011011101011011110011001101101010010001011011111110001111111010010101000010001101000110101001110001010;
#1 $display("%b", po);
# 1  pi=207'b001001111110001110110000000010110011010000011111101000111011110100010001110001101110110111110101000110001011101011110101011010111101010000100011001101100100101001110100011001000010110110000110000001001110011;
#1 $display("%b", po);
# 1  pi=207'b110100110001000101001101110000001011101001100010110110001000001101010110010110011101001101000111100101101010000111001110001010001100011010101101110111101000011100011110001010000011000011111110010101111001100;
#1 $display("%b", po);
# 1  pi=207'b111100110011100010101011111111011000001011101100110011101110001111001111011001111111101010111011011001100111010000011000101001110111010001110100110110011000010101111001100010110001000110111010110000101110001;
#1 $display("%b", po);
# 1  pi=207'b110110001001001000000111001000101100111101101000101001010100101110000000100010111101010011010001111001111111101110100111100011101000001000011111011110110101001001111001110110011110111111011011000010001100001;
#1 $display("%b", po);
# 1  pi=207'b101100001011001101100010001011101111110001100001101100010010110101000001110011101100111010110011000011101011000110000001110010001101010000001100011110001010111100111100100010111000100000000000011010001001010;
#1 $display("%b", po);
# 1  pi=207'b001111100101001111101001001101100110011110000010001011001001100011111011000101101100000111110101000000000101110001110100001110011110101011000000011011000101110110011001110101011101101110011101011101100111110;
#1 $display("%b", po);
# 1  pi=207'b110000010111000111011000010000110010010010011001110010111101100101100100101010010100111011100110101101001101110100110101111000101101001110110001011100101010101010111110111011100001000111000110000111010010110;
#1 $display("%b", po);
# 1  pi=207'b000100000001110011001110111011000100001001001111011111111000011111000110010000110110111011001111000100010110000111110000110101110101011101101001100111111010101001110100101001010100010010101101001000111000110;
#1 $display("%b", po);
# 1  pi=207'b110010010001011000101000101110011001100000011111100001100101011100011000100001111101110101010111011110010011110110000001001110010101011101001100010010110010011001001010000010101011100000001001111101111101101;
#1 $display("%b", po);
# 1  pi=207'b110011100011100001001001010011111100110000111110110010111100110110101011111110111100110110111111010010010100011111010011100100110011101100011111000111011101010110000010100100011001011101001110001001000001110;
#1 $display("%b", po);
# 1  pi=207'b000011000110000110000100101100000111100001100000110101101111111011100010011110010001101000010110100011010010000110110010000111010101101100100011111010110001110101100100010010111100010110011100111000011100110;
#1 $display("%b", po);
# 1  pi=207'b101011001001000111011000010101010110001000111001011001111110010100111111110100010010111010101011000100010111101110111110100001100000110001111000111100010110100110111011111100001111110101001110110011110010011;
#1 $display("%b", po);
# 1  pi=207'b001001000001010000000110011011101100001110010110010010111000010111010101011101101011100001011010101101100110100010101101001011100001100000001101110100110110111000111011111000001010011110101001000110011101011;
#1 $display("%b", po);
# 1  pi=207'b000110100011011000100011011000001100010110000001111010101100110000111010110110001001010100110111111111011011110111100101010101101011111011011010110010110100010000110100111000001010001010000101111011000101111;
#1 $display("%b", po);
# 1  pi=207'b000010110011101001001000010111100010000001011001110101110110111001001101011101001011110000000011011011101111101110110100001111000001101100010011101001000101001010011100001100010001000110100011101110111110001;
#1 $display("%b", po);
# 1  pi=207'b010101100011101111011001111111001011110110001101100010000011111010001011000001011000010101110001111110010111001100110101101101110001101001011001101010110100011000000101101001001100111011010110011001110111101;
#1 $display("%b", po);
# 1  pi=207'b110011100000111110000001010011110110010101000111100001010111111101101101011010101000000110001010110111010001010100100110000110100111111010010101000000001011001100010010001001000000001110000110111100101010001;
#1 $display("%b", po);
# 1  pi=207'b101010110111101110011010011011001010000101100010001110101101110100101111010010100011001110000010100011001000110000000010001101010001110101101010010001100001110110110110101011000000000100011010010101010100101;
#1 $display("%b", po);
# 1  pi=207'b101101110100100011101110000000001010010110111000011111000000001101101101001101101000111111110111100011101001111111111110001000011110001110101111010001110110010010111010010010001000110001111000001000000010101;
#1 $display("%b", po);
# 1  pi=207'b010010110110110101010101111101001011100000011100011010100111110000011111101111010100010001100001101100001100010000001001001001001010001011111001101010101111001111011101010101010111101110010111110011001101001;
#1 $display("%b", po);
# 1  pi=207'b101110101000001011101101011110000001000000100101011001010011110111010000111001010011000010011000000100011001011010110001101011000101101000010101111001001110010100000111001110110010101001011011010010010010010;
#1 $display("%b", po);
# 1  pi=207'b110111101110101111110001111000010101011011101001101011000011011001110010111110110001001010000000010100010110001011111101101110000110000011101001001100011001101110101001101100111000000011000111001100010010101;
#1 $display("%b", po);
# 1  pi=207'b101010011010011110110001111000110010000001101101111011001000111001011001100010101011010011001000010000011110101001101111000100100011000011001110010110001110101111010111110101111011000010111110100110110011110;
#1 $display("%b", po);
# 1  pi=207'b100100000010100111110100101000011001111111011000111000100010000100010000100011001000101101100011001000010100011111111100010101101000110100110011000111000000100101010010001000001111001010111011100111111011100;
#1 $display("%b", po);
# 1  pi=207'b001000111000101001110101100110011010011100111100110000011000010011111100001000100110100000111110110100000110111100101100100101011011011001111000010000100001000110011101111010010011111001001001101001111111110;
#1 $display("%b", po);
# 1  pi=207'b001010100111001010001100011001011010000000011011111101000111101101000110011010110111110100110010010001110100111110011010100010111101110001011110000100100000001001010010001110011101111000100000010111100011101;
#1 $display("%b", po);
# 1  pi=207'b101110010110100010000000011000111111001100010010100000011011000000010110000010111101111001110101110011111011111001011010100101010110001000100100001101100100110000011001010000100100000100101101110011110000001;
#1 $display("%b", po);
# 1  pi=207'b111110000101010100011110000011011010001110100111101100001111001000001110000000110101101000111100110100101100100001111010001110000001110111111111010110110110000010010111100000000101111111000110101001011000101;
#1 $display("%b", po);
# 1  pi=207'b110100011111111100111010001100011000101101011000111011011011110101111001011011011001010010100001011101000011011101001011101011100010111000001111100001001110010100001111111101110011000010101111110000010101011;
#1 $display("%b", po);
# 1  pi=207'b111001010011111111111011001111100011010100101110011100100000110010101110110101100110100110101100100100111100000001010100111001101111111001011100110100001100101000010000101100010111000010010010010011001111110;
#1 $display("%b", po);
# 1  pi=207'b000100100111010100001001110001000110010001011001011101110011000110000111110011010101000001011111001010011000110011110011000011101101001010010011110110001100000101010000110101110010101001011010100010100111110;
#1 $display("%b", po);
# 1  pi=207'b001111000100001111101000101100010101111110000010011111101111110000110010100110100011100001011100001010101000110101000100010100011010000101000110101100101011111010111001101000010110111001010100101000001000011;
#1 $display("%b", po);
# 1  pi=207'b110010101001111100011011001100000110110001010001001011001111011011001110010101001111110110001100011001001010010010110010000010101100101100010001100010010111010010111000000010000110010001111101100100000110101;
#1 $display("%b", po);
# 1  pi=207'b110001110001110101100000101110000100000110001010000101011010101011010110101010011001111000001010100000010111000010000101100011110111100011001000110110111010101111001000011111101111111000100100110111100101011;
#1 $display("%b", po);
# 1  pi=207'b000110110111000110111101110111000001010111110011011011010011101110000100001000100010110010100111010100010110011010011001100001110010110111111111111001111100101110101010000000101100000000001000010000001001101;
#1 $display("%b", po);
# 1  pi=207'b101110110011101111011011001110100010100010000111010110000101101011100100011110100011111001001011010010010101101111110101010001111100001010010011110111101010011111001101100011100011111100011000001010111010101;
#1 $display("%b", po);
# 1  pi=207'b110000101010010011001111110101010001101000011111111001110000001010101010010011011110100100110111000100101110011111100110100110110101101000100010000001101111111100101110001100100000110110111101011000101100110;
#1 $display("%b", po);
# 1  pi=207'b010110100110001111100000001111010110011101101010000111001001011101011010000100001110111100111010011100111100011000010100100001100010000101110110010110000000000001010010001110000001000011000110100100001110101;
#1 $display("%b", po);
# 1  pi=207'b011110001010000010111100111001100001001110000101000001101000111111101100111101111010000100011101001111001111000111110000000101011111001110100000110110010110000110011110000111010010001111010110001110010101001;
#1 $display("%b", po);
# 1  pi=207'b100011110000000101100111111110000010100010100110111010010110001110000100010100010111010000011011111111011101000110001111101011110000100101010011010011010110111111011100101001001110101001010110101100000010110;
#1 $display("%b", po);
# 1  pi=207'b011010110110111110110100011110010100010111011110100010000111101001000110011001001110110100001000010110000101011011110101110001110100100011000101110111000101100001110111011001000011000100001110101110110100111;
#1 $display("%b", po);
# 1  pi=207'b101111011100101001011010000001010110011011100000111100111110110110111001100101000100111000110010110101010110000011001101010000010011110001011110001010010111011011101111001000101010111011000010010000011111010;
#1 $display("%b", po);
# 1  pi=207'b110110101000110010111110110011011010111110100101100010111001001110101111010001100101010110100000001001100001001011001100010111100111111011100110111101011001110011010010000011101000000011010010000111011110011;
#1 $display("%b", po);
# 1  pi=207'b111010111101110101010001100111011101101100001010111000100011010001011011010000110101001111010101101100110001000100110010001010000000100011100001011011001010110110100000011001011101000100101111001111001111101;
#1 $display("%b", po);
# 1  pi=207'b001001001001100000100010100101101100111001000111010010111101001000000110000000101110101111100100001011110011101101101010000110110100000001100001100000111110110011011111101101111100011011100100110111110011100;
#1 $display("%b", po);
# 1  pi=207'b100101000010110010110111110110001011001010011000110011100000100000100111101000011010100110001001100100000010110010100011010000110100101111010010001000001010101110011111011010111101111011001010110001100000111;
#1 $display("%b", po);
# 1  pi=207'b000010111100111111110000101000010111000011111011100001111110101000100010001110010111111011101100010000100100001011100010000110101100010100101111101000000101010001000111111100111000110000100100110110011101000;
#1 $display("%b", po);
# 1  pi=207'b010111101010100111101010101000010010000101001011100110100010110010001100101011110100000010001111001001010100000110110010010101111110010001010111110010010101100011100110000111010110101100010000011110111011000;
#1 $display("%b", po);
# 1  pi=207'b001110110100100111010000100001000111010000101111001001101101001000010001001000101011110110010001100100100110010100010101101101100011000000011001001010100011101010001100110111101100000001101001101001101010110;
#1 $display("%b", po);
# 1  pi=207'b011111101111101100111101100111110011010010100111010001001100101001001000100001100100101111111001101010010001001001010010111110011110101000101010111010101111001001000111110100000010011000001011111111101101110;
#1 $display("%b", po);
# 1  pi=207'b111011010010100011000010010011100000101101110010011110101111010001010111111101111100101100001001000100011101100001000010101111000100010010110101101111001100100111011010001000010001010100101010110110001101110;
#1 $display("%b", po);
# 1  pi=207'b100000101000001111101111100001011011001110010110010000011010110100111001010000110100100110010011111000111110101011110000110101011100101000011110110111100111111010100001100011001111110110100001001101101010101;
#1 $display("%b", po);
# 1  pi=207'b001110010000010010000101000000110011010001111000111011001111001101110001011000001000001011100110001100000110111110010011001100010110011101010011110111010001000100101101100100011000010001110110000000010011101;
#1 $display("%b", po);
# 1  pi=207'b001101110101000110100101011111111010100011110001011110011010010110000101011110010101011101010000100000110110011111010101110010010111110100101111111011001100010010110100100111111100001001110111101101010111111;
#1 $display("%b", po);
# 1  pi=207'b001000111111010011010000011000000000100100110111100111101000111000001111110101001011010010001111110110101010110110001111001010010001000011101001000111101010000100011001001110011111001010000110110111110100010;
#1 $display("%b", po);
# 1  pi=207'b001010101001000100110010010111000110000111110111110100101000000111010101110010001100100001001101001010110001010001111101001000100111100100101100111101011000011000110011010011110101101001001001101001010000011;
#1 $display("%b", po);
# 1  pi=207'b111111010001011100110111101111101011010000000110101100010101100110110001000000000001101100010011111001001110110101111001101010010011011000101111100100101001011001001101000110111110110100100100101111111111011;
#1 $display("%b", po);
# 1  pi=207'b110010011101000101110110110010010101111010110100011110111011001011100001101000110101110010011110100101110010001100001011111010010000001101010100100000010001000101001110001000010000010000010111001101010010000;
#1 $display("%b", po);
# 1  pi=207'b000101001001000110010011101110000000100100010110100111001001101110111010001111001011001100111101010001110110110110011010010111100101010010001001101010101001000000011010010000001110110001111010001000010000010;
#1 $display("%b", po);
# 1  pi=207'b000111110101110011000010010011101000001001100100110111001101001001000101011100010001111111110000000010010010011010111111010011110001011000100010101101100001001110010111101001101001100011110011000010101001101;
#1 $display("%b", po);
# 1  pi=207'b100010011000010001011010010110111101100101111110100100010100111100100101110110000101100001101110011011101100110010001111111001110001011011110111110111111010011010010010110011110110100001001001110000001000111;
#1 $display("%b", po);
# 1  pi=207'b010010100001000011101110001111010010100000100000001101101011110010010100100101010100100011100000010001000001101111101010111100100000111010010011000111101101101001110101000110101100101101011010001001100000101;
#1 $display("%b", po);
# 1  pi=207'b101011100110011001111111000011010011111010010101100110001101000001100011001011111011100111110001111110110011100001111110010110101011100001100100011100010011101010001100101011110101001100111000011110100010011;
#1 $display("%b", po);
# 1  pi=207'b001000101110011011000011101100000111000011011101100100101011010000001010110110111001001110100100001010011101110100011000101111011111101000000110111000100000111101011010110110101001100000001101010010001000101;
#1 $display("%b", po);
# 1  pi=207'b111110010111001101101010010011001010100000100111111000100001101010001000001101110011111100101011011100100001011000001110110010100101101100001000110100100101001101001101001010010010000101011011110000110100001;
#1 $display("%b", po);
# 1  pi=207'b100011011111000101011101101011010010110101000100001010000011100011111010101111011000111011110101011100011101100101101010010010110101100010100101100111111011111011111000011100111010111011010001000010100100100;
#1 $display("%b", po);
# 1  pi=207'b111010110100100011011011011011011100110100101100101010000110011000110111000101111111111111100001110111011000101111110010001101111111101010010111001010100100000001101001101010010010101010010110010011010001011;
#1 $display("%b", po);
# 1  pi=207'b101101000100111001110101111111101010010110111110110010111010000001101101000010110001100101110001001100000010000010101001100101111111010100110001011100011111100000011101010100011000100101101111110100110101100;
#1 $display("%b", po);
# 1  pi=207'b001110101101101110010111111101010010111110110001011100101011011111001000010110011001011101100111110010011100111100110011110100100011110100000010100010010010011001011011100010111110010101001001010111010011000;
#1 $display("%b", po);
# 1  pi=207'b000010110011011111100111000010010110101001001000100010111110001100100100000011001001011111101001110010010000000111000101010101010010011100100010100010101101110100110111010101100111011110000000100000100100111;
#1 $display("%b", po);
# 1  pi=207'b011101000101100011010100110111000100101010000010001111000101011000101111000011110111111101010000010001100101111101101110111010010000111010011010011101111101011010001010001010001100100011011111110011010111000;
#1 $display("%b", po);
# 1  pi=207'b101110100101110001110101110000011011111001101111000111010110011010101000111111100101000101001001011010110011110110110011010111000110101110001001001001010011000010011011110100001011001100111101011101000010000;
#1 $display("%b", po);
# 1  pi=207'b010010000111100111011110110110000110110111110000000110001100110100000010001111010010111001000100101101001111110101011001000011011111111100110000100000101111111000010001101101001010011110010010110100100110011;
#1 $display("%b", po);
# 1  pi=207'b110010001011100000000011101001100001010001110111100000101111111110011001100110000011010010000100111101000000001010000000000101000000001011010110011010000001010100000001011110100110011110000110000110001101011;
#1 $display("%b", po);
# 1  pi=207'b001110100000101001001001001111100000000011101100011000001110000101100100111100000110001001100111011010011100010001000000001110111001010010100101100011010010100001111100000100001110000100101001111011011110101;
#1 $display("%b", po);
# 1  pi=207'b000010110111100001100111011010101111000000110011000110101101010101101100110000101101101100001000011010101001000100101011011111100100010101111001100110010011000110011001100001001100010111100100100101100001110;
#1 $display("%b", po);
# 1  pi=207'b010010100111010001100110111110100010001100011010100001101111010001001001010111111001000100001000001011110011001111010011101110001100001100000111000010100111110001001011111010011010100000001101111110111001000;
#1 $display("%b", po);
# 1  pi=207'b101111110110101111101010011100000010111110101101111100001000100100000011000001110100110111110000101010001001001001001111110100000111011001000111011101000000011011001100101100111110001000011011110101000111111;
#1 $display("%b", po);
# 1  pi=207'b101010111000011111110000001100111010011110000100000101011000010000000110100101110011111110111001010010010011100101000010000110101011110100000000110111111100011010010001011000011101110110001001111111000100011;
#1 $display("%b", po);
# 1  pi=207'b111110011010010001000100110000111000100110100100000010010101111111110010101010001001111001010011101110110101011011010010100100000110110010001001100111111101001111110100100011110011011011000111011101111010111;
#1 $display("%b", po);
# 1  pi=207'b000000111100100100000111010001101111100000110111000110000111100110100111011110100111001111110001010101001010011000001000010011001110100001101111011011110011001000110001011011011100010101010111111011010001000;
#1 $display("%b", po);
# 1  pi=207'b111110100111101011110001000101101001011011111100111110101011000011110110001000001101000001101111100010100001111001101011000010100011010111010011100111101010101101001101100110011110010010000010001110101011101;
#1 $display("%b", po);
# 1  pi=207'b010011100110001100100000100010100110101000001010111000011100100001101011010010110010011001111100010110110000100000010011110100011111110011001001111110111001110001000100111011000011111110101001011000100111010;
#1 $display("%b", po);
# 1  pi=207'b001100000101101100111000100100011111101011001111010101010100101101000100110110100011111111010111101000010000000100010111100001001111001100110000101010000000010111011111010000100101011011011001111011101000011;
#1 $display("%b", po);
# 1  pi=207'b001101100101101101111110110000111011110101110001000001000001111110110110000110001100111010100110011101111100011010100100010100110101010100010000001001100101001110111100010000010011110001101010011011110111001;
#1 $display("%b", po);
# 1  pi=207'b111000010101010010001010100110010101101100110111101101100000101101111110111010001111000010110001111001101000100011011011001101011100110000000001010101111001000111110111101010111001011011101100001101011110011;
#1 $display("%b", po);
# 1  pi=207'b010110010110110100001001010001111001011011100000010110011000000101100010001000001111011010001011111001010110110010001011100100111010001011001110111000000101011111101111100010001010101000000100100100000101000;
#1 $display("%b", po);
# 1  pi=207'b110011001000010101011111001110100011001100000001101111011101011000010110101010011000001101010011011110111000101100000000100010100010011111110110110101011000101110001101000011011011010011111101110111100011110;
#1 $display("%b", po);
# 1  pi=207'b111011011100100101110001111110111110110000100000100111001100101001110111110101101111011010001110011001011010001100011100111111000000001111011101101011000011111010011010010110101000011111100010010100010001101;
#1 $display("%b", po);
# 1  pi=207'b011011111111010001010100101001111101101010101111110000000110011111111101001000001101000001001111101011111110000010111111011010101100011101010010000110010010011101110011111110010101100001110000100000110011100;
#1 $display("%b", po);
# 1  pi=207'b010011010111011111010011101100111010000011011011111111000010001111111010111111011000110001101111010000010111110011101101100001101001001101111110110101101001100110110010100110001101001100011101001111100011001;
#1 $display("%b", po);
# 1  pi=207'b101101011010101111101001101010001110110100101001100011001000010100000110001001111111011111110101100110110110010001000001100011101101111101101011010010010010111001100011101001011101001011101011100111100000011;
#1 $display("%b", po);
# 1  pi=207'b010101001011000110011010000100000011010011001101100111001111101001110010100010000011011101001001100010011010011100110001011001111011010011000100011110101011100011001101101001100010101100101100010110010011010;
#1 $display("%b", po);
# 1  pi=207'b100101110100001011100100000111101000110011001110101011010111100110100100001101100111010111100101010110100100110111011010011011111000110011011100111001001110110000101110100101000001000101100100110110111010000;
#1 $display("%b", po);
# 1  pi=207'b100010111010000010110010010000010110101111100010101010111111110000001000000000110000000110011100000111011001001010010101001010110011110010100000010011010111111101011010101000010011100100001101000001010000001;
#1 $display("%b", po);
# 1  pi=207'b111110001100011111000001110110101000000001100111111000000100111101010010111011101011001100001000000000001101110101110010101100011100111110000111001101101011101101100110011000110111111001111001101110101100000;
#1 $display("%b", po);
# 1  pi=207'b000111110110000010111011100100010010110111110000000111100011011000000001100110111001110101100101011110111001010101111110111110011010110000110101010011101111010100110110001100010010101010101110000111001000010;
#1 $display("%b", po);
# 1  pi=207'b011100101010101000010110000101100101110100110101100101011111101000100100101001001001101100111111010010011001111111011101111000011001000110110101001110011011001101011011011101001001000110001010101111101100011;
#1 $display("%b", po);
# 1  pi=207'b010111001001110010110001100001010101101100111011100101010001011110100101011001110000110111101000100111101111100110101101001010111111101000111000100110011001110101100110001010111000011101010011111110000011000;
#1 $display("%b", po);
# 1  pi=207'b110001001110111001100110100111010100001111111001100000100001111100111110001110011101100101001010111001101110110001110111011001110011100111000010001000001101011001001010001101011110010101000111000011000100110;
#1 $display("%b", po);
# 1  pi=207'b001110010101100010001010011111000101111000011100100001000000011101000111110101100010010101100000110010101001101101000100011110000100101011010110010001110101000001000000111110111001111101001101010011101010100;
#1 $display("%b", po);
# 1  pi=207'b110001011101110101010100010111001010101110111101010001000010010011110111111100100000111010100000000110000110000010000110101110011100001000001101100101100111011010111100111101110001000111110001100000110100111;
#1 $display("%b", po);
# 1  pi=207'b100010000010101111010001010111010001011011110110000001011001001100110000001101100011110010101101100101111110000000101001011001000101010001110100111001001001010011001010011110100011001110111011001011010110010;
#1 $display("%b", po);
# 1  pi=207'b011001011101110111001101101100001000110111101010011000001110111100000010011010110010111010110010101000110001010001000000011001110001110010000010101001011110011111101111011111100011111010001111110111111100100;
#1 $display("%b", po);
# 1  pi=207'b110100001010101010011101000100110110000010101011101001101101110111011101110000111101011100110011101001011110011100110010101110101000100011001001011001011010000010000111110110101111010001011011001001000101101;
#1 $display("%b", po);
# 1  pi=207'b111110000011111011110011111111110010101110010001100101101100010101000110100001111101110101001110011101011010101111100001111010010001011010110000110011000100111110111111100000011101001110101000111111101011111;
#1 $display("%b", po);
# 1  pi=207'b010100100001110110001100000001101001110001110101111010110100011110101000000001011001100000011011110111110110100111100010011111000100100011110111111101110111111010111110001011000011000110001001100011100100011;
#1 $display("%b", po);
# 1  pi=207'b100010111010100101111101000101100111101111101111010010101011001101100100011111010111010101000011111111110011011100111110001101011011001111111110010110111001000101001111000010110010111101001011110110111100000;
#1 $display("%b", po);
# 1  pi=207'b001100011010110111101100110100011011000110101111111110101000100001011111001100010110101110000000001010000101010111010000010100010010111110111010000010100001111001000000010000111101011010001111010010000110011;
#1 $display("%b", po);
# 1  pi=207'b100010011100111001001000101100011111010111011101110001000000011101011100110000010001010101011100100111111010111000101000000011100100010010001100110101001110000010100011101100010011101011011011101101101101001;
#1 $display("%b", po);
# 1  pi=207'b100001100011110000101011110011001100000011010100101010100011111010011100011000011001100001000110111101010100101001000100000110011100001100000011101011101010100111101101110100010001111000001111011010100011101;
#1 $display("%b", po);
# 1  pi=207'b010001110101111110111001111011100111101110011101011011111001011101000011001100011110011011010011000101011111010111010011001110001110111001001000110111101110011100001100001111010010100101010101101100111010001;
#1 $display("%b", po);
# 1  pi=207'b010110001010110100010010001010111010010000110001111011001111010010111101101100101101010010010001001000111010110010101110101000111110010000010010100111100101101110001110001110101100011010001111100000111111110;
#1 $display("%b", po);
# 1  pi=207'b111100101001011001110101010010001010110111011101100100111001010100111111110101001110101111000100001011101111010010111110110010000110110101110000101011100000101110111100100001010010010111000000001110100011010;
#1 $display("%b", po);
# 1  pi=207'b101000001011000000001001111111110010101000011101010011000101111101101010011010000100101001110111001110100010001101111001001101001001111110011001111010101010001100111100001010001110000101101101011100110001101;
#1 $display("%b", po);
# 1  pi=207'b000101010100001011001110001010110010010001010010101001001111001111001111110101010011111011110001100111000100111111111010111010110001110111100110000100010000100010101100101010001001000110101001110010010010001;
#1 $display("%b", po);
# 1  pi=207'b100111101111000110001111010011011110110111100101100000100111100000110110100110010101010100101000110011000110100001010001011100010001100000000110010101110110001011011110000000110000001101100001101011001000011;
#1 $display("%b", po);
# 1  pi=207'b100000101100110011111101001001000110100010110011111111101001111111111000100101111101011100100001001111111110010011011000001111110001000011001100100001011000011110111110011001100010110000101110111010111110010;
#1 $display("%b", po);
# 1  pi=207'b101010111011101100010001110111101101100101010010000110001001110111110110101001100100101001010001010010101000011010111000110111011001010111000000001011001110111100110000011000101000010011100001101011011101000;
#1 $display("%b", po);
# 1  pi=207'b000000100101010101100011100100010000000101000101100000111011110100101101101001000101110101110110001000000100011111010110010111001010100101111110000000111100111010000110100111101000010101000011101100001001110;
#1 $display("%b", po);
# 1  pi=207'b100000110111110001001000010011110101100101010100000100100010000101001100001010111000101110000101011010110000010111001100110010111101101101010111000100011110100011111001001010110001111000100011001011001010111;
#1 $display("%b", po);
# 1  pi=207'b100011111011100001101000010011101111011111011011010000010101011101110001001101000100010011010110111001001000001010110100000111010110011010110111000111001101001100100111101101001001011111010011011101011111010;
#1 $display("%b", po);
# 1  pi=207'b110111010000000110100100011010000011101011101101111000001110000111101010101010010010010110100010001011011100111100010100011101111011011000101010110010110001100100011000011100000010001101111010111011111101101;
#1 $display("%b", po);
# 1  pi=207'b111010010110111100110010011101101101101100111100010001001011010101111011010010110111101011110100011000111001010100100100001110101011010100100111101101111111010101000001010110101010010010000000110000010100010;
#1 $display("%b", po);
# 1  pi=207'b011110100111001010111000101100100111001011001100111111011001010100011101101001101101011110000100101100101111111111110000010111100100101111000001010100111101111000101011101100111001011110010010110111011110100;
#1 $display("%b", po);
# 1  pi=207'b101111101111001001101110100001010001010111001010001101011110001110000101011011000110000000001100011111010110100000000111100010010111100011110101100110101111100101001101000101111010101010010011001001111001111;
#1 $display("%b", po);
# 1  pi=207'b010111010100011001001000010100100101101110111001111101101100101000101100011010011100111001110011000000110110001101011111011000100011110011011010110111010001100001100101101111111001110100100010010101011001111;
#1 $display("%b", po);
# 1  pi=207'b111011000011101001111001000100011000011001010100011110101101000110011101101101010011001001111011101101111000000001011100101001011110111001110000100100110011011000000100000011100100001101110001001001000010100;
#1 $display("%b", po);
# 1  pi=207'b100001111010010010100001100110100010110111011100011011111100110001100010000011100111101011010100001010101110110000000110100011101101000100110100101110000010100000011001100011000001010100110001111101101000110;
#1 $display("%b", po);
# 1  pi=207'b010101011100110011000010110100001110111010100110110101011011100000001000111110000111001111110101111101001000010011111100010010110110111001000110010000111010000000101010001011101101100100010101110010000000011;
#1 $display("%b", po);
# 1  pi=207'b000011010000111110001101000000001111011010110100110111111010010011010001101100101000000110001101010001010000100010010001001101101000000100010110111111110100100011011011111010101110000011101101100101110100001;
#1 $display("%b", po);
# 1  pi=207'b000100101101111100110111110101000010000011101000111101011010100111001100010100011100101100110110001110100010100100100000000001110110110001001010001100111010001001100111101110000100101101100101011111000100000;
#1 $display("%b", po);
# 1  pi=207'b001111101110101100011000011111110100111011010011010011111101101101000001110011100010110010111001001101100001000110111101101100110010000110100000110001011101111111000100111000001000001011101101110010101110010;
#1 $display("%b", po);
# 1  pi=207'b111100110110100000101010010100010111111100001111000100110011011010110100011001000001001110001010101100001101010011001111000110111111000100011101111110001111101110010101010101000000001110110101110101000011111;
#1 $display("%b", po);
# 1  pi=207'b111001110000101110001110000001100100100001101100101011101000011111010011101111100000111010001010101110000001111010100001101000001011111011100100000011010111101100000111011110101101000010101000010000010000001;
#1 $display("%b", po);
# 1  pi=207'b110101101001111101010011001000010100010011011001000101100101010111101000111100111011101011110110110011000100011000010011001011110110110110100101001100000100110000000010101011001100101011000111111000011001000;
#1 $display("%b", po);
# 1  pi=207'b110110010011100100010000111011010110011000010100010011000000110110101100011011000010100001110011100100110000111011110001110100001111111101110000100110100100111010000011111111000110001011110100100011100011001;
#1 $display("%b", po);
# 1  pi=207'b011101010111011111101011000111011100000111100110000010010000110100111000110111110101010101000110010000100100111000100001000110100010110101011110111011000101000011101011011000001100011111000011111111101000000;
#1 $display("%b", po);
# 1  pi=207'b111101110110100000010011101111101101111111010111111001110111001111010001011100110010001100011011111111100000010111110011011010110011000111001001101100000100010100101100111000011001010101111100110011010010010;
#1 $display("%b", po);
# 1  pi=207'b100001100100010010101000010111110110011100111111101101101011000101010010111010111000000101000101000110110101100111111111001110001010111100111001100111001001001011111110101110101100110000110100010111101101110;
#1 $display("%b", po);
# 1  pi=207'b011101101011011100001001101000000011100100111000100000001010110011001000011000011011100100100001101101001110101100110110101000101010011111101011010111001100000010000000110100111001111001010011111101000101011;
#1 $display("%b", po);
# 1  pi=207'b110100111101001000011011100110011111010101011101110100010110001001010110101100101000011010111110111001110101011010010100101010001011001010001000001011010110010011100101111000000001110111111010110001001101100;
#1 $display("%b", po);
# 1  pi=207'b110100101110010001001010001011111000001100010000110011110001100011010110000100111110111000000110000110010100110000001000000011101101000111010101101110110010110011011011000000001111001101110100000101111110011;
#1 $display("%b", po);
# 1  pi=207'b010011110110001101100001100110111010101000000000110111000000101111000101110011110010010000110110001101100111101001110110011000011110001110010010111110000101100011110001110001000000110000010010101100001101001;
#1 $display("%b", po);
# 1  pi=207'b010100011100011100100001010111111110101100011010111111110010000010111010000001011000100111000111111100111001011100010111101110100101010111011010100011010110010010111100001000101110000111101010000011100010000;
#1 $display("%b", po);
# 1  pi=207'b011010100101010100111000110110010000000111110010001010000000100010100100111111111000010011010010010011000100011100100100101100010001000001010110100010111000011000100101011000011101010010111100010010011011110;
#1 $display("%b", po);
# 1  pi=207'b111011110101110111000000010110110001111010110011011011101111110001111011011011000001001011111100111100110011001010100100110000100001000100101101111001110010110111111001110101010101101000011101010011000101001;
#1 $display("%b", po);
# 1  pi=207'b001110001000011110100110000110000101010100001010000000011100111010100011111010110000011011001110011010111101011010100101010101111100011001100011010001111101110101110110001010101111111000000111001011101110100;
#1 $display("%b", po);
# 1  pi=207'b110110011001010110000001101100101101100110000011100000110001111110101011010101000000111111010101010101100001011011011010000010001000101011010010000111001011000011011100001010000111101100010101101011001000000;
#1 $display("%b", po);
# 1  pi=207'b010001000111101011001111101111010101010001001001101110001010110010111000100100101111011000100010000111100011010101000101101001000010011001100100000110111101100011101110000111001001010101011011010100010001110;
#1 $display("%b", po);
# 1  pi=207'b011110100101110011001010111111110000101110111100000110111001110100110100110000100011110001011101000001001011010110001010010011101100001111100101110011011111100110101111101100110111011011000110011010011010001;
#1 $display("%b", po);
# 1  pi=207'b011101101011110010111110010000100100000010001110000011000111110111011100000110111010110001001100101111101011011001000101001010100100101011100111111000111011010100000100100000010100000001101000101010010011110;
#1 $display("%b", po);
# 1  pi=207'b001010101100011010010101101100101010010001110011010001100100110001000111101011110101110000010110111000000010101011010010101000010111100011111100101001110001110100001011111111010000110010001101000011101101111;
#1 $display("%b", po);
# 1  pi=207'b111001011100011011101111100111001111110100001111000010001001111101111110110100100010101100001000111111100101111101000010010100010000100001010010010110010000001111000001000101000011111101110011110011110101001;
#1 $display("%b", po);
# 1  pi=207'b111001001010100100110011111000000110010110110011010010111010100011011100001001001100101011010011001011111010000001100011111010000101111011010000110010101100101111001001100110111001000011110000101011111101011;
#1 $display("%b", po);
# 1  pi=207'b101001110100000100001110111100100110011101101101111111100101000101000010001011111010111010100111011001110011010000110110110110110011110111010000000101000111011110011110110100000010101011100001110100100001111;
#1 $display("%b", po);
# 1  pi=207'b001101011100011011110101100011111111011101000011001011011011110011010000011100111110110101110100110100101011011100100010110001000010001011011100010110101110100100111010111000010000011101110100010100101000000;
#1 $display("%b", po);
# 1  pi=207'b101001001011110001011001010011010001010111100111111101101001011001000001110011100010101010001111100101101001010010100100011100111001000011100110011011000111001000111111110000000100011110110111001100011000111;
#1 $display("%b", po);
# 1  pi=207'b110111011001110110111000000010000100110111100011011010110000011100100110010101100110110110110111001101110001111101000000111000101110100000101111011010000001011000100101001101010101100110001011011101010110100;
#1 $display("%b", po);
# 1  pi=207'b000011110010000110001110010011110100110100010010000000111010111100011010101011000010011001001001010011011110101111100110001110111100010110011000000110001001011110111110100101110001010010110100101101101110110;
#1 $display("%b", po);
# 1  pi=207'b010000101111000001000011110010001010001110100111100111111100011010111011101000101000110100110100110110111000000001111111101110011010100101000011010001000100100001101011110100111111011100110100011000001011100;
#1 $display("%b", po);
# 1  pi=207'b100011010010000101111100101110010111100001011001111001000100101101001000011001000101001101011001011110001010110101010001010011010101110010010011101010010011111011011100100010010011111001100001111110011010010;
#1 $display("%b", po);
# 1  pi=207'b110111101110111011101010110101110110011000110001010010110100110000010100111101111001100010011001101111010011100001010000001111011100111011100011111101010100101000110111101101001100111010010010000100111001011;
#1 $display("%b", po);
# 1  pi=207'b101100110010100110011101101011010111110101010010011001101000101110001100010100100010001111110101100011111000111101010010100100000000010110001001101011001000000011111000010011100101100010100100111000101111010;
#1 $display("%b", po);
# 1  pi=207'b110011000010110011010010001110110000000111110100101011010110010001010101010001011111000101100011101110000011000001101000100001001001100110101000101101101011100001010110111100010011111110001110011111101011101;
#1 $display("%b", po);
# 1  pi=207'b010100100111100101011111100011011001100101010111110111100000101001011100111100110110011001111011111001101000010010111011010000101010110001011011001010101001001001011110000010001110001001110001011101111000100;
#1 $display("%b", po);
# 1  pi=207'b111001111001110110111110010011000111100011100110011110011000010011010100100111001011100111001101001011111100000010100110001001111101010000101101001101101011100101111111101010100111110000111011110011010010101;
#1 $display("%b", po);
# 1  pi=207'b110111001100101010001000000111100010110101001000001111001100101101100001000110101000010111110100001110101011110111100011010010001101001100110110101101011011011001000100100101100101010100110100111010111000111;
#1 $display("%b", po);
# 1  pi=207'b111111011000001010110000010011101100010111000010111111010010101111101110100010101110001011001111010011101010011010000000101001101001110100101010010100101100100100110001001011010010010100010000010001110001101;
#1 $display("%b", po);
# 1  pi=207'b000011100011100001000110100101111100001111111100011101011011001100100011010100111011101110111001111111000110001100111100011100101000001001101001001101001011101010010110001111110010001111001100101101111010001;
#1 $display("%b", po);
# 1  pi=207'b111100110000001101000011111001011101000000100110110000011000011011100100110001000000011100111011101101001101011110110000000000100111001000100100111001010110111111100101000111101100101101000100000010010011010;
#1 $display("%b", po);
# 1  pi=207'b100000100010000010000011001101110011101000111011000101100001011110101011001101001111000101010100100100001011000001000101110101001011001101011010010110111000100111000111001110111011101101000000101101001011111;
#1 $display("%b", po);
# 1  pi=207'b110111110111000000001100000110110001110000011100001101110110010010011001100101111001011101011001111001011101110100101110011010101001100010101100101001100100100100100101100011000001101001101101010100010101011;
#1 $display("%b", po);
# 1  pi=207'b010001000110010000101110001100110000000111101110100111100000001110001110001001111010101110011010101001110100101110010101111001111100000001010111111110100111010000011011110010000011110001101111110101110001110;
#1 $display("%b", po);
# 1  pi=207'b110010000001100110101100111100111101011010101110110110111001100001011000111001111010011010111111010001100010100111111110101111101111001000111001100001110000010011111001010111011010000100001100100111011011110;
#1 $display("%b", po);
# 1  pi=207'b011000011110011101011100000011100110111100100011100101010011101100011111011100100010011001100000010111010000111111110101100000111010100011101010011011100010101111100010000001100111010010010101110000111010110;
#1 $display("%b", po);
# 1  pi=207'b100010111001001000000011110101000001000000111001011101110000111101000101011111100000110101000000000001100000100111101111001010111001011101101011011110100110011110100101110000101110110010001101001001101010110;
#1 $display("%b", po);
# 1  pi=207'b011011011011000110001100111011110111111000000011001011011111100011011000001101100000011100001001100000101001001011010000001011110011011110011110010100010010100110001101001001010000010010001101101100011111010;
#1 $display("%b", po);
# 1  pi=207'b000010101011110110100111011000100100000101111001011010011001110001101100001001000101011000000100101101100010010010111001110110101111101000111100010110110010110111111101101100011001110010011100101111000011000;
#1 $display("%b", po);
# 1  pi=207'b000001111010111110010100110011010110000110010101000111101111011110111100011011110111111000000011110111111000111000000111100001010111010001111101010011001100100010110010001100010001111001101011101100110000101;
#1 $display("%b", po);
# 1  pi=207'b111011011010011110111100101010100010011101111111001101000010111000100111011100110010100001110000101110011111100101110111010001111101111011010000011111010101110101110001001101001110110011000001011010110110000;
#1 $display("%b", po);
# 1  pi=207'b111111110110001100010110111000110110000100100000011111001110100100111101011000001010100111111101111100101110011001011110111011111001101000010110000101000010010010111101010111001110001010101110110101011101011;
#1 $display("%b", po);
# 1  pi=207'b101010110100111010010001110010110000101101011111111101100001111011110001001100101111100000111110101011000011111101110001101100101111010010010010010000111000010000101110110011000111010111100110111100000010010;
#1 $display("%b", po);
# 1  pi=207'b101011111101110011100100010110101000111011000010110101101100000100000010010100000111001001011101011110010111101111111000001111010100111110100100001000000011011010101011010010000011100010010111100111001011001;
#1 $display("%b", po);
# 1  pi=207'b110111011110110011001110001011001100100010101011011100001101100100000011010011010111011011110011011101110101000000101011111010110011101010010010100011101010111101000100110011110101110000010011001001001011110;
#1 $display("%b", po);
# 1  pi=207'b010010001111001010111000010000111010010000110000101111010010111011001010010001010100000010010111000011101000010110010000100011001100101110000100000101111000110011000010000101000010011100010000010010011111101;
#1 $display("%b", po);
# 1  pi=207'b110011110111000110111011011001100100111000001110011111011011000011101011111001000010111010100011000111101010110010001111100000011100101110110111100110010011010001111101001110101101011100100010111100111000100;
#1 $display("%b", po);
# 1  pi=207'b101111001010011000010110101001011101110101100001000011110010000001101000011111100101100100010001110111110000110110110001010011110001110001011001000011101011101110111111010100011101111000100010100000001001101;
#1 $display("%b", po);
# 1  pi=207'b000001110111000000011111011101101101111000111101000110000101011001110011001010001011000100000111110011100010001010101100111000010100110110001100001011000000000100001101111011111011000101001101011000111010000;
#1 $display("%b", po);
# 1  pi=207'b100111010010011011000001011110110011110000101001100011100001001110010111101110100000001000000010001111110000000011011110110101011100111100111011000111011000010101101010000010000011100011100001001101111011000;
#1 $display("%b", po);
# 1  pi=207'b010011111001100110110011001101111101110000000011000101111010101010100011000100001100110011110111011010110110100100100101000111011000011000110110100110011001101011101010000001110101110000010100100000010001011;
#1 $display("%b", po);
# 1  pi=207'b111001011000111111110011101101110111000011011011011100000100101100100101110110000001111010110001010001111101111110001001111000111010000000011111100111010111011001010000111011010010101010101010110110011100000;
#1 $display("%b", po);
# 1  pi=207'b111101000110101110100111111010001100111101001100001011110011011011111010000100100110110100011011111000011111010000100010100100001111110101000111101110110000010100100001000111000010110110101000001000001110010;
#1 $display("%b", po);
# 1  pi=207'b010101010011000110100100000000101100111111010100011101011001000100100111110001000101110001100011011101110110011011101010111111010111110000110011011101111110101101010110000100111110001001011111011010111000000;
#1 $display("%b", po);
# 1  pi=207'b111000111010111011010110100101011101010111011111101011001010110110111100110011110011011110011011010101100111001111001100010000000011011001101010110010100111000001111111011000000010001111011111000001011001000;
#1 $display("%b", po);
# 1  pi=207'b111011011010111011101100000100001111110000011101111010000110101001101011101001101110110110000010101101110010010010000111010000010000111001001100000101000011011100111100110111110010011110110000011101100111101;
#1 $display("%b", po);
# 1  pi=207'b101001010100110001100001101011100100110000001010001001100011110010000000010011010101110101100000111001111100111010000111011011010100011101101001011100010001100101110110110010011011101010110001010001100010011;
#1 $display("%b", po);
# 1  pi=207'b000100011101101011010110101101111001010000011010101010010001011010001111000001110000011000010011001100000101110011011101111100100101010010000100000110011101111000110100100101000010001011001110101100110101100;
#1 $display("%b", po);
# 1  pi=207'b000110011100101011000010011110111110100010001110001100010110110111000000101000011110100100110111111101101100111110111001100010110010000011111110110010011100110100101001010100010100010001001110010110010110000;
#1 $display("%b", po);
# 1  pi=207'b111110001110111110000101100110010111110000011110000101110111100101010000101010111111110110110000101000010100001100011100110101001100011100101010110001001111000010100011001000111001001001100100110111101010101;
#1 $display("%b", po);
# 1  pi=207'b111000011000000111110100010001101111110001011010100011010111100011111101100001100110101100000011000100001000111000010011010000111010100011010110101110001000011010011001000010100001100000110001011000001000110;
#1 $display("%b", po);
# 1  pi=207'b010111011111110000001101001011000110110111101111010111001101001100010011000100101011000101100011010010001101100111000011111100011001010101100110010000011110111111001101100101000011000100000001010100011011010;
#1 $display("%b", po);
# 1  pi=207'b111101111101010011001110111100000000011111011101100111111111010000001110001000010100111111010010100100000000000001101010110000010111101101000001100010110001010100110011111001110111011100010001000110010011001;
#1 $display("%b", po);
# 1  pi=207'b100010100111101000001111010001100110101011010101111100110111011011110101010101101001110011001011110101110110001000110001110110001011100000011110010011010100111000101110010000100110100111101011100101001101001;
#1 $display("%b", po);
# 1  pi=207'b100010011110011100100010110100110111101001011010110100001011111111100011111001010111001111011001000101111010011100101000100010101100000111011000001001011010111110001111011111000110110001101111011001111100100;
#1 $display("%b", po);
# 1  pi=207'b001010000010000100000110111001000110011010000111010101000001000000000100011111111011101111011101011100011111000111000001100000110010000110110100111110011110101110001100101000111000110010000111100101000000000;
#1 $display("%b", po);
# 1  pi=207'b100101100101100111010001010010001000011101011010000110001011010100001100110111100101001100010111110001111110001110001110111100100111001111101011000010110110011101011000010011001001110001001011100000101010001;
#1 $display("%b", po);
# 1  pi=207'b110000011110101100100111010110110000110110111011011111100011011001110001101110111101010110100010001111110000010011111101111011000001010100100011010011000110101000111001111100001111111010100110000010100000100;
#1 $display("%b", po);
# 1  pi=207'b011100011100100101101100001101001001110100100010101111001101101011100100110101110100010101010111011111100110111111111101110010110100010110110100010001100100101101001110000011101111111010010101111111100101011;
#1 $display("%b", po);
# 1  pi=207'b000010111011000001000011010011100110101100010111011101010110001110010111011001001101010001011000101011001001100101100010010000101100111010101101010011100000010101101011101110000111001110010011001110101011101;
#1 $display("%b", po);
# 1  pi=207'b101100110011111010000010011101001111111011111011111111000010010100011110000001100110010110100110110001001111011010110100100100100011110110000101011010100110100110100100100010110110100100110011011111000011001;
#1 $display("%b", po);
# 1  pi=207'b011101000111111010010101010010011010100100000110011011111011010010010111011111001000101111101100011001110110001111010101011101100101100110001101010010000100001000010110110010111010101101101010001010101101011;
#1 $display("%b", po);
# 1  pi=207'b110000110011010111110101110000001001001100011111110111100011011101101000101100010111110010110010100011110011010000100110000010111000001111010110111001110101110001011001011101000111111100001110101000011011000;
#1 $display("%b", po);
# 1  pi=207'b111010111110010111011111110010100101111110000101110011000011000110010101101101101100011000111100010110111001011111101010100001110011011010101100111111101010110010010001101010111111111001111101101101011110100;
#1 $display("%b", po);
# 1  pi=207'b101001001011001000101110010101110011110010100011000001001100101111001111000101000010010000001000110111001100100001110010110100111111111100000101001100001101111101001011101111001001010001010010110011000010111;
#1 $display("%b", po);
# 1  pi=207'b000001110011010010010010101111101100000001101110001011111010100000010111001100110110101110111001010100010111110000110111100110100100101000110101100101111010011010100100110001001111111101000100001110100101000;
#1 $display("%b", po);
# 1  pi=207'b001100101000011111001001011000101111110100111101001000100101010100101001010111001100010011101111001011011000101101000110110100111101100111011001111000101100011110010000000001101010100110100011011100110111000;
#1 $display("%b", po);
# 1  pi=207'b110101011100101100110010101000111100101101011101100111110111000010001000011100010001000001110000100000110111101100101100100101010111110111000000011000011111110011101011111000101111101011111100000000100110010;
#1 $display("%b", po);
# 1  pi=207'b110000000100000110110110110011110100001001001100010000000111001001111110100100111101011110001000011010001000000110011100110111111000010101011001011011101110000110101101000111100100010110100101101100100011000;
#1 $display("%b", po);
# 1  pi=207'b110100011100000001001000010110000011100011010001100000110110010000010101100011000011011010100100010111101111000011000011001010011010101100111001110011000001101001111110111111100100010111001010010101000110111;
#1 $display("%b", po);
# 1  pi=207'b010010011110111000100110110010110110100010011110011101001111011001101111000100000110100010000010010010001110101100111000011111000011111011011001111000010001010001111101100000111011110110011011010001101000110;
#1 $display("%b", po);
# 1  pi=207'b110011011010001000110110011001000110111001100000000101010110111101100110011001001100011100011000100000101000011010110110101100111000110100001110101101000010100011100101101100000010100010110110100011101110101;
#1 $display("%b", po);
# 1  pi=207'b000111001000011110101110110110001010101011010111001111010110011000100110001101100100100111000000011101000000110110111101111010110000100010101010100110111010011010101000111011001010010000010110000100000010101;
#1 $display("%b", po);
# 1  pi=207'b000000011101010000100001010111101001101000101010111001011111000101110000110011010011100100000111101111110110110010110100100111100001111001111110001000010110011110110010001011001110010010100101011101010001010;
#1 $display("%b", po);
# 1  pi=207'b100100101111000101000110100011000110001100110000000000010011000101100001101011000111010010101101000101111010110000001010010111101011011101110100101110110100110011101001010011100011001010100110100111111111000;
#1 $display("%b", po);
# 1  pi=207'b011100110001011101001111010010000001110111001010101101010111111001001000010000110010001101000010001111001011011111100001000101010011011000111001101111011010000100011001101111011101011111011001101111001101100;
#1 $display("%b", po);
# 1  pi=207'b001000111011111111111000010001010010111000110011101011000111001110101111111011101111101100000001011101010111111100010000000011100100011111001100001011001110010010000110111101001001000110111010000000100011100;
#1 $display("%b", po);
# 1  pi=207'b101000011011000010110111111010011000110100000100000010111001101101101001010101101110001101010010001100111100011001011110011101000011110000111111110100111011000101101110100110001100100101110000111111001110001;
#1 $display("%b", po);
# 1  pi=207'b101011001101000011110110111001100111011011101000101101101000010110011111101011110110101111111000101000001011010101100111010010000000101110001000001001101000010101011100000100001011000001000111010110000000110;
#1 $display("%b", po);
# 1  pi=207'b101111100011111011101001101001001010001111110000011100101111000100001111000100000100101000100110000000110010001000010010010100010110101100110110101100010101000100100101011101001101111101101000011000111010100;
#1 $display("%b", po);
# 1  pi=207'b101100110011111011111000001000001110110011100011001111000111001010111001000110010111011100101000100111100000101100010001010101001110000110110110011101101111010100111110101010000101010110000100011100011000001;
#1 $display("%b", po);
# 1  pi=207'b111111101011000001001011000100100001011100011001000100110100000000001001110110110111010001101110110000111011000010001001001000010101001011111111101010101000010100100111101111000111010111110001001101100010001;
#1 $display("%b", po);
# 1  pi=207'b011011000011011111101100110010010101010000011011011100011101001011100100110111111010111010010101010110000010101100101010111110111101100110110111000001101011101001001000000101110000010010001001001111110101011;
#1 $display("%b", po);
# 1  pi=207'b011111001011000011101011000000010110000001101101010101110101111010001000011111100101000110111000100100110111101000011001001001100011010010100010111101000101100001111001010100100110011000011100010001001001010;
#1 $display("%b", po);
# 1  pi=207'b101010000010101001101100000011000101110010110011100111000100010011011110000111111101001110100110001010110110110011110000100110000110000010010110110010000001010001001001101100010111000111011100000111001101001;
#1 $display("%b", po);
# 1  pi=207'b000101001100011101010001100001111110101011110011000100110011010100110001100001100111111101101101000011111100111000010010001010110000101101101100111101100101011101001000111000110010101110101000001111100110010;
#1 $display("%b", po);
# 1  pi=207'b101001111010101101100100011100010010100000101000111010100101001101110010000001101100000101010001010000101100010101010110111011010001001001100000000100111001011100111110100001010001000000000010011111111110111;
#1 $display("%b", po);
# 1  pi=207'b101111110011010101011100111000010101000111010001011111111101101000101000010100000001000010011110111000100010000100111010111100000000001101101100101111100111001011110111111000110111001000001010001100001000011;
#1 $display("%b", po);
# 1  pi=207'b000000110010011001100100001011000010011000010010000000001010111110011110101010110010101100111011101000101001011110110111000000000001000011000001100001011010011101011011010000101010111001001100000010110100100;
#1 $display("%b", po);
# 1  pi=207'b000000111011100000111010011101101001011110011101110100111110010101010101101100010011001110001110010111000011000111111111001110111100011001011011100011001000000100101001001011001010010110111001100110011011111;
#1 $display("%b", po);
# 1  pi=207'b001110110001010111110110101100010010011001000001111000000000001001001111101101111001010000110110011010001000010101101110001011100011000011111001001000111001011100110010010010001010000011000011011100111001101;
#1 $display("%b", po);
# 1  pi=207'b111101001100000100000010100110111111101100001101001100100010001100100001011100110000110111101111110101010110101111101011100001010000001111010000000010001110101010000101000010111110101101101001011110110100011;
#1 $display("%b", po);
# 1  pi=207'b001000011101000101110110010001000010000100010100010011001001000011101000111101101101101111110111110101011010011001110010100101010010100001000010010011100000111011011001000000001111000011011000010101110011001;
#1 $display("%b", po);
# 1  pi=207'b011100100000000001101101111110000101111111110010101000001101101011011010000101011111011111100101001101010000100111110001001011101100001011101110100000110011011011010111111001100000101100100101001001000110110;
#1 $display("%b", po);
# 1  pi=207'b010000111001001000101010110010101100101101111000101001110000011000010101000001010000100010101011110110111111111111000110001010101110000110000011111010111100010101110011000100100010001111111101010011111111111;
#1 $display("%b", po);
# 1  pi=207'b111010000010000111000001010000000110001110101111000111000110001100100100001010111001000010011101111010010000111001011111101000000001111100000110110111010000110000110000001000110011111101110111001111111110110;
#1 $display("%b", po);
# 1  pi=207'b101101000011001010100001010000001110111101001001101110001000001111000001011100010111000111011101001100111101010000110010000001011000110101100011101001110100100110101010011000100100110001001011101010001111110;
#1 $display("%b", po);
# 1  pi=207'b101110011011001011110101110100100111111010111101110011001100100101101000111100101110100111100010000111011011010010011000111010001100101010110001011010000001000001001111110001000010110010110110011011101011010;
#1 $display("%b", po);
# 1  pi=207'b000100111101101101100110010011100100111110011000000010000111001111000110001000101101101000101110100110011101000111011000011110011100110110110010001001101110111000000111000011110110101111000001100000011010011;
#1 $display("%b", po);
# 1  pi=207'b011010000010111111001101111101110101001010010111100101100111010101000001101010110111111000011101111111100000000001010001100100110000010111010111101100110101000010011100101101100010111001011100100100010011111;
#1 $display("%b", po);
# 1  pi=207'b011101101010000001110001111010100101001000101110101001001001111111110011000100010010010011101100010011010111011001100010110001011100000010010000011110011010010010100011011011100100101011111111011100100101110;
#1 $display("%b", po);
# 1  pi=207'b000100110111010010111101001100111110110110001101011110000000011010100111111110001011000001010010111011111010110111100011011010001010111001011001111110110110010001001010011111100000101100101010110010011001101;
#1 $display("%b", po);
# 1  pi=207'b001000110101101000001111111010000000000010010111110111010011100000111111010110101011000010000110100110001100001001101101101000111001110010101010111111000101000010101110001011110000110011000101010001011010101;
#1 $display("%b", po);
# 1  pi=207'b011111010110011010101101101000001011001111010000111010101010010000011100110101111001100101110110010101111100001110010000000100100000100000010001001010001110001101010010000110110000110101110100111110011010010;
#1 $display("%b", po);
# 1  pi=207'b000100110001101000000101100001000001111010110110001000010000001000001100010010101001010001111000110011000001111001101101101011011100010011011011101111110000010010100110000111111011010011111110111000000001000;
#1 $display("%b", po);
# 1  pi=207'b000000010111111001111110011001101100110011111101111100111110011000000011000000000111111010110010000111110000000100011001001111001010001110110101000101111000100111011111100010010010110101111000000111010100111;
#1 $display("%b", po);
# 1  pi=207'b011111011000100111011011110000111101001001001100000011101011101010000111110001100101000111000110011111001010011100011010001101010101010100101110110010001010000000000000000101111111010001101110000101111110000;
#1 $display("%b", po);
# 1  pi=207'b011011111011110111010000101011100011110000010111001110001011100011100011011011000101100100100001010111011111001001010100100111110101001101001000010000100110100101000111110001010000010010011010001000101101111;
#1 $display("%b", po);
# 1  pi=207'b011010011101001010000101111110001001001011101100010101101011110001000101101001110101101010010111011100010001110111101100011100101000001110001010000011011111100001011010111110101110011100111100000010011100011;
#1 $display("%b", po);
# 1  pi=207'b011111000110001110000000101101111000100110000100001011001010110110110001000101111111100100011010100000011001000000011000111100000000110110011111011001001101100000010011010000101001110100010011010010010101001;
#1 $display("%b", po);
# 1  pi=207'b001100110011110101010010011000010110100100111111000111010001110110011011011110111010100010001110101001101100001010111011111011011110011001100111010111000100100000011011000011101110101010010001011000000000010;
#1 $display("%b", po);
# 1  pi=207'b111001111011110000111010111000101110111011000110101100101000101100101010011000000101101111000100011010000110110110100010010001000100101100000000111111100010110011111100111000000111010101100011001001100010100;
#1 $display("%b", po);
# 1  pi=207'b010001110000001001000101101111111101110110000010010011000000001110100101101011111110100010000011110110011100011101100001100110010100101000111010100000110100001110110010011001101011100011100001011111101001100;
#1 $display("%b", po);
# 1  pi=207'b100101110101010011111000011000111101110111110101110010101000010010001110001110100100000110010100000111111001111010100101111000010101111100110110101001101101110010011101001111100110001001100011111000100100001;
#1 $display("%b", po);
# 1  pi=207'b100001001000001110000101010010101010010111011111011100111101110011101100000010000000100110011111110000001110000110101000100011100011010010101001010111010001001110110011111101111101010101111011001000011111011;
#1 $display("%b", po);
# 1  pi=207'b000111011011011111101010011100110011100110110011011001110111100011011011001100010000111100100101111001011001101001000000010101010001101100010110011010100000001010100111011010000011110001001001000000111010000;
#1 $display("%b", po);
# 1  pi=207'b000110000011000100010100001111101011010110110000010000001001000010001000011111110010000000101010000110100011010001010001100100010101010001101010000111000101111001001110111001000100101101100010100011010110001;
#1 $display("%b", po);
# 1  pi=207'b100100111010000111000000100111000000001110011001010111011111101100110101101010000100001001010010110101011100100010100110111110011100000001101010111111111001101110111001010111011101010011011101110100001011110;
#1 $display("%b", po);
# 1  pi=207'b110000001011110100101011001011001100100011000000101101111011101111111011010010001000111001011010101111111100010110111011100100011111010011011010010011101010100100101111011110011011100111011100010001101111110;
#1 $display("%b", po);
# 1  pi=207'b101100110010101111000110011111001000101110011001111000100000011100101001010111101111011110101000011011111100011111011000001111001111010010011011010110101100010111001101001010101100111111100110010111001100001;
#1 $display("%b", po);
# 1  pi=207'b111101101000011010110000100111001011010000111011011110011001000101000101000100100100111001110010011001110000110110100010000010000111111101101001100001100100111010011110101001101000011100011010100010001001111;
#1 $display("%b", po);
# 1  pi=207'b001010010000010000011010010110101011000001100001010000011000100010110011011110010010001111110000111101001100000010100110000001111110010001010000111001111100010011011001100111110100000011001101011000010000100;
#1 $display("%b", po);
# 1  pi=207'b101101010100100011111110110011110000111010011100101001101101111111111101010011010011000100111110000101001100010000001100110110101010000101011011000001101110110101000101000100100000011111101011010000010001111;
#1 $display("%b", po);
# 1  pi=207'b101000100010111101011011111010100010111001101010000001100011100111010100101100010010101011001111100011011010010011100001001101101001111011010111111001100000100000010111101000100100110100111100111101011111111;
#1 $display("%b", po);
# 1  pi=207'b011000101111110110100001000011000001111011110100100011000011010001100100011110000111000001001101000011111000101001001111111011101011111010110000111000010100100111010011001010000010001100011100010100010001001;
#1 $display("%b", po);
# 1  pi=207'b110000100111001001111100100101100010110000101011100100001001100001100001001101101010101001001110010101010000111100011101000010111101111000000000101100110101100100000000000101101001011011000101011011100001000;
#1 $display("%b", po);
# 1  pi=207'b111100100101100000101101101011111100100010001100111100111100111100010111111011001010100010000101100010110010010000100100001000011011000111011001000011001011101110111000100101111011011000100111101111010010111;
#1 $display("%b", po);
# 1  pi=207'b000011011111011100011010011110111110000101011011101110101000101010100001011100101010000010111001111110000001111110011100000000010100010001001011100101111101111110110111111000010001111101000001011010111100111;
#1 $display("%b", po);
# 1  pi=207'b111011000010001110001001010111101100001110100110010110101100011011110101010110110000010110110010111011001000100010010010010000101100001100101100000111111110110100110001001010011000110001111001110001010000111;
#1 $display("%b", po);
# 1  pi=207'b001111100000111001011000010011100110111111110001101100011111011001010111011101010000000101110111101111010101011001110010000001001111101101111100100011000010111111110011000001011111110010011101110100000011001;
#1 $display("%b", po);
# 1  pi=207'b100011000110101000100001101111110111100010111010110101000011100010100110101011110001100100011000000011111011101110100101111111111110100110100011110101001100010110110011111100010110110010100100011001000010011;
#1 $display("%b", po);
# 1  pi=207'b001001111101100011100010001010011001010010111110100110100000101010110010011110110110110011101111110011100111101101101000001011001101111101010100000011001101011101011011010001011110100111001100000110110100111;
#1 $display("%b", po);
# 1  pi=207'b110100000111101000101100001100010110110111011000111001001001111010110010101111011000100011101010000011110001001111100011110100011011110101000100000001011001000101011111101101011000001001110100101110010110110;
#1 $display("%b", po);
# 1  pi=207'b101000111000001100011010111000000001001111101010011011101000010000100011000010110010100110111100110011101001110010111000110001011111100010101111110100101100010011101111001110101001010010101001110001000110101;
#1 $display("%b", po);
# 1  pi=207'b110110110001011100000011011100100010011100000111101111000010110010101111010101001001000001100001110110010100001000010011111010010001000111000110010110011110110100001010110110110111110111100000001001110110001;
#1 $display("%b", po);
# 1  pi=207'b000001100100100110010101010010011000101100111010101010010010011111000011001100010001111111111001101011000101110110000010001100010011011100101001100010001000100000100100110100100110111001011110001111010101001;
#1 $display("%b", po);
# 1  pi=207'b100100011001000000000001010101011010011000110111010000111000110111110000000000011111111010000100010110010001111100001000100110110000101100001011101110000111011001010101000010011001010111100101110110010110010;
#1 $display("%b", po);
# 1  pi=207'b001001010010111100011010000110001101111000000001100111111101010010101010000001111101110111100111010000011001110110111111110100001110011110100010010110011101010111110111100101001100101110100101101001111101010;
#1 $display("%b", po);
# 1  pi=207'b011011101001010000101110100001011110000100001010101010000100011001111010010101101001010000111010111110100101011010111100011101110110111000010001000100011101111101110101101000001100000000111000000001111101101;
#1 $display("%b", po);
# 1  pi=207'b110011100001010101110000001011111001100000101100011000001010011111100000010110000000100000010010111010010010000001010010010000011100111111000011110001110110110100110111100000101110111111011000111000011011111;
#1 $display("%b", po);
# 1  pi=207'b100001000101101111010000001001001011100010110100001000001000110110010111010001010000110000010101011111001100011011011010011011010101101011011010000001101110101111111101111110100000011110110000111000101100000;
#1 $display("%b", po);
# 1  pi=207'b100111101010000000111100101010011011111011001100001000111101101010010110000110101110010011000000000001111111111110100000101000110011000111011100001110111111010010001111010101010011101111011110001001010010110;
#1 $display("%b", po);
# 1  pi=207'b000101110110001000100100001101110011110101000101111010011110000010100100001000100001010010100100100000100001001010011100010100000100100111101010011100100011000010111101010000001101111000000110000000011011010;
#1 $display("%b", po);
# 1  pi=207'b100001101100000001000011111111101101101101011010001101000010010100110110011100100100000111000011110010000100001000101001000111100010001011001101001111001100111101110110100101000010010011110011011110100010011;
#1 $display("%b", po);
# 1  pi=207'b001110101001001000011001111000111111110011100000010000100100110000000010000011001010101011101010110100110101001001010101111001011100101010011101010010111100010101011011100100111111001001101011000011111100101;
#1 $display("%b", po);
# 1  pi=207'b010011001111001100111011000101010100111111011100010101101010101011111010001011001111111110011111011111100000001011000100100100000110001100100101100111001110011000110110001100100000110001010111110010000110110;
#1 $display("%b", po);
# 1  pi=207'b101101110100100010100101110011100010110010001101101100101101001011001001011001010100110110001010011011101111000110010100100101100001000001000111011010101000101011101101110000100110001110100011000101000010001;
#1 $display("%b", po);
# 1  pi=207'b111011110111001101001110110011001100111010000101111111001111010010110011111001101011111010001111011010010000101011101010110011000100000011101001110101000111100000100010000110100111111110010101100011010101000;
#1 $display("%b", po);
# 1  pi=207'b011011101110100101011111111000011101010001100101110101111111100100011111110011111101111001010000110010000101100000001100100101010000110000110001101101001100101101010011101001111000101001011110011011011100000;
#1 $display("%b", po);
# 1  pi=207'b000001110001100100111001000010001101110000111111001001101000101101001100110111011010011001101111001110111101100010010110110100001011011101101010000001110010011101010101110011101100000111010010010111011100111;
#1 $display("%b", po);
# 1  pi=207'b101100011000010110101010111000011011101001111011110111110001000000111110000100100010001001100110110101010011011000100111101101101011001011110100111001100100111011111100000111100101011100100110110111111110101;
#1 $display("%b", po);
# 1  pi=207'b100011001111100101111010101001000010011010011100110010100100001111001100101001010011111010101101101001100000011111010111011101111101100100011100010110111101101000100011010111000100100010011110010010101000000;
#1 $display("%b", po);
# 1  pi=207'b100110110001101110100011111101011100001001100111000111000111101111011000001001111000110011010110111100011001100010101011001100010110000010001001110000011011100000100100011010011011001010001111010001101011001;
#1 $display("%b", po);
# 1  pi=207'b010100010010111100000111101010100001000000100000101100010100000100111011010010010001111110010101111100101010111101101111101110000011001111000001001000010011001001100110000011101001111100101100010001011001100;
#1 $display("%b", po);
# 1  pi=207'b001001111001001100110000000101010011010110001010001101001010110001100111010101001101010011010001101011100001101001111001001100111001111001101001101100111101010011001000100101101011011100110010000011111000101;
#1 $display("%b", po);
# 1  pi=207'b100000010100110100111000000011001101100001011010001001101111110100011100010000110000110100001111111101001010100000111000000001110101011010110110100011100110111100100100111110010100111111001110001011000000110;
#1 $display("%b", po);
# 1  pi=207'b110101000111011000011111100001011111010111111101101100001000011010000000110001001011000011011111111111110011100101001011101011101100001001110001100001101000100000001100010000100111010001001011000010100100100;
#1 $display("%b", po);
# 1  pi=207'b011000001001000100111100000000010001011111010111001100110111010111110110010010101110001101111100010111100010011111011111010111000010101101101100110010101111000000111000101100110010001010000011001011101100110;
#1 $display("%b", po);
# 1  pi=207'b010011101010111110011010001001100111110100001000100100010101110111110111000000001011111000010010011101000101110010111001111001011001111101010000010110101100001100110011000001101010001110000101110010110010100;
#1 $display("%b", po);
# 1  pi=207'b000100110011010010001110010110000001001010100001111001101010110110000101010110100111110001101011001100011000101101111111010010111010010000010110100100011111011100001011011100011010000110001001100101011001000;
#1 $display("%b", po);
# 1  pi=207'b000110000011000111000111111010011111110001101010100111100101000101101001011100010011010101111000001111110101000011000111010001011000011110111110000110101000101101101010010010011011111101010001100001001010111;
#1 $display("%b", po);
# 1  pi=207'b000100001111010010111000001111101010100100101110010110111110101000101000010000001100110101101010000101000110110111011110110000001010011101000100111111011111010100110111100000111100110001101010110010001001000;
#1 $display("%b", po);
# 1  pi=207'b010110100001111001101101010011110111001011000000101111110110011010010010011110111010111110101010011001110101100110011000001100010101111001111111111010000010010101010100100010101000000100100001001101001110110;
#1 $display("%b", po);
# 1  pi=207'b001100010100010000111111010101011100110000100011010010001000000011110001001000011100101010000011010100010110100110011000100110010110001000011111000100010000111010111110001111111011001010101101001011110100001;
#1 $display("%b", po);
# 1  pi=207'b110001110111011001100001100101110101111000111101000101010011101000010000000111110010110110010100111011000110000111001111001101101110101001001000100100000100001010010001101011000000000101000110111001011011100;
#1 $display("%b", po);
# 1  pi=207'b000011001011000101011001101000010000110001011110000001011000001000001011110110010111010111101011010001000110011100011000110000010110111011110100101000010000111000100011110101001110100001011110010011100011001;
#1 $display("%b", po);
# 1  pi=207'b101000111101101101010101000001110011000111111111001001101011101101101001010011001001100111001110011000101110001000111110110000101101011011101000000001101010001111011110000110101000110111110100110101011111011;
#1 $display("%b", po);
# 1  pi=207'b001000000101110010000001101000110111100000100001101100111111001101100101101001101100000000000110010000100111001110010110001010110000111000000101110100111011100001011010110110101010000101011100111100110101100;
#1 $display("%b", po);
# 1  pi=207'b011111000110111110000010111011100101100110001001010110100110010110101101111111110010011011111010010111100101010010111100111101111101000001100110110010010101001111111010011111111100011010110100010101111100001;
#1 $display("%b", po);
# 1  pi=207'b010000100011000101011111011010111110111000110110110010001010010100001100100100000000010000000000010110000111100110101100110000001001101011101111000101101101000001101101111000010000010101101011110010100001111;
#1 $display("%b", po);
# 1  pi=207'b000111010100011011111101101110111011100011100111110101100011111110001001001011011011011011000000000001010111111110110111010000000101101011100010010010111101111110001000011101100100001110001000111111110000100;
#1 $display("%b", po);
# 1  pi=207'b111100100111010111100111000111000111001001010101001001011101000011101011101110101000011100000101111010011010010011111001001001101111110100000111111111101110101100111100101011111101111100010111110111000011010;
#1 $display("%b", po);
# 1  pi=207'b101011101111101111100001001110100010011111111011011110011000011010111001010111001001100010001111100011111000010000011101000000111110011000110110110110010001000011101000001011110100101111100001000011111101010;
#1 $display("%b", po);
# 1  pi=207'b011111011001000101001001110001000101110001001110010011001010011101101111100101110101101100000101011000100100000000010111110100110001111001000100001000110011111010010100110001100100101000110101000001011110100;
#1 $display("%b", po);
# 1  pi=207'b010100111101100110110111000010011001000000000110011000100110000000100111100010111010100100110100111110000000010001000100111011011111100011101011000011001011011001100100010110110111001111100000101111110100000;
#1 $display("%b", po);
# 1  pi=207'b100010111111100111000001101010100001111100010011110001110101111011010111111100110110100010101001100111101000011111101100111101100000111001111101110001111011001110000110011001011101101001101010010010001001000;
#1 $display("%b", po);
# 1  pi=207'b011111000001001111100010101101010000010011110010001100011110100110100001011010101100011111100011110000000111101010001110000111000010110001111000100000001000101010001000010001111110001010001100101100010101011;
#1 $display("%b", po);
# 1  pi=207'b010000011010011110110101110010011000010011010101010100110000110101000111111011111111100100101000100100100010001000001110101101001000111111000101001101000100110101100110101100010011110110010101101101110001110;
#1 $display("%b", po);
# 1  pi=207'b110111100100110011101100011101000000011100101010111000010100000000000100100110011101010000010110100011100101010100011001111100000001010010001001111010111010111000001100110001110101011001100011111100001010000;
#1 $display("%b", po);
# 1  pi=207'b000001010101000000000000101000001100100110100010110110010100000010001011101110101101101111100101110111000111000010100100001011000100111000001001010010110011101101000010111101000100110001011001100001001011110;
#1 $display("%b", po);
# 1  pi=207'b100111010011010100110110110110001101100010100000001010111001010111100000001110101110101111100001011011100101011100000101101001001010111001010100011100100000010011110100101010000010001110101001101100111000000;
#1 $display("%b", po);
# 1  pi=207'b011110001000110111010010110010110010100111001011101110101101101000100000000111011111011111110101100010100010100100011000110011000100100101101100010100110001101000111000100000001011011100101011101101000001000;
#1 $display("%b", po);
# 1  pi=207'b111110101100100001101100000000100001000010101000111001010000000010010010010000100010001001100101001110001011111100000111100110011100110110100110001001101010111111011111011011111101111010000110111010011101101;
#1 $display("%b", po);
# 1  pi=207'b111100101010100000000100011111100110011101110001110010111110101011111011011111101001010100100000100101100110101111110001100001100100011011110010111000110011010011010010110101100110001101001001010101001000010;
#1 $display("%b", po);
# 1  pi=207'b100001000100011111111111111000100111000100111010000111100101001100011001100011100011000100010110110010110111010111010111000111111000110010111100010000000111000100011111110011010011000000110011111010110000001;
#1 $display("%b", po);
# 1  pi=207'b110111100000000010101000000001010110110110111101100110010101010000101010011011100100110101000011111110111000111000100000100011110111101101111110001110011001000000111101110101111000010011110110000000111111110;
#1 $display("%b", po);
# 1  pi=207'b110011111000010010001011001010001000101111101000010011011111011000110100000011110111011001001110100000100000001011111011110101100001001000010011110011010001110111011110101010110001001111010101001100011011010;
#1 $display("%b", po);
# 1  pi=207'b001101101000111000001101110100011001110001011010011111110101101110000010100011101000000010000111000100011110110110001010010100001000111111100110001111011110001100110001000011010101001001101100000010000111011;
#1 $display("%b", po);
# 1  pi=207'b100001001011110111111001000101011101100101000001100100111101000010010001100010011000000011011110011100000100111101001100011010101010111001100101001000100100101010111111010110011111011010010110010000010001011;
#1 $display("%b", po);
# 1  pi=207'b000110011011000011001101011101111111000000011010101011010000111111101110101100110100110110001011010001111000101111001000101000111111011100001100110111111010100000101101100001010100110100110000111010010010001;
#1 $display("%b", po);
# 1  pi=207'b110010110100001110011111100100001101100100010000111101111010001110101011111100111011101010101111100010111100011101011111010100010001101010110001101001011011001101000100101110011100111001001010001110101010110;
#1 $display("%b", po);
# 1  pi=207'b101110101100010010000000100010101001111011110110000000111001100100011010010111001011011011010001101001010100000100001100010101010011110000001110110010101111111110111110110010111000011011010001000000100111110;
#1 $display("%b", po);
# 1  pi=207'b010101111001101010101010101101101010100011110001101011010000101010011101011100110000001101110000001001011110111010010011101001010011110011001101101100010001000001110111010010100001011010110100111101100011111;
#1 $display("%b", po);
# 1  pi=207'b000000100101001010011001010100111111110000100001000111111010010011001001101011000011100010010111111011001110111110110011100111101100001000101111010100011010111001101001011101101000110100001110011101000100100;
#1 $display("%b", po);
# 1  pi=207'b111111101010110001000110100000100101101000010101000100111001110010100001010100110101011011000101110111000100000101000101110000011000100101010100100100100110001101100011101110100101110010011110010011100100011;
#1 $display("%b", po);
# 1  pi=207'b101100010111111110111001001000111101110101100111110111011010001110011100110101110011001011110011010111011100010000111101101101111000100110010011101111010110011100100110010011000010111010000101001111101110100;
#1 $display("%b", po);
# 1  pi=207'b001111101100000011101011001010001001000111000100100111010101001100001110001011000111110010110001111111101100011111011011001000000101011111010010001011011011000110110101001001101011000111101111100000101101111;
#1 $display("%b", po);
# 1  pi=207'b101001111001110010110010110000110001011101001111111010100110011101101001001111001011000101010010111001011100001111101110010011101101001010011100011000011010010000010101111001111111011010101110010101101001010;
#1 $display("%b", po);
# 1  pi=207'b010011000100100010101010011100010111000110111001111110000110000100110011010000110110100111101011011100101111010011000100000110011010001111011110011011110011100010010111011010000001011100100000001000110001000;
#1 $display("%b", po);
# 1  pi=207'b000011010101011101001010110011000100000001110110110001110110110111100111011100010100000010110100101111010000100000000101011001101011010000110000110101011010011111011100011100111001111010100101011111100111111;
#1 $display("%b", po);
# 1  pi=207'b100100000010010001101111110101000000011000000011101010100000100010101011100000000111111011101010000000111001001010111101100101011110000110010011110100011011010011011100101010101110001111110101111111010011110;
#1 $display("%b", po);
# 1  pi=207'b011001011101100001010101101001110101111100110010100001010010110000001110110100111111101111010110101110101000110001100110111110100101010010010000101011001111010110000010011101011000110011101011010000000010101;
#1 $display("%b", po);
# 1  pi=207'b000011001010000010110101000101101101011101000101101011101010000110100101011101000101011001100101011001111101101101100011101101010010111111000101100111011000010101000101000001000011111000000011011010101001100;
#1 $display("%b", po);
# 1  pi=207'b000011001000100011110001100110101100101101110010011000101101111110001111111100010000001111000100011000000110010010011000111001011110100010110000011010010111001100001111011001000101111000000001100011101000000;
#1 $display("%b", po);
# 1  pi=207'b010110010101110010101101001011000001001111000011111111010011101100110101111000011100010011110100000000000110111000000111100101000110110010001001010111110101010010000101111001010010101000101000000101111011100;
#1 $display("%b", po);
# 1  pi=207'b100000000001100101111100000110000111110110010011001100101010001010111101010111110010111000010101100101101000010111010101101000111101001110011100101110110100000010001100110001001000011000001010010010101000101;
#1 $display("%b", po);
# 1  pi=207'b110101110100111011011011111101110100010101000000001101110001101000100110110011000111001110001010001101001101110110100100000011010101000000000000010101000000100111110000011110001011111001011101000011101001100;
#1 $display("%b", po);
# 1  pi=207'b011011111010100000110101110111011001110110110101010110011010110001011011011110101011101000011100010000000101011000110011000001101001111001110110111001100010110001000000111110111011011100111110101110010101110;
#1 $display("%b", po);
# 1  pi=207'b010010110111001100100011100110001101100101111001110110011110110101001100101101101101110100000011010010101011111111111010001011100110011011001110001110110011110110101010011101000000111011101000000111000101011;
#1 $display("%b", po);
# 1  pi=207'b110111100000010010111001101010110001111110010101100001011100001010010010101100101111111001001000101001111001010000001000110011110110010010010010100001010010111100011000100001101000110000000100111101110111011;
#1 $display("%b", po);
# 1  pi=207'b001100111010011101100011110111010011111111101111111100111100111110001011000110010000011110101111001011001000011100001001011010110111001001111010101010000110101001000010101010111111010110110110100101010110110;
#1 $display("%b", po);
# 1  pi=207'b001000101100010000110111110011111010011000001110101100101110101011010010010000101011001111010110101100101010110101110101000100011110100011000000001101001001000111010100100100000000100111001111111111000000000;
#1 $display("%b", po);
# 1  pi=207'b100101101011100100001011001101111001001011010010111000110101011000001100000110101110110000101010110111111011111010110110000011000100010000101111010000001100000101111101000111001100100110011100111010111110000;
#1 $display("%b", po);
# 1  pi=207'b001111101001110001000010101001110010110101101101010001011011111011111001010001010010101100000101000011000100011100010101001001111100111111100101000011101111000110111110011010010001111111000110000110010101100;
#1 $display("%b", po);
# 1  pi=207'b000110111111010010010101011111100001010111011111101011001100001000110110011001010010101111101011011001011101111110000000000000001101110011101111001010010110101100000111011101100001011010100111101101110101110;
#1 $display("%b", po);
# 1  pi=207'b000001100111100000001100001010000001111011010001100100000111100101010001000111101000011011110111000010111101100111011101101000101010011110001111110110110011100101100101100110100111100110010011011011011001100;
#1 $display("%b", po);
# 1  pi=207'b110001010010101111110110010011111001011011110011010010001110101010111001101011001111001100101111100101110010000111011100111110110111110110001001011101101000101110101011000010010000000001011000101110110011010;
#1 $display("%b", po);
# 1  pi=207'b000000001100010101001110001110011100010110110101100010000110001111101101011000101001110110101011100011001100110000110001101001100010100011111101101101110001001110001111101000001100110010001100100101101111111;
#1 $display("%b", po);
# 1  pi=207'b110001000011000001010011010111011011001101010011111100111011101000010010011000110001000000110101000000000110100110000000110000101111011101001000101110000101101111101011011100110110101010100110001001001010110;
#1 $display("%b", po);
# 1  pi=207'b110100110110011100100111101101011011001000000001110001100011101101100000001000101111101000010100110110100000110100010111110001101100110011001010011101000011011100101100101110001110100101111011100100100010010;
#1 $display("%b", po);
# 1  pi=207'b010110100110110111001101101100101010101101110100010000101110111001011010001101000111101111000001111101100011001110101111011110000001101111001010101010010101111000101100010001110100011111100100100000011010010;
#1 $display("%b", po);
# 1  pi=207'b010011111010100110001011000101101000111101101110001010101001010101000001000001001100001001010110011111100101011011100100100001100000001000101000100101001000100100000011010101101101100001000010111101010110111;
#1 $display("%b", po);
# 1  pi=207'b101011100001001010000000010100100000110101011100110111111001100001111001101111100010010111001010010111101111100010011010101010100101100000100100101110100110010011010110000111110100001111000110001110001101100;
#1 $display("%b", po);
# 1  pi=207'b101100100111101110111101010010101011000101010001111100010100011010101101010011101110000010010111001001100110101110100000111011000010100110001111010110000000100111100111010110100001111010100011101000110000000;
#1 $display("%b", po);
# 1  pi=207'b001100111101101100110101110111110111101001011100101101000101011000111000010110110100001110100001100111001100101110100110011011010101000110100110000001010001101110100111111100100101011101011000111001110011010;
#1 $display("%b", po);
# 1  pi=207'b100101110001001111010110110100100000000101001101100110111100011010110100000111110000010110101011101100011001010010001001110010111000101001010111010110001101100101100101100011001111011000110101001010011001010;
#1 $display("%b", po);
# 1  pi=207'b000111000011110101100011111010111001101111011000010101101110001001010111111011101101010011110100001000011011100010110001000000111110000001001110111101010111001100111011010110110000111110101100100001101110001;
#1 $display("%b", po);
# 1  pi=207'b011101001111100100011001100011010110100111011010001001110010011010111000100101010010010101110000001111110011000100010010100111101100111110101100011010101111011011011101010011001111001100011111100010001011110;
#1 $display("%b", po);
# 1  pi=207'b111101100011100000011101110101110000010011100100011001011101010001001111011010111000001000000100011101110110010001100010000001001010000010000000001101000110100110001100011110110011000001011010100111010110111;
#1 $display("%b", po);
# 1  pi=207'b001010110011000110001101010011011101111001111001100111000010000111011000010100001001000100110101100001011001101100000011000100001101101100011100001001101101011110011100001000101000010001100101010000001000000;
#1 $display("%b", po);
# 1  pi=207'b110110111001111101011111111010100111000100111010000111101011011010101100101111011001000010011001001111100100111011110111111111001111101100000111101001010001100100100100111111111001110111100001011110110111001;
#1 $display("%b", po);
# 1  pi=207'b110010001101000010111110001010011010110010000101000110110000101011000111101010001101001011011001000010111100100110111011101101000110011001000010110101101000011100010011001001000100101000100000010111011110111;
#1 $display("%b", po);
# 1  pi=207'b110101111001011111010011011101010101010110100101111101100000101011010010001100111011111110110000111000101110011000110000010111001000000001110100110001111111111011101011110101100110110001101101100011010101100;
#1 $display("%b", po);
# 1  pi=207'b001110110010001101001010101010010100010101011101011010111000100110100111011011110010100000000010001110101110000011111001111111000111101111000011111101001111111111001110000011111111001100011100011101100011001;
#1 $display("%b", po);
# 1  pi=207'b101011000101100011001111100111111111111111010100001001111011101010100110000101010111101010011101100011111110100101010110001011000001000001010010100100100111000101100110011111001110010110000101010011001101100;
#1 $display("%b", po);
# 1  pi=207'b100111110100011010101110100100011100010101100001001101100101110010011111001100111110111010000110110111101001110100110000100011011011001000000001111000010111001010101010011110000110000100001100100110111000001;
#1 $display("%b", po);
# 1  pi=207'b010101010101001101100100101010000110100010101001101011100100010100110100111101100110011001111011001101001111110011100100100110110101010111111111110111010001000000000011110000100011001111110010001011000110110;
#1 $display("%b", po);
# 1  pi=207'b000100001101011110100111110010011111010011100000010010010010111110010001110001000100001011111101110011110111111001100001001001101100111010100001001000110010001101010111100101101111110101000110001011100001101;
#1 $display("%b", po);
# 1  pi=207'b111000101111000010011100011001001011001011001001010100100101101110110111010010010000001111000101001111010100111011010011111000100100111110011100011010111100101110010001010101111110111011100101111001011101110;
#1 $display("%b", po);
# 1  pi=207'b110111111111000011101111011101111001010001010001101011011100000011011011111111110000000000101001011000110000000101110001011101011000110110101101001000001101000000110101101100111001010000101111010000001111101;
#1 $display("%b", po);
# 1  pi=207'b000011010011011001110100111100000101101010110110110100101101101101101011101100100010101110101100101111011100001110110100101110101000100001001001010001110101000010110010110001001111000010111011000000100011110;
#1 $display("%b", po);
# 1  pi=207'b110010011100000001110000101011010110001001110111011001111111101010000001000010000001110000010100111000011101110110100110100001101100001110110011011000001010100010111010111110001011111000010000011101010011010;
#1 $display("%b", po);
# 1  pi=207'b001011010011001001010100110101001001110000100000100010101100011101000011011110110111010010101101010000111011010101110011010101001110111001010000101101111001100110010001001001001111011101111000000011111101110;
#1 $display("%b", po);
# 1  pi=207'b001111101011110110110001111010000100011011100111100110010001010101001010101010100100011001110110001011110110111110100000100101001011101100011100101011111001011111101101101111010010110110000010110110101110001;
#1 $display("%b", po);
# 1  pi=207'b010100100100100001111100110100110001001001001110010100100110101001000100111110100100011000001110101010101000101011101101100110101000001101101110110000110111000101011001111110100011000111110111010110110011010;
#1 $display("%b", po);
# 1  pi=207'b011110010110101111010110000101000111110010110011110010011001000000101111101011100111001110111001100101010111001110011110100011001001001001010011011010100111111101000001010000001010101111000111000101110010111;
#1 $display("%b", po);
# 1  pi=207'b010101000110110010110100011011010111111111001000010000101001110110011101100001111111100001011100010111100111010101011000101111111000111101001001101100011100001011011000101000110110000010101010011111010011011;
#1 $display("%b", po);
# 1  pi=207'b001010011111000010101101010100101100010000001011001000010011100110010111111101010110110010001001100011010101010010100011011100111011001010000000101000101010000100011001101001101101011101001110011001011101001;
#1 $display("%b", po);
# 1  pi=207'b111001011011111110011001101101111101000100101101001011100000010111001000010110001011100101001100010010110111100110111101011000100011101001101100010100110100001101101010011100011010000010100100001000111111011;
#1 $display("%b", po);
# 1  pi=207'b101101100000101101100000100110111101010100011111011001001111010001101001110000000011010100010010110100011111011111000111111010010100100010000110001000001001100000010010010010011110001001010100101010010010101;
#1 $display("%b", po);
# 1  pi=207'b011001001111001101101001010000000100100001111001111011011011011010000010000100100100011001010110001101110100011000000011111001000111011011001111011000101101000010100111111100100011101011100110111100110110110;
#1 $display("%b", po);
# 1  pi=207'b111001101101111101000111100011100101110111111010110000111110110111010110110101000110000000111000011000100000111010011100000000001011000100010111111110001010100010000011110111110001111100100111001010011100010;
#1 $display("%b", po);
# 1  pi=207'b011101100000110101110101010000101101100101100011001010001100100100110010110100000110011001110110011101111011111001100011101111011010110011100110101111111000110100111011000001100000100000000011100110000110110;
#1 $display("%b", po);
# 1  pi=207'b100110010110010010010111101101010000011101011110100111110001001111101011010100110011001011011111100110100011011011101101001000101000101010001000001111000000111001101111000001100001110101111010011110111100101;
#1 $display("%b", po);
# 1  pi=207'b100011110000101111011000111110101000110001111100100010111100100110010001111101011110100101110001010001001011011110001011011000111010011101110000011101101011100111100101001011011000011101110011000101001001011;
#1 $display("%b", po);
# 1  pi=207'b100100100101001010010001011111111001000001101011010101111000001000110001011110111110000110111010101111000100110101110110010001010101111111010010001010110101100101000110111011001000100011100010000000011101011;
#1 $display("%b", po);
# 1  pi=207'b010110001001010000010101101101011100011001100111010110000111110000000001110100010001111110110001110110111110001111101110101100110111100111011001111101110100010101111010011001001111011110110101111001000100111;
#1 $display("%b", po);
# 1  pi=207'b011000110100101101011001011100010000111101000110011001110010000111100111010111101101010001101010011100010001001001100101101011010110000111010101011101001001100111011110111000001001000101111110111110001111010;
#1 $display("%b", po);
# 1  pi=207'b001111100011110100101011110111100101101101110001010000111001001000011110011100100000010100011000000010010010110101011001001111000010001010011011000101011100011100001000001010111100111011000000011111101110100;
#1 $display("%b", po);
# 1  pi=207'b110011000001110010110110111101000011111000010111001011100111110111000111110110001001100110110100000100010110111011011100101000010100110110011111000110011100011111101010010100100000111001000111000000100100010;
#1 $display("%b", po);
# 1  pi=207'b010011010010100111111001101001001000001100001101011110000101001001101100101000010011010010101011000010010010111010011001011110000110010101010111000100000100010100000101101010101111011011001101111101111000110;
#1 $display("%b", po);
# 1  pi=207'b101101011011100000101100001101100100011011100010000001110100000111100100101100000111000000110001011110001101111011100111001010010100110101011111100011010101100110011110110001000001110010010110110001100111101;
#1 $display("%b", po);
# 1  pi=207'b001010101100000000001110010011100011010111000111101110100111000110000011000111000111101000110010100011011011111110101010001010011011001110001000010101001000100101101100000101001001111000000100010001110110111;
#1 $display("%b", po);
# 1  pi=207'b111001001101110011101001001111111101111010110011101100110010110011100110101101111000001011001010101100100110010001110000110100100101010010110111011000100110000111110011100110111101110000110011011110010100100;
#1 $display("%b", po);
# 1  pi=207'b010010000101010000100110011010111101100011001001100101101111100001011011110100001100100101101110110000111000010110000100111101100011110001001010101011011000101100010001000110010000000101000101111010100111001;
#1 $display("%b", po);
# 1  pi=207'b011011101110010111100101010101111010111101001100001000001001000110110010011100001100001101010011110100000011011001101010110010100100100100110111000010111000001011011001101110111001110100001000000000101010111;
#1 $display("%b", po);
# 1  pi=207'b010001111100001001100110010011001100000100000111000111011010010110111101110011010010010101000011011001100100110011001110111011001001010010011000011100010001110111100000010011110110100000010100001100110101001;
#1 $display("%b", po);
# 1  pi=207'b000111000010101110110111001111110011111110000011011010000001101011011111010111011100001101010011111010001111010000001000000000100000001001010111010001101110100111111111001001111111010101000101110011100111011;
#1 $display("%b", po);
# 1  pi=207'b010101001000001011001001001101101001101000101100110100110100011101111100001100011110110110110010110110100110100011101000011111000101011011100101010100000111001011111111010110110110001010101001101100001000011;
#1 $display("%b", po);
# 1  pi=207'b010100110100100101010001011010111101001101011110010001101100101010100110110110010110101010110101110010010111100111011011111001010111100111010101000111011101011000011101000001110011101111101111001001111001100;
#1 $display("%b", po);
# 1  pi=207'b101010000011110111110100010111010001010000111100111110100111100100100010000011000101011010010101001011010111011010101011110111001001010100001010000111001110011010000011111011101100100110001001111100010100001;
#1 $display("%b", po);
# 1  pi=207'b110000100110100111101001000101001011111010111101001011011111110001101101101101011101000111001000000110101011101100110011000100000011000000010001100000110001000101010101100011111000110000010000001100111010111;
#1 $display("%b", po);
# 1  pi=207'b100001001000011110101011001000101010110111100011101011011011010001011010010110000011111000111110001000111000001010110011000010011100110000100011110101000001001011011101110111111000100000001110111010001111000;
#1 $display("%b", po);
# 1  pi=207'b011001001101101100100111000010001001001000010010011011100000100000100011101100010011010100111000000110011010110011010111111001000011110111101001101001001011011000011100001100000111000110010100010000110111011;
#1 $display("%b", po);
# 1  pi=207'b011101001101100111010100011100111001001001000111001000111100011010100111110110110000011111001101111100011001101000001110001110110010000010101101011010100011010010000000111011000110101010101100101011010100001;
#1 $display("%b", po);
# 1  pi=207'b110111100111110001001011101101100101110110000011001001100100011000101101100001100111001000000010000010111010011010111110100011001011011111100111110001011000011010010110001010101001101110101010011100010010101;
#1 $display("%b", po);
# 1  pi=207'b011101111010010110100110101001011000011100001001111001000001011111010111000001011110110100010011010011100001011101010011100101101101101110000000110000001111011001000101000010101101010001100110100001111101000;
#1 $display("%b", po);
# 1  pi=207'b111000010110011000011100010010001010110011111111110100111011110001110001001001100101111010101101011011010100000110100111110001001000011001001010111110001111011000010000000100001101111011001100100010100001111;
#1 $display("%b", po);
# 1  pi=207'b110010110010000001110111001011101011100111100111101011011001101110001101100001001111010100111010100001010101110101100101000110011010001011110001000100110000011110011110110011001110010010110101101010100011100;
#1 $display("%b", po);
# 1  pi=207'b111001100011100001001111110011000011111100010101100101101111000110000101001010011101110001111101011011111001000000111001111001110111100000000001101111010111101110110111111111000000010011001111110001111010000;
#1 $display("%b", po);
# 1  pi=207'b110101000101111100101000001111111110111000010001011101110110000011010000000100110010011001001001010110001011011010100000111111010000001011101101010111001001101000111100011001101011110001011101110110100000000;
#1 $display("%b", po);
# 1  pi=207'b000100011000100100111110010101111111001100001110110110001010100010001011111010010100101011101100111000001101100010000111010111111101011111011000000010011010001011101000000100000000011110011000001011100110111;
#1 $display("%b", po);
# 1  pi=207'b000111011000001101000110001100001010000010100001111110111101010110110011001110001110101000010010110010101010101101111011011101100001001101100110111101111000111100101010010011010001110111110110111001111010110;
#1 $display("%b", po);
# 1  pi=207'b111110011001001111011110110001111000011010001110101110000100011110000001110011000110101110101101100001101011101100100101101100010101011100010110101010100001000111011001101010000110010011100000111000100110010;
#1 $display("%b", po);
# 1  pi=207'b100111010011111100110100110111011110100000010011001100100101000100100011101101010101111000101000010111110010110100000100111011100100001010001111010011101100001100110011100001010010011100110101010110111000100;
#1 $display("%b", po);
# 1  pi=207'b101110110011111101111011110110101001100101010010111011100110001011101101101110010001110111000111011001011000110100101111010100011110110100110000001011101001111101101011110001101101100001000011011011111110000;
#1 $display("%b", po);
# 1  pi=207'b101110000011010011010101111010011000110001111110010110000000010010111111010011001100010100101111010101010011001011010001100110010000100101010010011110001111001110000011100100010000111001011111010110000100100;
#1 $display("%b", po);
# 1  pi=207'b111001010000111111010110101010011110001110110011011010011100111001011111011011011100100000100111111010011100001110010110011011110101100110111000001100010110000111010000010000110000000000010100010010111110010;
#1 $display("%b", po);
# 1  pi=207'b111001100011000110101001011010011000111000000100010111101101000100100101100111100000000011100101011000001010111001000100111000001110010001010101000101110001001111000011010011110110010111111101001101100011111;
#1 $display("%b", po);
# 1  pi=207'b110011011011100101010111100010100101101000110110000000110010000011100000011101100001110011110011111101011000101011111011011000010100100111011001001110110101001110111101100000111010000100010000001001011001111;
#1 $display("%b", po);
# 1  pi=207'b100101011010110110111100110111110111101001100001010000110110000010010000010011100011010011011000011010110011101001001011101101011110111110111110100000100100100011101111111011101101111001011010010010111011101;
#1 $display("%b", po);
# 1  pi=207'b101001111010101111010001000101111110111110000001010011100011100000011000111110011111101100110000110101011011011011101011100010110011100001011110101111110111001101000001010100100101010100010011001110010001001;
#1 $display("%b", po);
# 1  pi=207'b111110011111111010011100000010111010101010001011010110100110101100111111100101100011100011110001001001101110000110000101001111111000110111010110110110000100110000000110100001010101010111000011001000101101011;
#1 $display("%b", po);
# 1  pi=207'b100111000100100010111010110101010010010000011110110000111010111001011111000001111110000111101100101111110010111101110100100011101010011001001111101001110001001011100100100100001111100010011001010100110000001;
#1 $display("%b", po);
# 1  pi=207'b010010101101110011001111000111101111110011100111101010100000101000100000100011101101110001001000101010011001000110010011110010101010011010011001000100011001000101100110100001011000000110011001101001101111110;
#1 $display("%b", po);
# 1  pi=207'b110010100111100001100110000011000000011010110110000100110111110001101101110001111100101110110000001111101011011010011000100101001001001101110110001110011011110110110111000101010001000110000000100010011110010;
#1 $display("%b", po);
# 1  pi=207'b000001010010011100000101001110000110000010000010010100100101010000010101001001100111011001010100111110110010111001101010001100101010101100001010100001001100011010100011100111111111000110101110111111101111111;
#1 $display("%b", po);
# 1  pi=207'b110111100100010110001000111011100111100011000011111100101101111101100011000011001010101101111101011000111111101001000101000010100110111100010011100111111010101111101111000111110110110110010000000101001111100;
#1 $display("%b", po);
# 1  pi=207'b110101000010111010110100110110100000010000100100110100001101111001000101110101100110110000001001010101111001001000000101000000111000100001110110011100001111010110111111101011011111111001001011110010100000001;
#1 $display("%b", po);
# 1  pi=207'b111011101010101001010001101000011100101000110100111110111010001101101011111111100000011011011111011110101111010011000001010111011100101100101101111110001111000011100000100011111011011000101001010000111011011;
#1 $display("%b", po);
# 1  pi=207'b100011110000100101010111100000000100111110011101001010111011111100100100010101001011000000100001001100010000111010001000111001000100000111000000000101110000110101101000000000110011000001010011011000010101011;
#1 $display("%b", po);
# 1  pi=207'b010100100010001011010101000011000001000110000110110001011100110110011010001011101101111110100100010000000110110101011101100101010000000111001110111011100000100011100111000101001101001110100011100011100101011;
#1 $display("%b", po);
# 1  pi=207'b010111110100011010000000100010010111111110001011101111101111001001011110010110010110011000110001001011011011000111000101011101001110100101000110100110100100111101100011100001000011010010001101100111010001111;
#1 $display("%b", po);
# 1  pi=207'b100110101110000001010001111111100110100100100100001100000100011101011000111100100100111100101001010100000001111110001100001000111001000100110101011000111100100011011100010101010110011001001001011001100001100;
#1 $display("%b", po);
# 1  pi=207'b011011001010010000111110000100100111100001111111001010001011100101010111111100101001100000001010111110100100111010100011001000100010010100001100111101101110010000101111100111011010111110000011100111001111010;
#1 $display("%b", po);
# 1  pi=207'b110101000000110110101111110101101001000111100110000101011011011011111011011110000001000100101011010011110100101110010000111011001110011010101010111010111000100001110100000011100010011111110000000011110100110;
#1 $display("%b", po);
# 1  pi=207'b110011010110000011110100111010110010010100100100110111100011101101110101001010011000100001001110011100001011110010110000111111010101111111010010000001001010111100010001110010000101100101011010111011100110001;
#1 $display("%b", po);
# 1  pi=207'b101111001100001111001000011000011100100000010000110100101001000101111000101010010000111101110011001000000000100001001011010000010001001110001010100101100010011110111001110110101010010010010111011000100101100;
#1 $display("%b", po);
# 1  pi=207'b011000011111001001000111100101011000111000100011110110011110101111000011111101010100001111100110000101001000001101100001101110111100100110111000110011101000011110010101011101101000001011001001011000110001001;
#1 $display("%b", po);
# 1  pi=207'b010000000010100000111011011110000110011011000011010011111011110110110111100011010000101001010011100011111111010111110111111011101101010110111101010100110011010100101101110001011100111110010100101110000000000;
#1 $display("%b", po);
# 1  pi=207'b001011111010111011010011000010011101100001100001000111111100111010010010000101110000110011110010100101001010101111010000001011011000000010111101110000001011110100011101100000110111001111010100011010110100100;
#1 $display("%b", po);
# 1  pi=207'b111010100110000110011100100111010100011011111001010011010111011010101000010001011001000101100000111011101010111011000101100010001100000110001111100000111111001011011010010101110001111001101001110000111010010;
#1 $display("%b", po);
# 1  pi=207'b011000000010101011110100100111000000011001000001100101110010010110001010101000110100111001100110100011100000000101101001010010111011010110000111011010110010110011111110110011011100010101111000001001101010011;
#1 $display("%b", po);
# 1  pi=207'b101110010110100111010110111001001101000010001000110000001000011101011100111000000100011111010101100100000110101111101101100001100010111110000110001110101000000000010101101111000100011111011110110010011000000;
#1 $display("%b", po);
# 1  pi=207'b011001011111100010101110110001111000111100000010000100100010111111101101111110111010001110110001000110010100101110100000101011101111011101110101011011110101011111000110101010000001111010100001010000110011110;
#1 $display("%b", po);
# 1  pi=207'b111110010000001111101011011101010111110001000000010001010110001110001111010100100111000101001100101110001001110001011011001100111011101110011011010111001011100111011110010110100100011111010001010100010000011;
#1 $display("%b", po);
# 1  pi=207'b001000001011100100000011010101101010000110001101010010111111011111011010011000110101101001111101001100111101101001100110010101001011011111100110110110010000001110010000101100100101000100110110000010100110100;
#1 $display("%b", po);
# 1  pi=207'b001101110011001001001010101001010010110111010110000000100101101100001000011001000100110010010100111111000100000010100111101100101000010101110011010110000010000010110100001111001111111111000000111100101100110;
#1 $display("%b", po);
# 1  pi=207'b000101110011100010101100001001011101100111100000101111100011001100100010011010011101001010110010010111111000010110111011110000011110000010001010010111101010010010111111101101010111010101000000111000110111110;
#1 $display("%b", po);
# 1  pi=207'b011111111100101011010011100011001011010110101001111001110110110100001010000110011001101001000100111111110100100101001001011100100001000101010110100011111000111111101110111000101111010010100001000010001000111;
#1 $display("%b", po);
# 1  pi=207'b001110001110111111100110110010100010101101110110010010001101000110001010010001011010011011111001110101101111011000111101100001000000000011000110101011100000000110111110011100000111000100001001011110110110100;
#1 $display("%b", po);
# 1  pi=207'b001110101110010001000011100101101001100001010010110011000111001000000111100110011000101110101000001011010011011011101111100110111010000011001010101110110010011011101100111100000001001111111100011001101011100;
#1 $display("%b", po);
# 1  pi=207'b011111100100101100011100001001000110111010110101111010110110010101100010001011000101000101000011000001111111101101011000111001111010100100000010011111110100101110100111010101101001010100000001000010100110000;
#1 $display("%b", po);
# 1  pi=207'b011111001010110111110111100000111100101110000011101000010000010110101011010111110110010010101101110011001001000010011110010111001001110111101010111000000010110010001001101110010111100101110010111100100010000;
#1 $display("%b", po);
# 1  pi=207'b001011001010111111111010000111100010111011001110101100111111010000101101111110011110100110110100010000110000000110110010010111011101001010001101100111101111001101000001101110101111001101101011101110100001011;
#1 $display("%b", po);
# 1  pi=207'b110011100000001000101001010111101000010011100111000011100001100101111111010100010010100011101100110111110011001101100110101100101000011000110101110000010101001100101100001100000010010100010000000101010000100;
#1 $display("%b", po);
# 1  pi=207'b100011110101100100110101100010000111010011000001000111111011111100100001010010101000001010010110000001000001110001011110011010111011000000111100100111011100010111000101110111100110010110011011101011100011111;
#1 $display("%b", po);
# 1  pi=207'b111111100101010000010010000101100111011001101000111000100000000010010101111110110111101111000111010101010111111100011011110110001111100110010010100111100110001010100111000111110101100001110111001101011100010;
#1 $display("%b", po);
# 1  pi=207'b100011100001101001011111010010111101110011010011101011100110001101010111111101101110011000111100100001001110000111110010001100000100111101110110001110111010110001110111100010111001001000101101000110111110100;
#1 $display("%b", po);
# 1  pi=207'b110011101010100010000100001001110010000111011000101111100100011111010111100110001010011010100101110001000011000110000101000100010100111001111011111001011111110101000100110101000110100010110110000000110000100;
#1 $display("%b", po);
# 1  pi=207'b011011111000101100000011000010011110001011110001011001010101101100010011101110000100100000100111110111001111011010011100000001111010100010101111101011101011001001101110001100100111011000111010011011111011000;
#1 $display("%b", po);
# 1  pi=207'b111011000111101000001110001100000101101110111000100010101011011100111101000011000111001111000000010101100010110111110110001000001110110110100001010010100011011010010000011010111011010001001101110001011110101;
#1 $display("%b", po);
# 1  pi=207'b000110000110010000110010001011111111101010001000101111010101111001100111101011111010100011101100001000110000010100011110001110001011111110111000001110100101011101100100010111111100110111010011010011101100110;
#1 $display("%b", po);
# 1  pi=207'b010110001011111000110011001011011101001110100000100101110010000001011101000111001100011101101101100010001110100100100101011001000011101110010100011001111001010000000001000000100101001001000101100111101010000;
#1 $display("%b", po);
# 1  pi=207'b101111011001110111110101110000111100110100000000001001010001011000110110110111101100101010101010110000000111010000101011111100010000001101110011110111011011001100001101101000111110111100100011101001111101110;
#1 $display("%b", po);
# 1  pi=207'b001100010000010101101000011000101100000011100001111000100111011001011101000101000100010111001101101010110110101010111100011111110001111111001000100011010101110111110001100000101111011000110000100101100111011;
#1 $display("%b", po);
# 1  pi=207'b100000011101101010110100111101001100110001110001111101000101110001110010111110010101011111000000001001001110101010100010101010100101110110011011111111101111000110101001111011011001000001111000010010001000000;
#1 $display("%b", po);
# 1  pi=207'b110000100001010110011110001111111001011110010110000001110110000010001101010100111100110111010001011010111000111111111010011001101110100101110001110101000100011101101000110110100010000000110001101111101010011;
#1 $display("%b", po);
# 1  pi=207'b110100001001110011011111000011111010000000100101101110111110000001101101101100000110011000011001000111101100010000101101000110001110011100011011110010100101110110011000010101000110110110101011011000001110100;
#1 $display("%b", po);
# 1  pi=207'b110010101010011111101110010110101110000111001001010110111011101011111000111011000000110001010010110100110111110110000101011100100110100110111001111010000011010011000010111100111101011010110100111001101000010;
#1 $display("%b", po);
# 1  pi=207'b101100001100100110110001011011001000001011000100010110110011100011010101110001101111011110101110000110011011100011000111100010001000110110100011010111001100001000110110110001000110100011100010000101100100001;
#1 $display("%b", po);
# 1  pi=207'b101111001000111111111100101101001101000110011000111011011010001000011001110011110011101101000111010010111000100000110111001111111100100111100111100111110000101000011111001010111001100100110110100110011001101;
#1 $display("%b", po);
# 1  pi=207'b001101111100001011001010110010100100101111100001111110100101111101111101001100100010001100001111000101111101010011001000100100110010111100001101100100100111011111001100010110011101010111011100011001000100000;
#1 $display("%b", po);
# 1  pi=207'b110111111010110110000110111010010010010101100110101000110010000111001101101111001011001011000010000001100001000010001100010010010100110000110110100101000000101110110100000010011000010010101011010011011010010;
#1 $display("%b", po);
# 1  pi=207'b001101101000111001100100111011111000110001010000111100111010100110110010101010100100101011011101100001000110101100000110001011111000100011101101011110010001000001110011010101000110011101111010100000110101001;
#1 $display("%b", po);
# 1  pi=207'b011110000101111100110101000100010101101001111100011100111100010111011111000100001101110011000011111101011110100000010101110000111010011100010111010110001000101111110100110110110101101010000101010101111100111;
#1 $display("%b", po);
# 1  pi=207'b010111101000000100101010111110010001011011110001001011011110011100101101110110010000011111011111010111001111001010010111010011011101010011101010101010010001111101011011011000101101001110110001100101101011011;
#1 $display("%b", po);
# 1  pi=207'b101110111011000010010111110011000001010000100010111110111000001011000101110001110100011000100000000001101000110010000111101011101000110010111001111101010000010011110110010001110011101000110010101010011011100;
#1 $display("%b", po);
# 1  pi=207'b111110011011001000100010100100100010010010111101000010000001101101000111000110000001010110100011101100110101001110110010110101111011101001110000010011000011001101111010100001111000000101011010111101110101100;
#1 $display("%b", po);
# 1  pi=207'b110111111111000001101110111111111111000101010110001101111010000001000100110100101111001110110010011000101110111111101001001000010110101111101101110100000101101011101000111010001010000010010011010000011000110;
#1 $display("%b", po);
# 1  pi=207'b011010001001100001011011000010111000110100011001101001001000110111011101000101100000000010100000011011101001101100101101011110111110000100101100101001101110110011000011010101011110000110101000101000110010111;
#1 $display("%b", po);
# 1  pi=207'b001001110000011111111101100001100011010010101101101110011100011011111000100000110110110111101001110000000010110111111010000001011100001111111011000100110101101110111111101001111010001111100101011111011111000;
#1 $display("%b", po);
# 1  pi=207'b110111010010111010100100010110001000001000111111111111010000010110010111100001011000111011111000001000000111110000101011001001100000000011010010011110000100101101110001100001101010010110110111101101110111111;
#1 $display("%b", po);
# 1  pi=207'b100101001000001010011100101001011110101101011100110000100011101111110100111010100100010101011110011010001000110100111000010011001001111000100011111000100100111110000000011110010111111010111101011011000011100;
#1 $display("%b", po);
# 1  pi=207'b111011011000001110111101100111110101010000001000010110110100010011100010011010111011110010111111010110111111010101110100000001011101101101000000111000101000011011000101111001000001011001100101010000001101001;
#1 $display("%b", po);
# 1  pi=207'b100010011011110001110110010111011100111010011001011101011001110101111110011111001001001101011010100010101111000001010000011110110010001100101000000101001001101001010110000000111100111100010111000001000010011;
#1 $display("%b", po);
# 1  pi=207'b101100111010101000100100010000000010001110001010011011011011000010101110000011111010111101001001001010000010100101110011101111110100110101110000000001100100011011011101111110100111010101000111110011001111010;
#1 $display("%b", po);
# 1  pi=207'b100001000000000101011110011110010101110111101101001110000100010010000000110111111000100011010011011101100010110011001100100000000100001111111110100000101111101011000011000110101100001010000010111100110010110;
#1 $display("%b", po);
# 1  pi=207'b100000111111101101111100100001101100011001000110111101011001011111100000000110101010001010010000110100111100001001100001110001000101100101111010101000111100000101000100001111110101001111101101010101010101000;
#1 $display("%b", po);
# 1  pi=207'b110110101111111001011001101100101101110100010101101101010010000110110100110000010100011110111000000101100110111111111101000101111000001011001100111011101100000001100100101100101100000001110100001001110000000;
#1 $display("%b", po);
# 1  pi=207'b110010011001101010110000111001111110001010110010001001110010111010000100101011110101011110000101100001001000011010101101001101100111100111101100100111000000010010100011111001100001001000011101001111100010000;
#1 $display("%b", po);
# 1  pi=207'b111011110110110101010101110000111011101100010110100111100000011000001011010000101110001000100011001010111110101110100100100011011010011010001001011010111111011110000111001010011000110000011100001000000101111;
#1 $display("%b", po);
# 1  pi=207'b010110011001001010010110100000100110111000101001111100100010110011001111010110011110110111000011110100010011100100110010010000101011101111000100010100001000001000010010010010101110001001010001000101111101001;
#1 $display("%b", po);
# 1  pi=207'b111111111111111110010111100111011001001011111100101100100010000100111100000001111111001001111010100001111010110101110100101001000011101111110001011111111011000111110000110111100000011111010011111011001111010;
#1 $display("%b", po);
# 1  pi=207'b111011101000010011001100100011111010100110001010110111101011101110000001111110011010110010000001001111110111001110100110100000110011001001010100001010100001101010110001010011100000100010110001100001110001111;
#1 $display("%b", po);
# 1  pi=207'b111111111100001100100100100011000100001110100000101001010011010010110001101010110010100100010101110010001100000110101100111111100100000011001010101011111001010010101000011111111101001110001000101111000110001;
#1 $display("%b", po);
# 1  pi=207'b100111000111101111101100011001001100000000001001101010011111011111011001011011010011111000100000100111100011011100010100000000001111100110001011000000000010011100000100110111100110111110110011101000111100010;
#1 $display("%b", po);
# 1  pi=207'b010110011001010000011010001100000000111101111100100000111000011011101001011100001111000001001001101111001110111000010101000011001000001110110011111101000000010100111111001101001011101111110001001000101110010;
#1 $display("%b", po);
# 1  pi=207'b110011110111011011000110011101101100111001100110110101011001101000000110110100100010110111011010010001111111110111111010010010111010110111011001010101101000100100100000111010010000010011111111110000001010011;
#1 $display("%b", po);
# 1  pi=207'b110111000010011101111010010011110011100001100100111100011100110001111011101111101111001011110110110100111011100100101110101111101111000100101001010001100111011001111101000100101101001000110110010100110100001;
#1 $display("%b", po);
# 1  pi=207'b001010011010110111100010111001110110001010010101100011111101000111001111000011010001101011010101100001000101011111101011000011000110000110110100111011100110100010111011001010010001001011100010011011110111010;
#1 $display("%b", po);
# 1  pi=207'b110111100001111100010100111100000110110011101110111111010111001000000000101110100100101010011000000001110110000110101100010111000101010000000011011001110011001000111000010101001111110000111110001000001110001;
#1 $display("%b", po);
# 1  pi=207'b101111101100111111011011000000111000111100111010011001001100000111000111001111011100010101001010010111111111111110110100000110111101011100001001000110010110010110001110110101000111001101010011000000100110100;
#1 $display("%b", po);
# 1  pi=207'b100010001000100110111001100001101111010101011110001011000011110000100100001111011101101101001111110000100001101101000111100000000011100111001010011010000000100011011110100111011001010100000100010000111101100;
#1 $display("%b", po);
# 1  pi=207'b010101100000010110001111101101011111101001101001011000100101111110000010011000001000111010001010001111010000100001100101011101111110001111100101011000111110100011101111011000101001100111100111001111111010111;
#1 $display("%b", po);
# 1  pi=207'b101001011111001101011011111101000000010010101000111001010010110011100110111010010001010010111000101010101000111011100101101010100100000010010001000000111010011011011100011001011110100111011011101011001010100;
#1 $display("%b", po);
# 1  pi=207'b000001100111101011111000000000000101101011011100100010111110110000100010010100100100111100000111000101111011110010110101110011010011111011000101000101111010101110111101011110000011000110010001010100011111111;
#1 $display("%b", po);
# 1  pi=207'b101100101100011101010011110111111100111011010001110010111101010000101101011001110000110101011011000010011111000110100010001010110101011011000010101100100110111010001100110001101101011101001101101101101001010;
#1 $display("%b", po);
# 1  pi=207'b001011111100000111011101101011010100000000000011101101111101101110101110100101111000000110010011101100011010110101000110100000110100101011101111111000000100011101110101010101011010111111101011001010010110000;
#1 $display("%b", po);
# 1  pi=207'b001010100011000111000011011110101010010000011101000110110110010010110101000000110111010010100001100001111010001111100111110100110000110111011101101010000100100111110100110000010011010101111000110001100011110;
#1 $display("%b", po);
# 1  pi=207'b011011000010011011100010101110010101001010001101100100000111001000101001100110110110110000000101111101000011000111101010001100101010010101110101010111001101010010110100010111001101001001000001111000011101101;
#1 $display("%b", po);
# 1  pi=207'b010010101001011101000010101110001011101010001000000110001111011110011110011000011110110111010000110101010000101110001101100000101110100011100010001000111011110001010001100110101010010100000010011001011001101;
#1 $display("%b", po);
# 1  pi=207'b000010011110100010010100110011011100010110001111100100000101000000101011111010100110101101110000000110001000010111010011001011011111001101100000000001110011010101110100010110011000100111001100111001110001010;
#1 $display("%b", po);
# 1  pi=207'b011011011011000111100001000011001011101011100010011011000010001110001110100110101011000001001010110110000111001001011110110111000100001111010011010100000100011001010001001100011010000110111111101001110010101;
#1 $display("%b", po);
# 1  pi=207'b010100110101101000101111111111111011111110001110000010101011001111111101101100100001001100100100110100010001000000010100000001110101000101010001100101000101011100001110000100001010110111100011001101110000010;
#1 $display("%b", po);
# 1  pi=207'b001010010011111011111111011101101011111111001111011010111111101011001111110001110010000100101000110101001001010111100000000111011110111100010000100101111101000010101100100000011000011010001101011111001100101;
#1 $display("%b", po);
# 1  pi=207'b000011010101111001100010100101001000100000010001101000101011100011010110101010011001101011111011100110000110100001000010101100100110010001001101001001101101001101110010100101101001111010111000100111000100110;
#1 $display("%b", po);
# 1  pi=207'b100001010110110101000101101000011011110111110010000110111111111100110000100111010001101011100111101110000001000011111101000110010000001010101000110001100110011111100001101111100001110111101001100010111011010;
#1 $display("%b", po);
# 1  pi=207'b100010010101000110110011001100100101011101011101001000100100101000001111011011110110000000001100110001111101111010000110000001100001001110000000001111111100101111110011011101001001110011010101111010001111010;
#1 $display("%b", po);
# 1  pi=207'b100010010101001010001111111001000110111111010010110110001110111010101101000010010011110010111010000010110111100101010111101011001111011001110010111000100100100010100011110010111100010011111000110011011101101;
#1 $display("%b", po);
# 1  pi=207'b010011000110101111110111111001001100101011101010001010101011001011101010100100100110101110101111011011111011000111100011001111001000010010110010111101000110110000000110100101111101100001000001000001011111110;
#1 $display("%b", po);
# 1  pi=207'b100001010111100110000101100011100011010100110011000011110000111111001011101001000010011011010001011110011101000101111110100101011011101010010111001011000001110001000100001011100000000100110110001100101001000;
#1 $display("%b", po);
# 1  pi=207'b001011010110110100001110011001001110111101111001010011011100101100001110100001010110100101100010111100011010010110010010101111011111011001111110010111011001010001101110101000000101011111011001110001000010110;
#1 $display("%b", po);
# 1  pi=207'b111000000010000001110011000101100111100110111111100101011011011010010011000001011011001100101000011000000010101000100000001100111011000110101111001111010010010101100000100000010000110010100001100001101000101;
#1 $display("%b", po);
# 1  pi=207'b011000101001101101100101101101110100011010110011111111101100000011010111001110000001111111111001010000101100001101110010110101011010101101001100100100110100101101110110011010011100110000100100101100110011111;
#1 $display("%b", po);
# 1  pi=207'b010010000011110001000011000011101100001000000010011000101110001101111001000100001100001100100100101101111110010110000011001101010110111010001110101001001101110010000000000101101111111100100100100000111100100;
#1 $display("%b", po);
# 1  pi=207'b010110001110110111110101010010010111110110011010111111100110110110111101111001001111110100111100100011010000110011100000011001000001101011001001100010001110001100100110100100000111100101101001101101010001110;
#1 $display("%b", po);
# 1  pi=207'b001000001001010010000001111111111101001110000010001010010101101011111111100100111100001110001100101111001110010000111010100101001001001101001000000000011110001010111101000100111111101100011110110001001010101;
#1 $display("%b", po);
# 1  pi=207'b010011100111000010001000011000010001001110000000101111011101111001010001010011110100110110100010100111101010000100100100110100011100101100110111001111000111000101010100000111001010110010001000001110110100000;
#1 $display("%b", po);
# 1  pi=207'b110101110001110101010001110000100100100101000001000011010011101110110011100000101011101110010100001111100011101110010001111011111101001000100101010100000101011100111111011000001100101110011000110110001011001;
#1 $display("%b", po);
# 1  pi=207'b111001000101101101011101001111100010010110011101110111111010011101101001010001100101110010001100100101101011011110101110110011100100100000001011100101010101010010000110011111011000111110000111011101011111101;
#1 $display("%b", po);
# 1  pi=207'b101001110100110100010000011101111111110111011001001110111100010000100000110001110011100100111100011000100110101110100011100110101101100001101101001010001111010000110000001111010110000011101000001100100111001;
#1 $display("%b", po);
# 1  pi=207'b000010111000101110101010000001100100101110011011010001100000011101001111110110010010001101100100001000010010001100110001011011011010010010110100101100001011101010001010101100100101110001101000110111101111001;
#1 $display("%b", po);
# 1  pi=207'b001000001001101011001111101010110101010110011001000010101100001110001110110000100010100000001101110001010101001011100100001100011000110001101001110101001010100010100100110011101111100000101001101001110001110;
#1 $display("%b", po);
# 1  pi=207'b011000110111000101010101111001011101100110101011111100110110101110110000100001111101111000100010011101101101101001111110011001011000110111001101100111010000100101011001000000111100100000110011101010111111110;
#1 $display("%b", po);
# 1  pi=207'b101101111101000110001110011111001111100011110100110100011000100101001001110101110000001010101011110111111100101100000000010111011001100010101000011011111010011100001001100110011001101101111010101010101001110;
#1 $display("%b", po);
# 1  pi=207'b000010110001000000110101101100101010100000101011000001111000100111001001011110000111100111001100001101110101010011101010100010001101101100011000000011110001100000001100001101010110010100110110111010100011010;
#1 $display("%b", po);
# 1  pi=207'b111100010111011011001111100111110000000001101010110000001110110001000010100010000100000010001101001100101000100010101100000010000011110000010011101001010001001100001111101100101000000101010110000100000000100;
#1 $display("%b", po);
# 1  pi=207'b100100111110110000111000000001011101000110110001010000111001101101001011000000101110110111011001101011001101000100011101111000011011000010110100001000011010110010101011101011110111000010111001010011100010011;
#1 $display("%b", po);
# 1  pi=207'b000111001010101011000001111100111011100101110001111101100011000111101101011110010100001000001010101100100010101010000010100010011000010010001011100011111000001110110000111100100100001001010001110010011111110;
#1 $display("%b", po);
# 1  pi=207'b000111011001111001000100111101011111111010001000110111100101101011000101100010000011100011001101001110001011001100101010001000100100011111010010010010110000100110000100101111111010001111001010011100000101000;
#1 $display("%b", po);
# 1  pi=207'b101011010100101101011001011001100010101110010110000001101110000001011001000101001011000100111111001110100010101100111011000100010001111111011010100110100000001011100010111110010011110101001110101000010100001;
#1 $display("%b", po);
# 1  pi=207'b111110110010011011011011010111100110101101101000101100000001001010000011100110100101001010101110000010011010000011100101110100100001001111000001101000001111111010110001000010111111010110011111111100100000100;
#1 $display("%b", po);
# 1  pi=207'b100101110110001111000100100001011000001001000101000001100101000001100000110100001111100110010111110100001010111100010011011110110001100110110000000001001000001100110001100101001010101111011110001010011011010;
#1 $display("%b", po);
# 1  pi=207'b111101101011111001000110100001010111111111001100011011000110111011001001111011011111001000100011011101110101100010111101001000001101010011111010111100010001010010101100100101110010111111001001110101101110111;
#1 $display("%b", po);
# 1  pi=207'b011010110110000011000110100010111011100101110011011100110010010110011111100000110001000101001101101000101010100000011110101100111110011011010110100101011100100100101100001000000010100001011111010100110001011;
#1 $display("%b", po);
end
endmodule
