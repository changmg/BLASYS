module adder32(\in1[0] , \in1[1] , \in1[2] , \in1[3] , \in1[4] , \in1[5] , \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] , \in1[11] , \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] , \in1[17] , \in1[18] , \in1[19] , \in1[20] 
, \in1[21] , \in1[22] , \in1[23] , \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] , \in1[29] , \in1[30] , \in1[31] , \in2[0] , \in2[1] , \in2[2] , \in2[3] , \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] 
, \in2[10] , \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] , \in2[16] , \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] , \in2[22] , \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] , \in2[28] , \in2[29] , \in2[30] 
, \in2[31] , \res[0] , \res[1] , \res[2] , \res[3] , \res[4] , \res[5] , \res[6] , \res[7] , \res[8] , \res[9] , \res[10] , \res[11] , \res[12] , \res[13] , \res[14] , \res[15] , \res[16] , \res[17] , \res[18] , \res[19] 
, \res[20] , \res[21] , \res[22] , \res[23] , \res[24] , \res[25] , \res[26] , \res[27] , \res[28] , \res[29] , \res[30] , \res[31] , \res[32] );
  input \in1[0] ;
  input \in1[10] ;
  input \in1[11] ;
  input \in1[12] ;
  input \in1[13] ;
  input \in1[14] ;
  input \in1[15] ;
  input \in1[16] ;
  input \in1[17] ;
  input \in1[18] ;
  input \in1[19] ;
  input \in1[1] ;
  input \in1[20] ;
  input \in1[21] ;
  input \in1[22] ;
  input \in1[23] ;
  input \in1[24] ;
  input \in1[25] ;
  input \in1[26] ;
  input \in1[27] ;
  input \in1[28] ;
  input \in1[29] ;
  input \in1[2] ;
  input \in1[30] ;
  input \in1[31] ;
  input \in1[3] ;
  input \in1[4] ;
  input \in1[5] ;
  input \in1[6] ;
  input \in1[7] ;
  input \in1[8] ;
  input \in1[9] ;
  input \in2[0] ;
  input \in2[10] ;
  input \in2[11] ;
  input \in2[12] ;
  input \in2[13] ;
  input \in2[14] ;
  input \in2[15] ;
  input \in2[16] ;
  input \in2[17] ;
  input \in2[18] ;
  input \in2[19] ;
  input \in2[1] ;
  input \in2[20] ;
  input \in2[21] ;
  input \in2[22] ;
  input \in2[23] ;
  input \in2[24] ;
  input \in2[25] ;
  input \in2[26] ;
  input \in2[27] ;
  input \in2[28] ;
  input \in2[29] ;
  input \in2[2] ;
  input \in2[30] ;
  input \in2[31] ;
  input \in2[3] ;
  input \in2[4] ;
  input \in2[5] ;
  input \in2[6] ;
  input \in2[7] ;
  input \in2[8] ;
  input \in2[9] ;
  output \res[0] ;
  output \res[10] ;
  output \res[11] ;
  output \res[12] ;
  output \res[13] ;
  output \res[14] ;
  output \res[15] ;
  output \res[16] ;
  output \res[17] ;
  output \res[18] ;
  output \res[19] ;
  output \res[1] ;
  output \res[20] ;
  output \res[21] ;
  output \res[22] ;
  output \res[23] ;
  output \res[24] ;
  output \res[25] ;
  output \res[26] ;
  output \res[27] ;
  output \res[28] ;
  output \res[29] ;
  output \res[2] ;
  output \res[30] ;
  output \res[31] ;
  output \res[32] ;
  output \res[3] ;
  output \res[4] ;
  output \res[5] ;
  output \res[6] ;
  output \res[7] ;
  output \res[8] ;
  output \res[9] ;
  top U0 ( .pi00( \in1[0] ) , .pi01( \in1[1] ) , .pi02( \in1[2] ) , .pi03( \in1[3] ) , .pi04( \in1[4] ) , .pi05( \in1[5] ) , .pi06( \in1[6] ) , .pi07( \in1[7] ) , .pi08( \in1[8] ) , .pi09( \in1[9] ) , .pi10( \in1[10] ) , .pi11( \in1[11] ) , .pi12( \in1[12] ) , .pi13( \in1[13] ) , .pi14( \in1[14] ) , .pi15( \in1[15] ) , .pi16( \in1[16] ) , .pi17( \in1[17] ) , .pi18( \in1[18] ) , .pi19( \in1[19] ) , .pi20( \in1[20] ) , .pi21( \in1[21] ) , .pi22( \in1[22] ) , .pi23( \in1[23] ) , .pi24( \in1[24] ) , .pi25( \in1[25] ) , .pi26( \in1[26] ) , .pi27( \in1[27] ) , .pi28( \in1[28] ) , .pi29( \in1[29] ) , .pi30( \in1[30] ) , .pi31( \in1[31] ) , .pi32( \in2[0] ) , .pi33( \in2[1] ) , .pi34( \in2[2] ) , .pi35( \in2[3] ) , .pi36( \in2[4] ) , .pi37( \in2[5] ) , .pi38( \in2[6] ) , .pi39( \in2[7] ) , .pi40( \in2[8] ) , .pi41( \in2[9] ) , .pi42( \in2[10] ) , .pi43( \in2[11] ) , .pi44( \in2[12] ) , .pi45( \in2[13] ) , .pi46( \in2[14] ) , .pi47( \in2[15] ) , .pi48( \in2[16] ) , .pi49( \in2[17] ) , .pi50( \in2[18] ) , .pi51( \in2[19] ) , .pi52( \in2[20] ) , .pi53( \in2[21] ) , .pi54( \in2[22] ) , .pi55( \in2[23] ) , .pi56( \in2[24] ) , .pi57( \in2[25] ) , .pi58( \in2[26] ) , .pi59( \in2[27] ) , .pi60( \in2[28] ) , .pi61( \in2[29] ) , .pi62( \in2[30] ) , .pi63( \in2[31] ) , .po00( \res[0] ) , .po01( \res[1] ) , .po02( \res[2] ) , .po03( \res[3] ) , .po04( \res[4] ) , .po05( \res[5] ) , .po06( \res[6] ) , .po07( \res[7] ) , .po08( \res[8] ) , .po09( \res[9] ) , .po10( \res[10] ) , .po11( \res[11] ) , .po12( \res[12] ) , .po13( \res[13] ) , .po14( \res[14] ) , .po15( \res[15] ) , .po16( \res[16] ) , .po17( \res[17] ) , .po18( \res[18] ) , .po19( \res[19] ) , .po20( \res[20] ) , .po21( \res[21] ) , .po22( \res[22] ) , .po23( \res[23] ) , .po24( \res[24] ) , .po25( \res[25] ) , .po26( \res[26] ) , .po27( \res[27] ) , .po28( \res[28] ) , .po29( \res[29] ) , .po30( \res[30] ) , .po31( \res[31] ) , .po32( \res[32] ) );
endmodule

module top(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63, po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32;
  wire n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, tpo00, tpo01, tpo02, tpo03, tpo04, tpo05, tpo06, tpo07, tpo08, tpo09, tpo10, tpo11, tpo12, tpo13, tpo14, tpo15, tpo16, tpo17, tpo18, tpo19, tpo20, tpo21, tpo22, tpo23, tpo24, tpo25, tpo26, tpo27, tpo28, tpo29, tpo30, tpo31, tpo32;
  assign po00 = tpo00;
  assign po01 = tpo01;
  assign po02 = tpo02;
  assign po03 = ~tpo03;
  assign po04 = tpo04;
  assign po05 = ~tpo05;
  assign po06 = tpo06;
  assign po07 = ~tpo07;
  assign po08 = tpo08;
  assign po09 = ~tpo09;
  assign po10 = tpo10;
  assign po11 = ~tpo11;
  assign po12 = tpo12;
  assign po13 = ~tpo13;
  assign po14 = tpo14;
  assign po15 = ~tpo15;
  assign po16 = tpo16;
  assign po17 = ~tpo17;
  assign po18 = tpo18;
  assign po19 = ~tpo19;
  assign po20 = tpo20;
  assign po21 = ~tpo21;
  assign po22 = tpo22;
  assign po23 = ~tpo23;
  assign po24 = tpo24;
  assign po25 = ~tpo25;
  assign po26 = tpo26;
  assign po27 = ~tpo27;
  assign po28 = tpo28;
  assign po29 = ~tpo29;
  assign po30 = ~tpo30;
  assign po31 = ~tpo31;
  assign po32 = ~tpo32;
  adder32_0 U0 ( .pi00( pi07 ), .pi01( pi08 ), .pi02( pi09 ), .pi03( pi10 ), .pi04( pi11 ), .pi05( pi39 ), .pi06( pi40 ), .pi07( pi41 ), .pi08( pi42 ), .pi09( pi43 ), .pi10( n1 ), .po0( tpo07 ), .po1( tpo08 ), .po2( tpo09 ), .po3( tpo10 ), .po4( tpo11 ), .po5( n2 ) );
  adder32_1 U1 ( .pi0( pi12 ), .pi1( pi13 ), .pi2( pi14 ), .pi3( pi44 ), .pi4( pi45 ), .pi5( pi46 ), .pi6( n2 ), .po0( tpo12 ), .po1( tpo13 ), .po2( tpo14 ), .po3( n3 ) );
  adder32_2 U2 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi02 ), .pi3( pi32 ), .pi4( pi33 ), .pi5( pi34 ), .po0( tpo00 ), .po1( tpo01 ), .po2( tpo02 ), .po3( n0 ) );
  adder32_3 U3 ( .pi0( pi03 ), .pi1( pi04 ), .pi2( pi05 ), .pi3( pi06 ), .pi4( pi35 ), .pi5( pi36 ), .pi6( pi37 ), .pi7( pi38 ), .pi8( n0 ), .po0( tpo03 ), .po1( tpo04 ), .po2( tpo05 ), .po3( tpo06 ), .po4( n1 ) );
  adder32_4 U4 ( .pi0( pi24 ), .pi1( pi25 ), .pi2( pi26 ), .pi3( pi27 ), .pi4( pi56 ), .pi5( pi57 ), .pi6( pi58 ), .pi7( pi59 ), .pi8( n8 ), .po0( tpo24 ), .po1( tpo25 ), .po2( tpo26 ), .po3( tpo27 ), .po4( n9 ) );
  adder32_5 U5 ( .pi0( pi28 ), .pi1( pi29 ), .pi2( pi30 ), .pi3( pi31 ), .pi4( pi60 ), .pi5( pi61 ), .pi6( pi62 ), .pi7( pi63 ), .pi8( n9 ), .po0( tpo28 ), .po1( tpo29 ), .po2( tpo30 ), .po3( tpo31 ), .po4( tpo32 ) );
  adder32_6 U6 ( .pi0( pi15 ), .pi1( pi16 ), .pi2( pi47 ), .pi3( pi48 ), .pi4( n3 ), .po0( tpo15 ), .po1( n4 ), .po2( n5 ), .po3( tpo16 ) );
  adder32_7 U7 ( .pi0( pi17 ), .pi1( pi18 ), .pi2( pi19 ), .pi3( pi49 ), .pi4( pi50 ), .pi5( pi51 ), .pi6( n4 ), .pi7( n5 ), .po0( tpo17 ), .po1( tpo18 ), .po2( tpo19 ), .po3( n6 ), .po4( n7 ) );
  adder32_8 U8 ( .pi00( pi20 ), .pi01( pi21 ), .pi02( pi22 ), .pi03( pi23 ), .pi04( pi52 ), .pi05( pi53 ), .pi06( pi54 ), .pi07( pi55 ), .pi08( n6 ), .pi09( n7 ), .po0( tpo20 ), .po1( tpo21 ), .po2( tpo22 ), .po3( tpo23 ), .po4( n8 ) );
endmodule
