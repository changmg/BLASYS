module mac(\a[0] , \a[1] , \a[2] , \a[3] , \b[0] , \b[1] , \b[2] , \b[3] , \c[0] , \c[1] , \c[2] , \c[3] , \r[0] , \r[1] , \r[2] , \r[3] , \r[4] , \r[5] , \r[6] , \r[7] );
  input \a[0] ;
  input \a[1] ;
  input \a[2] ;
  input \a[3] ;
  input \b[0] ;
  input \b[1] ;
  input \b[2] ;
  input \b[3] ;
  input \c[0] ;
  input \c[1] ;
  input \c[2] ;
  input \c[3] ;
  output \r[0] ;
  output \r[1] ;
  output \r[2] ;
  output \r[3] ;
  output \r[4] ;
  output \r[5] ;
  output \r[6] ;
  output \r[7] ;
  top U0 ( .pi00( \a[0] ) , .pi01( \a[1] ) , .pi02( \a[2] ) , .pi03( \a[3] ) , .pi04( \b[0] ) , .pi05( \b[1] ) , .pi06( \b[2] ) , .pi07( \b[3] ) , .pi08( \c[0] ) , .pi09( \c[1] ) , .pi10( \c[2] ) , .pi11( \c[3] ) , .po0( \r[0] ) , .po1( \r[1] ) , .po2( \r[2] ) , .po3( \r[3] ) , .po4( \r[4] ) , .po5( \r[5] ) , .po6( \r[6] ) , .po7( \r[7] ) );
endmodule

module top(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, po0, po1, po2, po3, po4, po5, po6, po7);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, tpo0, tpo1, tpo2, tpo3, tpo4, tpo5, tpo6, tpo7;
  assign po0 = tpo0;
  assign po1 = tpo1;
  assign po2 = tpo2;
  assign po3 = tpo3;
  assign po4 = tpo4;
  assign po5 = tpo5;
  assign po6 = tpo6;
  assign po7 = ~tpo7;
  mac_0 U0 ( .pi0( n3 ), .pi1( n4 ), .pi2( n7 ), .pi3( n8 ), .pi4( n9 ), .po0( tpo4 ), .po1( tpo5 ), .po2( n10 ) );
  mac_1 U1 ( .pi0( pi02 ), .pi1( pi03 ), .pi2( pi06 ), .pi3( pi07 ), .pi4( n0 ), .pi5( n5 ), .pi6( n6 ), .pi7( n10 ), .po0(  ), .po1(  ), .po2(  ), .po3(  ), .po4( n7 ), .po5( n9 ), .po6( tpo6 ), .po7( tpo7 ) );
  mac_2 U2 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi04 ), .pi3( pi05 ), .pi4( pi06 ), .pi5( pi08 ), .pi6( pi09 ), .pi7( n1 ), .pi8( n2 ), .po0( tpo0 ), .po1( tpo1 ), .po2( n0 ), .po3( tpo2 ), .po4( n3 ), .po5( tpo3 ), .po6( n4 ) );
  mac_3 U3 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi02 ), .pi3( pi03 ), .pi4( pi04 ), .pi5( pi05 ), .pi6( pi07 ), .pi7( pi10 ), .pi8( pi11 ), .po0(  ), .po1(  ), .po2(  ), .po3(  ), .po4( n1 ), .po5( n2 ), .po6( n5 ), .po7( n6 ), .po8( n8 ) );
endmodule
