module max_38_2(pi0 , pi1 , pi2 , pi3 , pi4 , po0 , po1 , po2 , po3 , po4 );
  input pi0 , pi1 , pi2 , pi3 , pi4 ;
  output po0 , po1 , po2 , po3 , po4 ;
  wire new_n6, new_n7, new_n8, new_n9, new_n10, new_n11, new_n12, new_n13, new_n14, new_n15, new_n16;
  assign new_n6 = pi0 & ~pi2 ;
  assign new_n7 = ~pi0 & pi2 ;
  assign new_n8 = ~pi1 & pi3 ;
  assign new_n9 = ~new_n7 & ~new_n8 ;
  assign new_n10 = pi1 & ~pi3 ;
  assign new_n11 = pi0 & pi4 ;
  assign new_n12 = pi2 & ~pi4 ;
  assign new_n13 = ~new_n11 & ~new_n12 ;
  assign new_n14 = pi1 & pi4 ;
  assign new_n15 = pi3 & ~pi4 ;
  assign new_n16 = ~new_n14 & ~new_n15 ;
  assign po0 = new_n6 ;
  assign po1 = new_n9 ;
  assign po2 = new_n10 ;
  assign po3 = new_n13 ;
  assign po4 = new_n16 ;
endmodule
