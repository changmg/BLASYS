module max_39(pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 , po0 , po1 , po2 , po3 , po4 , po5 );
  input pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 ;
  output po0 , po1 , po2 , po3 , po4 , po5 ;
  wire new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36, new_n37, new_n38, new_n39;
  assign new_n12 = pi02 & ~pi06 ;
  assign new_n13 = ~pi01 & pi05 ;
  assign new_n14 = ~pi00 & pi04 ;
  assign new_n15 = ~pi09 & ~new_n14 ;
  assign new_n16 = ~pi08 & new_n15 ;
  assign new_n17 = pi01 & ~pi05 ;
  assign new_n18 = pi00 & ~pi04 ;
  assign new_n19 = ~new_n17 & ~new_n18 ;
  assign new_n20 = ~new_n16 & new_n19 ;
  assign new_n21 = ~new_n13 & ~new_n20 ;
  assign new_n22 = ~new_n12 & ~new_n21 ;
  assign new_n23 = ~pi03 & pi07 ;
  assign new_n24 = ~pi02 & pi06 ;
  assign new_n25 = ~new_n23 & ~new_n24 ;
  assign new_n26 = ~new_n22 & new_n25 ;
  assign new_n27 = pi03 & ~pi07 ;
  assign new_n28 = pi00 & pi10 ;
  assign new_n29 = pi04 & ~pi10 ;
  assign new_n30 = ~new_n28 & ~new_n29 ;
  assign new_n31 = pi01 & pi10 ;
  assign new_n32 = pi05 & ~pi10 ;
  assign new_n33 = ~new_n31 & ~new_n32 ;
  assign new_n34 = pi02 & pi10 ;
  assign new_n35 = pi06 & ~pi10 ;
  assign new_n36 = ~new_n34 & ~new_n35 ;
  assign new_n37 = pi03 & pi10 ;
  assign new_n38 = pi07 & ~pi10 ;
  assign new_n39 = ~new_n37 & ~new_n38 ;
  assign po0 = new_n26 ;
  assign po1 = new_n27 ;
  assign po2 = new_n30 ;
  assign po3 = new_n33 ;
  assign po4 = new_n36 ;
  assign po5 = new_n39 ;
endmodule
