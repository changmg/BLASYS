module max_12_1(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , po0 , po1 , po2 , po3 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 ;
  output po0 , po1 , po2 , po3 ;
  wire new_n8, new_n9, new_n10, new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22;
  assign new_n8 = ~pi1 & pi3 ;
  assign new_n9 = ~pi0 & pi2 ;
  assign new_n10 = ~pi6 & ~new_n9 ;
  assign new_n11 = ~pi5 & new_n10 ;
  assign new_n12 = pi1 & ~pi3 ;
  assign new_n13 = pi0 & ~pi2 ;
  assign new_n14 = ~new_n12 & ~new_n13 ;
  assign new_n15 = ~new_n11 & new_n14 ;
  assign new_n16 = ~new_n8 & ~new_n15 ;
  assign new_n17 = pi0 & pi4 ;
  assign new_n18 = pi2 & ~pi4 ;
  assign new_n19 = ~new_n17 & ~new_n18 ;
  assign new_n20 = pi1 & pi4 ;
  assign new_n21 = pi3 & ~pi4 ;
  assign new_n22 = ~new_n20 & ~new_n21 ;
  assign po0 = pi4 ;
  assign po1 = new_n16 ;
  assign po2 = new_n19 ;
  assign po3 = new_n22 ;
endmodule
