module adder16(\in1[0] , \in1[1] , \in1[2] , \in1[3] , \in1[4] , \in1[5] , \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] , \in1[11] , \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in2[0] , \in2[1] , \in2[2] , \in2[3] , \in2[4] 
, \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] , \in2[10] , \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] , \res[0] , \res[1] , \res[2] , \res[3] , \res[4] , \res[5] , \res[6] , \res[7] , \res[8] , \res[9] 
, \res[10] , \res[11] , \res[12] , \res[13] , \res[14] , \res[15] , \res[16] );
  input \in1[0] ;
  input \in1[10] ;
  input \in1[11] ;
  input \in1[12] ;
  input \in1[13] ;
  input \in1[14] ;
  input \in1[15] ;
  input \in1[1] ;
  input \in1[2] ;
  input \in1[3] ;
  input \in1[4] ;
  input \in1[5] ;
  input \in1[6] ;
  input \in1[7] ;
  input \in1[8] ;
  input \in1[9] ;
  input \in2[0] ;
  input \in2[10] ;
  input \in2[11] ;
  input \in2[12] ;
  input \in2[13] ;
  input \in2[14] ;
  input \in2[15] ;
  input \in2[1] ;
  input \in2[2] ;
  input \in2[3] ;
  input \in2[4] ;
  input \in2[5] ;
  input \in2[6] ;
  input \in2[7] ;
  input \in2[8] ;
  input \in2[9] ;
  output \res[0] ;
  output \res[10] ;
  output \res[11] ;
  output \res[12] ;
  output \res[13] ;
  output \res[14] ;
  output \res[15] ;
  output \res[16] ;
  output \res[1] ;
  output \res[2] ;
  output \res[3] ;
  output \res[4] ;
  output \res[5] ;
  output \res[6] ;
  output \res[7] ;
  output \res[8] ;
  output \res[9] ;
  top U0 ( .pi00( \in1[0] ) , .pi01( \in1[1] ) , .pi02( \in1[2] ) , .pi03( \in1[3] ) , .pi04( \in1[4] ) , .pi05( \in1[5] ) , .pi06( \in1[6] ) , .pi07( \in1[7] ) , .pi08( \in1[8] ) , .pi09( \in1[9] ) , .pi10( \in1[10] ) , .pi11( \in1[11] ) , .pi12( \in1[12] ) , .pi13( \in1[13] ) , .pi14( \in1[14] ) , .pi15( \in1[15] ) , .pi16( \in2[0] ) , .pi17( \in2[1] ) , .pi18( \in2[2] ) , .pi19( \in2[3] ) , .pi20( \in2[4] ) , .pi21( \in2[5] ) , .pi22( \in2[6] ) , .pi23( \in2[7] ) , .pi24( \in2[8] ) , .pi25( \in2[9] ) , .pi26( \in2[10] ) , .pi27( \in2[11] ) , .pi28( \in2[12] ) , .pi29( \in2[13] ) , .pi30( \in2[14] ) , .pi31( \in2[15] ) , .po00( \res[0] ) , .po01( \res[1] ) , .po02( \res[2] ) , .po03( \res[3] ) , .po04( \res[4] ) , .po05( \res[5] ) , .po06( \res[6] ) , .po07( \res[7] ) , .po08( \res[8] ) , .po09( \res[9] ) , .po10( \res[10] ) , .po11( \res[11] ) , .po12( \res[12] ) , .po13( \res[13] ) , .po14( \res[14] ) , .po15( \res[15] ) , .po16( \res[16] ) );
endmodule

module top(pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16);
  input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16;
  wire n0, n1, n2, tpo00, tpo01, tpo02, tpo03, tpo04, tpo05, tpo06, tpo07, tpo08, tpo09, tpo10, tpo11, tpo12, tpo13, tpo14, tpo15, tpo16;
  assign po00 = tpo00;
  assign po01 = ~tpo01;
  assign po02 = tpo02;
  assign po03 = ~tpo03;
  assign po04 = tpo04;
  assign po05 = ~tpo05;
  assign po06 = ~tpo06;
  assign po07 = ~tpo07;
  assign po08 = tpo08;
  assign po09 = ~tpo09;
  assign po10 = tpo10;
  assign po11 = ~tpo11;
  assign po12 = tpo12;
  assign po13 = ~tpo13;
  assign po14 = ~tpo14;
  assign po15 = ~tpo15;
  assign po16 = ~tpo16;
  adder16_0 U0 ( .pi0( pi00 ), .pi1( pi01 ), .pi2( pi02 ), .pi3( pi16 ), .pi4( pi17 ), .pi5( pi18 ), .po0( tpo00 ), .po1( tpo01 ), .po2( tpo02 ), .po3( n0 ) );
  adder16_1 U1 ( .pi00( pi03 ), .pi01( pi04 ), .pi02( pi05 ), .pi03( pi06 ), .pi04( pi07 ), .pi05( pi19 ), .pi06( pi20 ), .pi07( pi21 ), .pi08( pi22 ), .pi09( pi23 ), .pi10( n0 ), .po0( tpo03 ), .po1( tpo04 ), .po2( tpo05 ), .po3( tpo06 ), .po4( tpo07 ), .po5( n1 ) );
  adder16_2 U2 ( .pi00( pi08 ), .pi01( pi09 ), .pi02( pi10 ), .pi03( pi11 ), .pi04( pi12 ), .pi05( pi24 ), .pi06( pi25 ), .pi07( pi26 ), .pi08( pi27 ), .pi09( pi28 ), .pi10( n1 ), .po0( tpo08 ), .po1( tpo09 ), .po2( tpo10 ), .po3( tpo11 ), .po4( tpo12 ), .po5( n2 ) );
  adder16_3 U3 ( .pi0( pi13 ), .pi1( pi14 ), .pi2( pi15 ), .pi3( pi29 ), .pi4( pi30 ), .pi5( pi31 ), .pi6( n2 ), .po0( tpo13 ), .po1( tpo14 ), .po2( tpo15 ), .po3( tpo16 ) );
endmodule
