module max_40_tb;
reg [12:0] pi;
wire [5:0] po;
max_40 dut(pi[12], pi[11], pi[10], pi[9], pi[8], pi[7], pi[6], pi[5], pi[4], pi[3], pi[2], pi[1], pi[0], po[5], po[4], po[3], po[2], po[1], po[0]);
initial
begin
# 1  pi=13'b0000000000000;
#1 $display("%b", po);
# 1  pi=13'b0000000000001;
#1 $display("%b", po);
# 1  pi=13'b0000000000010;
#1 $display("%b", po);
# 1  pi=13'b0000000000011;
#1 $display("%b", po);
# 1  pi=13'b0000000000100;
#1 $display("%b", po);
# 1  pi=13'b0000000000101;
#1 $display("%b", po);
# 1  pi=13'b0000000000110;
#1 $display("%b", po);
# 1  pi=13'b0000000000111;
#1 $display("%b", po);
# 1  pi=13'b0000000001000;
#1 $display("%b", po);
# 1  pi=13'b0000000001001;
#1 $display("%b", po);
# 1  pi=13'b0000000001010;
#1 $display("%b", po);
# 1  pi=13'b0000000001011;
#1 $display("%b", po);
# 1  pi=13'b0000000001100;
#1 $display("%b", po);
# 1  pi=13'b0000000001101;
#1 $display("%b", po);
# 1  pi=13'b0000000001110;
#1 $display("%b", po);
# 1  pi=13'b0000000001111;
#1 $display("%b", po);
# 1  pi=13'b0000000010000;
#1 $display("%b", po);
# 1  pi=13'b0000000010001;
#1 $display("%b", po);
# 1  pi=13'b0000000010010;
#1 $display("%b", po);
# 1  pi=13'b0000000010011;
#1 $display("%b", po);
# 1  pi=13'b0000000010100;
#1 $display("%b", po);
# 1  pi=13'b0000000010101;
#1 $display("%b", po);
# 1  pi=13'b0000000010110;
#1 $display("%b", po);
# 1  pi=13'b0000000010111;
#1 $display("%b", po);
# 1  pi=13'b0000000011000;
#1 $display("%b", po);
# 1  pi=13'b0000000011001;
#1 $display("%b", po);
# 1  pi=13'b0000000011010;
#1 $display("%b", po);
# 1  pi=13'b0000000011011;
#1 $display("%b", po);
# 1  pi=13'b0000000011100;
#1 $display("%b", po);
# 1  pi=13'b0000000011101;
#1 $display("%b", po);
# 1  pi=13'b0000000011110;
#1 $display("%b", po);
# 1  pi=13'b0000000011111;
#1 $display("%b", po);
# 1  pi=13'b0000000100000;
#1 $display("%b", po);
# 1  pi=13'b0000000100001;
#1 $display("%b", po);
# 1  pi=13'b0000000100010;
#1 $display("%b", po);
# 1  pi=13'b0000000100011;
#1 $display("%b", po);
# 1  pi=13'b0000000100100;
#1 $display("%b", po);
# 1  pi=13'b0000000100101;
#1 $display("%b", po);
# 1  pi=13'b0000000100110;
#1 $display("%b", po);
# 1  pi=13'b0000000100111;
#1 $display("%b", po);
# 1  pi=13'b0000000101000;
#1 $display("%b", po);
# 1  pi=13'b0000000101001;
#1 $display("%b", po);
# 1  pi=13'b0000000101010;
#1 $display("%b", po);
# 1  pi=13'b0000000101011;
#1 $display("%b", po);
# 1  pi=13'b0000000101100;
#1 $display("%b", po);
# 1  pi=13'b0000000101101;
#1 $display("%b", po);
# 1  pi=13'b0000000101110;
#1 $display("%b", po);
# 1  pi=13'b0000000101111;
#1 $display("%b", po);
# 1  pi=13'b0000000110000;
#1 $display("%b", po);
# 1  pi=13'b0000000110001;
#1 $display("%b", po);
# 1  pi=13'b0000000110010;
#1 $display("%b", po);
# 1  pi=13'b0000000110011;
#1 $display("%b", po);
# 1  pi=13'b0000000110100;
#1 $display("%b", po);
# 1  pi=13'b0000000110101;
#1 $display("%b", po);
# 1  pi=13'b0000000110110;
#1 $display("%b", po);
# 1  pi=13'b0000000110111;
#1 $display("%b", po);
# 1  pi=13'b0000000111000;
#1 $display("%b", po);
# 1  pi=13'b0000000111001;
#1 $display("%b", po);
# 1  pi=13'b0000000111010;
#1 $display("%b", po);
# 1  pi=13'b0000000111011;
#1 $display("%b", po);
# 1  pi=13'b0000000111100;
#1 $display("%b", po);
# 1  pi=13'b0000000111101;
#1 $display("%b", po);
# 1  pi=13'b0000000111110;
#1 $display("%b", po);
# 1  pi=13'b0000000111111;
#1 $display("%b", po);
# 1  pi=13'b0000001000000;
#1 $display("%b", po);
# 1  pi=13'b0000001000001;
#1 $display("%b", po);
# 1  pi=13'b0000001000010;
#1 $display("%b", po);
# 1  pi=13'b0000001000011;
#1 $display("%b", po);
# 1  pi=13'b0000001000100;
#1 $display("%b", po);
# 1  pi=13'b0000001000101;
#1 $display("%b", po);
# 1  pi=13'b0000001000110;
#1 $display("%b", po);
# 1  pi=13'b0000001000111;
#1 $display("%b", po);
# 1  pi=13'b0000001001000;
#1 $display("%b", po);
# 1  pi=13'b0000001001001;
#1 $display("%b", po);
# 1  pi=13'b0000001001010;
#1 $display("%b", po);
# 1  pi=13'b0000001001011;
#1 $display("%b", po);
# 1  pi=13'b0000001001100;
#1 $display("%b", po);
# 1  pi=13'b0000001001101;
#1 $display("%b", po);
# 1  pi=13'b0000001001110;
#1 $display("%b", po);
# 1  pi=13'b0000001001111;
#1 $display("%b", po);
# 1  pi=13'b0000001010000;
#1 $display("%b", po);
# 1  pi=13'b0000001010001;
#1 $display("%b", po);
# 1  pi=13'b0000001010010;
#1 $display("%b", po);
# 1  pi=13'b0000001010011;
#1 $display("%b", po);
# 1  pi=13'b0000001010100;
#1 $display("%b", po);
# 1  pi=13'b0000001010101;
#1 $display("%b", po);
# 1  pi=13'b0000001010110;
#1 $display("%b", po);
# 1  pi=13'b0000001010111;
#1 $display("%b", po);
# 1  pi=13'b0000001011000;
#1 $display("%b", po);
# 1  pi=13'b0000001011001;
#1 $display("%b", po);
# 1  pi=13'b0000001011010;
#1 $display("%b", po);
# 1  pi=13'b0000001011011;
#1 $display("%b", po);
# 1  pi=13'b0000001011100;
#1 $display("%b", po);
# 1  pi=13'b0000001011101;
#1 $display("%b", po);
# 1  pi=13'b0000001011110;
#1 $display("%b", po);
# 1  pi=13'b0000001011111;
#1 $display("%b", po);
# 1  pi=13'b0000001100000;
#1 $display("%b", po);
# 1  pi=13'b0000001100001;
#1 $display("%b", po);
# 1  pi=13'b0000001100010;
#1 $display("%b", po);
# 1  pi=13'b0000001100011;
#1 $display("%b", po);
# 1  pi=13'b0000001100100;
#1 $display("%b", po);
# 1  pi=13'b0000001100101;
#1 $display("%b", po);
# 1  pi=13'b0000001100110;
#1 $display("%b", po);
# 1  pi=13'b0000001100111;
#1 $display("%b", po);
# 1  pi=13'b0000001101000;
#1 $display("%b", po);
# 1  pi=13'b0000001101001;
#1 $display("%b", po);
# 1  pi=13'b0000001101010;
#1 $display("%b", po);
# 1  pi=13'b0000001101011;
#1 $display("%b", po);
# 1  pi=13'b0000001101100;
#1 $display("%b", po);
# 1  pi=13'b0000001101101;
#1 $display("%b", po);
# 1  pi=13'b0000001101110;
#1 $display("%b", po);
# 1  pi=13'b0000001101111;
#1 $display("%b", po);
# 1  pi=13'b0000001110000;
#1 $display("%b", po);
# 1  pi=13'b0000001110001;
#1 $display("%b", po);
# 1  pi=13'b0000001110010;
#1 $display("%b", po);
# 1  pi=13'b0000001110011;
#1 $display("%b", po);
# 1  pi=13'b0000001110100;
#1 $display("%b", po);
# 1  pi=13'b0000001110101;
#1 $display("%b", po);
# 1  pi=13'b0000001110110;
#1 $display("%b", po);
# 1  pi=13'b0000001110111;
#1 $display("%b", po);
# 1  pi=13'b0000001111000;
#1 $display("%b", po);
# 1  pi=13'b0000001111001;
#1 $display("%b", po);
# 1  pi=13'b0000001111010;
#1 $display("%b", po);
# 1  pi=13'b0000001111011;
#1 $display("%b", po);
# 1  pi=13'b0000001111100;
#1 $display("%b", po);
# 1  pi=13'b0000001111101;
#1 $display("%b", po);
# 1  pi=13'b0000001111110;
#1 $display("%b", po);
# 1  pi=13'b0000001111111;
#1 $display("%b", po);
# 1  pi=13'b0000010000000;
#1 $display("%b", po);
# 1  pi=13'b0000010000001;
#1 $display("%b", po);
# 1  pi=13'b0000010000010;
#1 $display("%b", po);
# 1  pi=13'b0000010000011;
#1 $display("%b", po);
# 1  pi=13'b0000010000100;
#1 $display("%b", po);
# 1  pi=13'b0000010000101;
#1 $display("%b", po);
# 1  pi=13'b0000010000110;
#1 $display("%b", po);
# 1  pi=13'b0000010000111;
#1 $display("%b", po);
# 1  pi=13'b0000010001000;
#1 $display("%b", po);
# 1  pi=13'b0000010001001;
#1 $display("%b", po);
# 1  pi=13'b0000010001010;
#1 $display("%b", po);
# 1  pi=13'b0000010001011;
#1 $display("%b", po);
# 1  pi=13'b0000010001100;
#1 $display("%b", po);
# 1  pi=13'b0000010001101;
#1 $display("%b", po);
# 1  pi=13'b0000010001110;
#1 $display("%b", po);
# 1  pi=13'b0000010001111;
#1 $display("%b", po);
# 1  pi=13'b0000010010000;
#1 $display("%b", po);
# 1  pi=13'b0000010010001;
#1 $display("%b", po);
# 1  pi=13'b0000010010010;
#1 $display("%b", po);
# 1  pi=13'b0000010010011;
#1 $display("%b", po);
# 1  pi=13'b0000010010100;
#1 $display("%b", po);
# 1  pi=13'b0000010010101;
#1 $display("%b", po);
# 1  pi=13'b0000010010110;
#1 $display("%b", po);
# 1  pi=13'b0000010010111;
#1 $display("%b", po);
# 1  pi=13'b0000010011000;
#1 $display("%b", po);
# 1  pi=13'b0000010011001;
#1 $display("%b", po);
# 1  pi=13'b0000010011010;
#1 $display("%b", po);
# 1  pi=13'b0000010011011;
#1 $display("%b", po);
# 1  pi=13'b0000010011100;
#1 $display("%b", po);
# 1  pi=13'b0000010011101;
#1 $display("%b", po);
# 1  pi=13'b0000010011110;
#1 $display("%b", po);
# 1  pi=13'b0000010011111;
#1 $display("%b", po);
# 1  pi=13'b0000010100000;
#1 $display("%b", po);
# 1  pi=13'b0000010100001;
#1 $display("%b", po);
# 1  pi=13'b0000010100010;
#1 $display("%b", po);
# 1  pi=13'b0000010100011;
#1 $display("%b", po);
# 1  pi=13'b0000010100100;
#1 $display("%b", po);
# 1  pi=13'b0000010100101;
#1 $display("%b", po);
# 1  pi=13'b0000010100110;
#1 $display("%b", po);
# 1  pi=13'b0000010100111;
#1 $display("%b", po);
# 1  pi=13'b0000010101000;
#1 $display("%b", po);
# 1  pi=13'b0000010101001;
#1 $display("%b", po);
# 1  pi=13'b0000010101010;
#1 $display("%b", po);
# 1  pi=13'b0000010101011;
#1 $display("%b", po);
# 1  pi=13'b0000010101100;
#1 $display("%b", po);
# 1  pi=13'b0000010101101;
#1 $display("%b", po);
# 1  pi=13'b0000010101110;
#1 $display("%b", po);
# 1  pi=13'b0000010101111;
#1 $display("%b", po);
# 1  pi=13'b0000010110000;
#1 $display("%b", po);
# 1  pi=13'b0000010110001;
#1 $display("%b", po);
# 1  pi=13'b0000010110010;
#1 $display("%b", po);
# 1  pi=13'b0000010110011;
#1 $display("%b", po);
# 1  pi=13'b0000010110100;
#1 $display("%b", po);
# 1  pi=13'b0000010110101;
#1 $display("%b", po);
# 1  pi=13'b0000010110110;
#1 $display("%b", po);
# 1  pi=13'b0000010110111;
#1 $display("%b", po);
# 1  pi=13'b0000010111000;
#1 $display("%b", po);
# 1  pi=13'b0000010111001;
#1 $display("%b", po);
# 1  pi=13'b0000010111010;
#1 $display("%b", po);
# 1  pi=13'b0000010111011;
#1 $display("%b", po);
# 1  pi=13'b0000010111100;
#1 $display("%b", po);
# 1  pi=13'b0000010111101;
#1 $display("%b", po);
# 1  pi=13'b0000010111110;
#1 $display("%b", po);
# 1  pi=13'b0000010111111;
#1 $display("%b", po);
# 1  pi=13'b0000011000000;
#1 $display("%b", po);
# 1  pi=13'b0000011000001;
#1 $display("%b", po);
# 1  pi=13'b0000011000010;
#1 $display("%b", po);
# 1  pi=13'b0000011000011;
#1 $display("%b", po);
# 1  pi=13'b0000011000100;
#1 $display("%b", po);
# 1  pi=13'b0000011000101;
#1 $display("%b", po);
# 1  pi=13'b0000011000110;
#1 $display("%b", po);
# 1  pi=13'b0000011000111;
#1 $display("%b", po);
# 1  pi=13'b0000011001000;
#1 $display("%b", po);
# 1  pi=13'b0000011001001;
#1 $display("%b", po);
# 1  pi=13'b0000011001010;
#1 $display("%b", po);
# 1  pi=13'b0000011001011;
#1 $display("%b", po);
# 1  pi=13'b0000011001100;
#1 $display("%b", po);
# 1  pi=13'b0000011001101;
#1 $display("%b", po);
# 1  pi=13'b0000011001110;
#1 $display("%b", po);
# 1  pi=13'b0000011001111;
#1 $display("%b", po);
# 1  pi=13'b0000011010000;
#1 $display("%b", po);
# 1  pi=13'b0000011010001;
#1 $display("%b", po);
# 1  pi=13'b0000011010010;
#1 $display("%b", po);
# 1  pi=13'b0000011010011;
#1 $display("%b", po);
# 1  pi=13'b0000011010100;
#1 $display("%b", po);
# 1  pi=13'b0000011010101;
#1 $display("%b", po);
# 1  pi=13'b0000011010110;
#1 $display("%b", po);
# 1  pi=13'b0000011010111;
#1 $display("%b", po);
# 1  pi=13'b0000011011000;
#1 $display("%b", po);
# 1  pi=13'b0000011011001;
#1 $display("%b", po);
# 1  pi=13'b0000011011010;
#1 $display("%b", po);
# 1  pi=13'b0000011011011;
#1 $display("%b", po);
# 1  pi=13'b0000011011100;
#1 $display("%b", po);
# 1  pi=13'b0000011011101;
#1 $display("%b", po);
# 1  pi=13'b0000011011110;
#1 $display("%b", po);
# 1  pi=13'b0000011011111;
#1 $display("%b", po);
# 1  pi=13'b0000011100000;
#1 $display("%b", po);
# 1  pi=13'b0000011100001;
#1 $display("%b", po);
# 1  pi=13'b0000011100010;
#1 $display("%b", po);
# 1  pi=13'b0000011100011;
#1 $display("%b", po);
# 1  pi=13'b0000011100100;
#1 $display("%b", po);
# 1  pi=13'b0000011100101;
#1 $display("%b", po);
# 1  pi=13'b0000011100110;
#1 $display("%b", po);
# 1  pi=13'b0000011100111;
#1 $display("%b", po);
# 1  pi=13'b0000011101000;
#1 $display("%b", po);
# 1  pi=13'b0000011101001;
#1 $display("%b", po);
# 1  pi=13'b0000011101010;
#1 $display("%b", po);
# 1  pi=13'b0000011101011;
#1 $display("%b", po);
# 1  pi=13'b0000011101100;
#1 $display("%b", po);
# 1  pi=13'b0000011101101;
#1 $display("%b", po);
# 1  pi=13'b0000011101110;
#1 $display("%b", po);
# 1  pi=13'b0000011101111;
#1 $display("%b", po);
# 1  pi=13'b0000011110000;
#1 $display("%b", po);
# 1  pi=13'b0000011110001;
#1 $display("%b", po);
# 1  pi=13'b0000011110010;
#1 $display("%b", po);
# 1  pi=13'b0000011110011;
#1 $display("%b", po);
# 1  pi=13'b0000011110100;
#1 $display("%b", po);
# 1  pi=13'b0000011110101;
#1 $display("%b", po);
# 1  pi=13'b0000011110110;
#1 $display("%b", po);
# 1  pi=13'b0000011110111;
#1 $display("%b", po);
# 1  pi=13'b0000011111000;
#1 $display("%b", po);
# 1  pi=13'b0000011111001;
#1 $display("%b", po);
# 1  pi=13'b0000011111010;
#1 $display("%b", po);
# 1  pi=13'b0000011111011;
#1 $display("%b", po);
# 1  pi=13'b0000011111100;
#1 $display("%b", po);
# 1  pi=13'b0000011111101;
#1 $display("%b", po);
# 1  pi=13'b0000011111110;
#1 $display("%b", po);
# 1  pi=13'b0000011111111;
#1 $display("%b", po);
# 1  pi=13'b0000100000000;
#1 $display("%b", po);
# 1  pi=13'b0000100000001;
#1 $display("%b", po);
# 1  pi=13'b0000100000010;
#1 $display("%b", po);
# 1  pi=13'b0000100000011;
#1 $display("%b", po);
# 1  pi=13'b0000100000100;
#1 $display("%b", po);
# 1  pi=13'b0000100000101;
#1 $display("%b", po);
# 1  pi=13'b0000100000110;
#1 $display("%b", po);
# 1  pi=13'b0000100000111;
#1 $display("%b", po);
# 1  pi=13'b0000100001000;
#1 $display("%b", po);
# 1  pi=13'b0000100001001;
#1 $display("%b", po);
# 1  pi=13'b0000100001010;
#1 $display("%b", po);
# 1  pi=13'b0000100001011;
#1 $display("%b", po);
# 1  pi=13'b0000100001100;
#1 $display("%b", po);
# 1  pi=13'b0000100001101;
#1 $display("%b", po);
# 1  pi=13'b0000100001110;
#1 $display("%b", po);
# 1  pi=13'b0000100001111;
#1 $display("%b", po);
# 1  pi=13'b0000100010000;
#1 $display("%b", po);
# 1  pi=13'b0000100010001;
#1 $display("%b", po);
# 1  pi=13'b0000100010010;
#1 $display("%b", po);
# 1  pi=13'b0000100010011;
#1 $display("%b", po);
# 1  pi=13'b0000100010100;
#1 $display("%b", po);
# 1  pi=13'b0000100010101;
#1 $display("%b", po);
# 1  pi=13'b0000100010110;
#1 $display("%b", po);
# 1  pi=13'b0000100010111;
#1 $display("%b", po);
# 1  pi=13'b0000100011000;
#1 $display("%b", po);
# 1  pi=13'b0000100011001;
#1 $display("%b", po);
# 1  pi=13'b0000100011010;
#1 $display("%b", po);
# 1  pi=13'b0000100011011;
#1 $display("%b", po);
# 1  pi=13'b0000100011100;
#1 $display("%b", po);
# 1  pi=13'b0000100011101;
#1 $display("%b", po);
# 1  pi=13'b0000100011110;
#1 $display("%b", po);
# 1  pi=13'b0000100011111;
#1 $display("%b", po);
# 1  pi=13'b0000100100000;
#1 $display("%b", po);
# 1  pi=13'b0000100100001;
#1 $display("%b", po);
# 1  pi=13'b0000100100010;
#1 $display("%b", po);
# 1  pi=13'b0000100100011;
#1 $display("%b", po);
# 1  pi=13'b0000100100100;
#1 $display("%b", po);
# 1  pi=13'b0000100100101;
#1 $display("%b", po);
# 1  pi=13'b0000100100110;
#1 $display("%b", po);
# 1  pi=13'b0000100100111;
#1 $display("%b", po);
# 1  pi=13'b0000100101000;
#1 $display("%b", po);
# 1  pi=13'b0000100101001;
#1 $display("%b", po);
# 1  pi=13'b0000100101010;
#1 $display("%b", po);
# 1  pi=13'b0000100101011;
#1 $display("%b", po);
# 1  pi=13'b0000100101100;
#1 $display("%b", po);
# 1  pi=13'b0000100101101;
#1 $display("%b", po);
# 1  pi=13'b0000100101110;
#1 $display("%b", po);
# 1  pi=13'b0000100101111;
#1 $display("%b", po);
# 1  pi=13'b0000100110000;
#1 $display("%b", po);
# 1  pi=13'b0000100110001;
#1 $display("%b", po);
# 1  pi=13'b0000100110010;
#1 $display("%b", po);
# 1  pi=13'b0000100110011;
#1 $display("%b", po);
# 1  pi=13'b0000100110100;
#1 $display("%b", po);
# 1  pi=13'b0000100110101;
#1 $display("%b", po);
# 1  pi=13'b0000100110110;
#1 $display("%b", po);
# 1  pi=13'b0000100110111;
#1 $display("%b", po);
# 1  pi=13'b0000100111000;
#1 $display("%b", po);
# 1  pi=13'b0000100111001;
#1 $display("%b", po);
# 1  pi=13'b0000100111010;
#1 $display("%b", po);
# 1  pi=13'b0000100111011;
#1 $display("%b", po);
# 1  pi=13'b0000100111100;
#1 $display("%b", po);
# 1  pi=13'b0000100111101;
#1 $display("%b", po);
# 1  pi=13'b0000100111110;
#1 $display("%b", po);
# 1  pi=13'b0000100111111;
#1 $display("%b", po);
# 1  pi=13'b0000101000000;
#1 $display("%b", po);
# 1  pi=13'b0000101000001;
#1 $display("%b", po);
# 1  pi=13'b0000101000010;
#1 $display("%b", po);
# 1  pi=13'b0000101000011;
#1 $display("%b", po);
# 1  pi=13'b0000101000100;
#1 $display("%b", po);
# 1  pi=13'b0000101000101;
#1 $display("%b", po);
# 1  pi=13'b0000101000110;
#1 $display("%b", po);
# 1  pi=13'b0000101000111;
#1 $display("%b", po);
# 1  pi=13'b0000101001000;
#1 $display("%b", po);
# 1  pi=13'b0000101001001;
#1 $display("%b", po);
# 1  pi=13'b0000101001010;
#1 $display("%b", po);
# 1  pi=13'b0000101001011;
#1 $display("%b", po);
# 1  pi=13'b0000101001100;
#1 $display("%b", po);
# 1  pi=13'b0000101001101;
#1 $display("%b", po);
# 1  pi=13'b0000101001110;
#1 $display("%b", po);
# 1  pi=13'b0000101001111;
#1 $display("%b", po);
# 1  pi=13'b0000101010000;
#1 $display("%b", po);
# 1  pi=13'b0000101010001;
#1 $display("%b", po);
# 1  pi=13'b0000101010010;
#1 $display("%b", po);
# 1  pi=13'b0000101010011;
#1 $display("%b", po);
# 1  pi=13'b0000101010100;
#1 $display("%b", po);
# 1  pi=13'b0000101010101;
#1 $display("%b", po);
# 1  pi=13'b0000101010110;
#1 $display("%b", po);
# 1  pi=13'b0000101010111;
#1 $display("%b", po);
# 1  pi=13'b0000101011000;
#1 $display("%b", po);
# 1  pi=13'b0000101011001;
#1 $display("%b", po);
# 1  pi=13'b0000101011010;
#1 $display("%b", po);
# 1  pi=13'b0000101011011;
#1 $display("%b", po);
# 1  pi=13'b0000101011100;
#1 $display("%b", po);
# 1  pi=13'b0000101011101;
#1 $display("%b", po);
# 1  pi=13'b0000101011110;
#1 $display("%b", po);
# 1  pi=13'b0000101011111;
#1 $display("%b", po);
# 1  pi=13'b0000101100000;
#1 $display("%b", po);
# 1  pi=13'b0000101100001;
#1 $display("%b", po);
# 1  pi=13'b0000101100010;
#1 $display("%b", po);
# 1  pi=13'b0000101100011;
#1 $display("%b", po);
# 1  pi=13'b0000101100100;
#1 $display("%b", po);
# 1  pi=13'b0000101100101;
#1 $display("%b", po);
# 1  pi=13'b0000101100110;
#1 $display("%b", po);
# 1  pi=13'b0000101100111;
#1 $display("%b", po);
# 1  pi=13'b0000101101000;
#1 $display("%b", po);
# 1  pi=13'b0000101101001;
#1 $display("%b", po);
# 1  pi=13'b0000101101010;
#1 $display("%b", po);
# 1  pi=13'b0000101101011;
#1 $display("%b", po);
# 1  pi=13'b0000101101100;
#1 $display("%b", po);
# 1  pi=13'b0000101101101;
#1 $display("%b", po);
# 1  pi=13'b0000101101110;
#1 $display("%b", po);
# 1  pi=13'b0000101101111;
#1 $display("%b", po);
# 1  pi=13'b0000101110000;
#1 $display("%b", po);
# 1  pi=13'b0000101110001;
#1 $display("%b", po);
# 1  pi=13'b0000101110010;
#1 $display("%b", po);
# 1  pi=13'b0000101110011;
#1 $display("%b", po);
# 1  pi=13'b0000101110100;
#1 $display("%b", po);
# 1  pi=13'b0000101110101;
#1 $display("%b", po);
# 1  pi=13'b0000101110110;
#1 $display("%b", po);
# 1  pi=13'b0000101110111;
#1 $display("%b", po);
# 1  pi=13'b0000101111000;
#1 $display("%b", po);
# 1  pi=13'b0000101111001;
#1 $display("%b", po);
# 1  pi=13'b0000101111010;
#1 $display("%b", po);
# 1  pi=13'b0000101111011;
#1 $display("%b", po);
# 1  pi=13'b0000101111100;
#1 $display("%b", po);
# 1  pi=13'b0000101111101;
#1 $display("%b", po);
# 1  pi=13'b0000101111110;
#1 $display("%b", po);
# 1  pi=13'b0000101111111;
#1 $display("%b", po);
# 1  pi=13'b0000110000000;
#1 $display("%b", po);
# 1  pi=13'b0000110000001;
#1 $display("%b", po);
# 1  pi=13'b0000110000010;
#1 $display("%b", po);
# 1  pi=13'b0000110000011;
#1 $display("%b", po);
# 1  pi=13'b0000110000100;
#1 $display("%b", po);
# 1  pi=13'b0000110000101;
#1 $display("%b", po);
# 1  pi=13'b0000110000110;
#1 $display("%b", po);
# 1  pi=13'b0000110000111;
#1 $display("%b", po);
# 1  pi=13'b0000110001000;
#1 $display("%b", po);
# 1  pi=13'b0000110001001;
#1 $display("%b", po);
# 1  pi=13'b0000110001010;
#1 $display("%b", po);
# 1  pi=13'b0000110001011;
#1 $display("%b", po);
# 1  pi=13'b0000110001100;
#1 $display("%b", po);
# 1  pi=13'b0000110001101;
#1 $display("%b", po);
# 1  pi=13'b0000110001110;
#1 $display("%b", po);
# 1  pi=13'b0000110001111;
#1 $display("%b", po);
# 1  pi=13'b0000110010000;
#1 $display("%b", po);
# 1  pi=13'b0000110010001;
#1 $display("%b", po);
# 1  pi=13'b0000110010010;
#1 $display("%b", po);
# 1  pi=13'b0000110010011;
#1 $display("%b", po);
# 1  pi=13'b0000110010100;
#1 $display("%b", po);
# 1  pi=13'b0000110010101;
#1 $display("%b", po);
# 1  pi=13'b0000110010110;
#1 $display("%b", po);
# 1  pi=13'b0000110010111;
#1 $display("%b", po);
# 1  pi=13'b0000110011000;
#1 $display("%b", po);
# 1  pi=13'b0000110011001;
#1 $display("%b", po);
# 1  pi=13'b0000110011010;
#1 $display("%b", po);
# 1  pi=13'b0000110011011;
#1 $display("%b", po);
# 1  pi=13'b0000110011100;
#1 $display("%b", po);
# 1  pi=13'b0000110011101;
#1 $display("%b", po);
# 1  pi=13'b0000110011110;
#1 $display("%b", po);
# 1  pi=13'b0000110011111;
#1 $display("%b", po);
# 1  pi=13'b0000110100000;
#1 $display("%b", po);
# 1  pi=13'b0000110100001;
#1 $display("%b", po);
# 1  pi=13'b0000110100010;
#1 $display("%b", po);
# 1  pi=13'b0000110100011;
#1 $display("%b", po);
# 1  pi=13'b0000110100100;
#1 $display("%b", po);
# 1  pi=13'b0000110100101;
#1 $display("%b", po);
# 1  pi=13'b0000110100110;
#1 $display("%b", po);
# 1  pi=13'b0000110100111;
#1 $display("%b", po);
# 1  pi=13'b0000110101000;
#1 $display("%b", po);
# 1  pi=13'b0000110101001;
#1 $display("%b", po);
# 1  pi=13'b0000110101010;
#1 $display("%b", po);
# 1  pi=13'b0000110101011;
#1 $display("%b", po);
# 1  pi=13'b0000110101100;
#1 $display("%b", po);
# 1  pi=13'b0000110101101;
#1 $display("%b", po);
# 1  pi=13'b0000110101110;
#1 $display("%b", po);
# 1  pi=13'b0000110101111;
#1 $display("%b", po);
# 1  pi=13'b0000110110000;
#1 $display("%b", po);
# 1  pi=13'b0000110110001;
#1 $display("%b", po);
# 1  pi=13'b0000110110010;
#1 $display("%b", po);
# 1  pi=13'b0000110110011;
#1 $display("%b", po);
# 1  pi=13'b0000110110100;
#1 $display("%b", po);
# 1  pi=13'b0000110110101;
#1 $display("%b", po);
# 1  pi=13'b0000110110110;
#1 $display("%b", po);
# 1  pi=13'b0000110110111;
#1 $display("%b", po);
# 1  pi=13'b0000110111000;
#1 $display("%b", po);
# 1  pi=13'b0000110111001;
#1 $display("%b", po);
# 1  pi=13'b0000110111010;
#1 $display("%b", po);
# 1  pi=13'b0000110111011;
#1 $display("%b", po);
# 1  pi=13'b0000110111100;
#1 $display("%b", po);
# 1  pi=13'b0000110111101;
#1 $display("%b", po);
# 1  pi=13'b0000110111110;
#1 $display("%b", po);
# 1  pi=13'b0000110111111;
#1 $display("%b", po);
# 1  pi=13'b0000111000000;
#1 $display("%b", po);
# 1  pi=13'b0000111000001;
#1 $display("%b", po);
# 1  pi=13'b0000111000010;
#1 $display("%b", po);
# 1  pi=13'b0000111000011;
#1 $display("%b", po);
# 1  pi=13'b0000111000100;
#1 $display("%b", po);
# 1  pi=13'b0000111000101;
#1 $display("%b", po);
# 1  pi=13'b0000111000110;
#1 $display("%b", po);
# 1  pi=13'b0000111000111;
#1 $display("%b", po);
# 1  pi=13'b0000111001000;
#1 $display("%b", po);
# 1  pi=13'b0000111001001;
#1 $display("%b", po);
# 1  pi=13'b0000111001010;
#1 $display("%b", po);
# 1  pi=13'b0000111001011;
#1 $display("%b", po);
# 1  pi=13'b0000111001100;
#1 $display("%b", po);
# 1  pi=13'b0000111001101;
#1 $display("%b", po);
# 1  pi=13'b0000111001110;
#1 $display("%b", po);
# 1  pi=13'b0000111001111;
#1 $display("%b", po);
# 1  pi=13'b0000111010000;
#1 $display("%b", po);
# 1  pi=13'b0000111010001;
#1 $display("%b", po);
# 1  pi=13'b0000111010010;
#1 $display("%b", po);
# 1  pi=13'b0000111010011;
#1 $display("%b", po);
# 1  pi=13'b0000111010100;
#1 $display("%b", po);
# 1  pi=13'b0000111010101;
#1 $display("%b", po);
# 1  pi=13'b0000111010110;
#1 $display("%b", po);
# 1  pi=13'b0000111010111;
#1 $display("%b", po);
# 1  pi=13'b0000111011000;
#1 $display("%b", po);
# 1  pi=13'b0000111011001;
#1 $display("%b", po);
# 1  pi=13'b0000111011010;
#1 $display("%b", po);
# 1  pi=13'b0000111011011;
#1 $display("%b", po);
# 1  pi=13'b0000111011100;
#1 $display("%b", po);
# 1  pi=13'b0000111011101;
#1 $display("%b", po);
# 1  pi=13'b0000111011110;
#1 $display("%b", po);
# 1  pi=13'b0000111011111;
#1 $display("%b", po);
# 1  pi=13'b0000111100000;
#1 $display("%b", po);
# 1  pi=13'b0000111100001;
#1 $display("%b", po);
# 1  pi=13'b0000111100010;
#1 $display("%b", po);
# 1  pi=13'b0000111100011;
#1 $display("%b", po);
# 1  pi=13'b0000111100100;
#1 $display("%b", po);
# 1  pi=13'b0000111100101;
#1 $display("%b", po);
# 1  pi=13'b0000111100110;
#1 $display("%b", po);
# 1  pi=13'b0000111100111;
#1 $display("%b", po);
# 1  pi=13'b0000111101000;
#1 $display("%b", po);
# 1  pi=13'b0000111101001;
#1 $display("%b", po);
# 1  pi=13'b0000111101010;
#1 $display("%b", po);
# 1  pi=13'b0000111101011;
#1 $display("%b", po);
# 1  pi=13'b0000111101100;
#1 $display("%b", po);
# 1  pi=13'b0000111101101;
#1 $display("%b", po);
# 1  pi=13'b0000111101110;
#1 $display("%b", po);
# 1  pi=13'b0000111101111;
#1 $display("%b", po);
# 1  pi=13'b0000111110000;
#1 $display("%b", po);
# 1  pi=13'b0000111110001;
#1 $display("%b", po);
# 1  pi=13'b0000111110010;
#1 $display("%b", po);
# 1  pi=13'b0000111110011;
#1 $display("%b", po);
# 1  pi=13'b0000111110100;
#1 $display("%b", po);
# 1  pi=13'b0000111110101;
#1 $display("%b", po);
# 1  pi=13'b0000111110110;
#1 $display("%b", po);
# 1  pi=13'b0000111110111;
#1 $display("%b", po);
# 1  pi=13'b0000111111000;
#1 $display("%b", po);
# 1  pi=13'b0000111111001;
#1 $display("%b", po);
# 1  pi=13'b0000111111010;
#1 $display("%b", po);
# 1  pi=13'b0000111111011;
#1 $display("%b", po);
# 1  pi=13'b0000111111100;
#1 $display("%b", po);
# 1  pi=13'b0000111111101;
#1 $display("%b", po);
# 1  pi=13'b0000111111110;
#1 $display("%b", po);
# 1  pi=13'b0000111111111;
#1 $display("%b", po);
# 1  pi=13'b0001000000000;
#1 $display("%b", po);
# 1  pi=13'b0001000000001;
#1 $display("%b", po);
# 1  pi=13'b0001000000010;
#1 $display("%b", po);
# 1  pi=13'b0001000000011;
#1 $display("%b", po);
# 1  pi=13'b0001000000100;
#1 $display("%b", po);
# 1  pi=13'b0001000000101;
#1 $display("%b", po);
# 1  pi=13'b0001000000110;
#1 $display("%b", po);
# 1  pi=13'b0001000000111;
#1 $display("%b", po);
# 1  pi=13'b0001000001000;
#1 $display("%b", po);
# 1  pi=13'b0001000001001;
#1 $display("%b", po);
# 1  pi=13'b0001000001010;
#1 $display("%b", po);
# 1  pi=13'b0001000001011;
#1 $display("%b", po);
# 1  pi=13'b0001000001100;
#1 $display("%b", po);
# 1  pi=13'b0001000001101;
#1 $display("%b", po);
# 1  pi=13'b0001000001110;
#1 $display("%b", po);
# 1  pi=13'b0001000001111;
#1 $display("%b", po);
# 1  pi=13'b0001000010000;
#1 $display("%b", po);
# 1  pi=13'b0001000010001;
#1 $display("%b", po);
# 1  pi=13'b0001000010010;
#1 $display("%b", po);
# 1  pi=13'b0001000010011;
#1 $display("%b", po);
# 1  pi=13'b0001000010100;
#1 $display("%b", po);
# 1  pi=13'b0001000010101;
#1 $display("%b", po);
# 1  pi=13'b0001000010110;
#1 $display("%b", po);
# 1  pi=13'b0001000010111;
#1 $display("%b", po);
# 1  pi=13'b0001000011000;
#1 $display("%b", po);
# 1  pi=13'b0001000011001;
#1 $display("%b", po);
# 1  pi=13'b0001000011010;
#1 $display("%b", po);
# 1  pi=13'b0001000011011;
#1 $display("%b", po);
# 1  pi=13'b0001000011100;
#1 $display("%b", po);
# 1  pi=13'b0001000011101;
#1 $display("%b", po);
# 1  pi=13'b0001000011110;
#1 $display("%b", po);
# 1  pi=13'b0001000011111;
#1 $display("%b", po);
# 1  pi=13'b0001000100000;
#1 $display("%b", po);
# 1  pi=13'b0001000100001;
#1 $display("%b", po);
# 1  pi=13'b0001000100010;
#1 $display("%b", po);
# 1  pi=13'b0001000100011;
#1 $display("%b", po);
# 1  pi=13'b0001000100100;
#1 $display("%b", po);
# 1  pi=13'b0001000100101;
#1 $display("%b", po);
# 1  pi=13'b0001000100110;
#1 $display("%b", po);
# 1  pi=13'b0001000100111;
#1 $display("%b", po);
# 1  pi=13'b0001000101000;
#1 $display("%b", po);
# 1  pi=13'b0001000101001;
#1 $display("%b", po);
# 1  pi=13'b0001000101010;
#1 $display("%b", po);
# 1  pi=13'b0001000101011;
#1 $display("%b", po);
# 1  pi=13'b0001000101100;
#1 $display("%b", po);
# 1  pi=13'b0001000101101;
#1 $display("%b", po);
# 1  pi=13'b0001000101110;
#1 $display("%b", po);
# 1  pi=13'b0001000101111;
#1 $display("%b", po);
# 1  pi=13'b0001000110000;
#1 $display("%b", po);
# 1  pi=13'b0001000110001;
#1 $display("%b", po);
# 1  pi=13'b0001000110010;
#1 $display("%b", po);
# 1  pi=13'b0001000110011;
#1 $display("%b", po);
# 1  pi=13'b0001000110100;
#1 $display("%b", po);
# 1  pi=13'b0001000110101;
#1 $display("%b", po);
# 1  pi=13'b0001000110110;
#1 $display("%b", po);
# 1  pi=13'b0001000110111;
#1 $display("%b", po);
# 1  pi=13'b0001000111000;
#1 $display("%b", po);
# 1  pi=13'b0001000111001;
#1 $display("%b", po);
# 1  pi=13'b0001000111010;
#1 $display("%b", po);
# 1  pi=13'b0001000111011;
#1 $display("%b", po);
# 1  pi=13'b0001000111100;
#1 $display("%b", po);
# 1  pi=13'b0001000111101;
#1 $display("%b", po);
# 1  pi=13'b0001000111110;
#1 $display("%b", po);
# 1  pi=13'b0001000111111;
#1 $display("%b", po);
# 1  pi=13'b0001001000000;
#1 $display("%b", po);
# 1  pi=13'b0001001000001;
#1 $display("%b", po);
# 1  pi=13'b0001001000010;
#1 $display("%b", po);
# 1  pi=13'b0001001000011;
#1 $display("%b", po);
# 1  pi=13'b0001001000100;
#1 $display("%b", po);
# 1  pi=13'b0001001000101;
#1 $display("%b", po);
# 1  pi=13'b0001001000110;
#1 $display("%b", po);
# 1  pi=13'b0001001000111;
#1 $display("%b", po);
# 1  pi=13'b0001001001000;
#1 $display("%b", po);
# 1  pi=13'b0001001001001;
#1 $display("%b", po);
# 1  pi=13'b0001001001010;
#1 $display("%b", po);
# 1  pi=13'b0001001001011;
#1 $display("%b", po);
# 1  pi=13'b0001001001100;
#1 $display("%b", po);
# 1  pi=13'b0001001001101;
#1 $display("%b", po);
# 1  pi=13'b0001001001110;
#1 $display("%b", po);
# 1  pi=13'b0001001001111;
#1 $display("%b", po);
# 1  pi=13'b0001001010000;
#1 $display("%b", po);
# 1  pi=13'b0001001010001;
#1 $display("%b", po);
# 1  pi=13'b0001001010010;
#1 $display("%b", po);
# 1  pi=13'b0001001010011;
#1 $display("%b", po);
# 1  pi=13'b0001001010100;
#1 $display("%b", po);
# 1  pi=13'b0001001010101;
#1 $display("%b", po);
# 1  pi=13'b0001001010110;
#1 $display("%b", po);
# 1  pi=13'b0001001010111;
#1 $display("%b", po);
# 1  pi=13'b0001001011000;
#1 $display("%b", po);
# 1  pi=13'b0001001011001;
#1 $display("%b", po);
# 1  pi=13'b0001001011010;
#1 $display("%b", po);
# 1  pi=13'b0001001011011;
#1 $display("%b", po);
# 1  pi=13'b0001001011100;
#1 $display("%b", po);
# 1  pi=13'b0001001011101;
#1 $display("%b", po);
# 1  pi=13'b0001001011110;
#1 $display("%b", po);
# 1  pi=13'b0001001011111;
#1 $display("%b", po);
# 1  pi=13'b0001001100000;
#1 $display("%b", po);
# 1  pi=13'b0001001100001;
#1 $display("%b", po);
# 1  pi=13'b0001001100010;
#1 $display("%b", po);
# 1  pi=13'b0001001100011;
#1 $display("%b", po);
# 1  pi=13'b0001001100100;
#1 $display("%b", po);
# 1  pi=13'b0001001100101;
#1 $display("%b", po);
# 1  pi=13'b0001001100110;
#1 $display("%b", po);
# 1  pi=13'b0001001100111;
#1 $display("%b", po);
# 1  pi=13'b0001001101000;
#1 $display("%b", po);
# 1  pi=13'b0001001101001;
#1 $display("%b", po);
# 1  pi=13'b0001001101010;
#1 $display("%b", po);
# 1  pi=13'b0001001101011;
#1 $display("%b", po);
# 1  pi=13'b0001001101100;
#1 $display("%b", po);
# 1  pi=13'b0001001101101;
#1 $display("%b", po);
# 1  pi=13'b0001001101110;
#1 $display("%b", po);
# 1  pi=13'b0001001101111;
#1 $display("%b", po);
# 1  pi=13'b0001001110000;
#1 $display("%b", po);
# 1  pi=13'b0001001110001;
#1 $display("%b", po);
# 1  pi=13'b0001001110010;
#1 $display("%b", po);
# 1  pi=13'b0001001110011;
#1 $display("%b", po);
# 1  pi=13'b0001001110100;
#1 $display("%b", po);
# 1  pi=13'b0001001110101;
#1 $display("%b", po);
# 1  pi=13'b0001001110110;
#1 $display("%b", po);
# 1  pi=13'b0001001110111;
#1 $display("%b", po);
# 1  pi=13'b0001001111000;
#1 $display("%b", po);
# 1  pi=13'b0001001111001;
#1 $display("%b", po);
# 1  pi=13'b0001001111010;
#1 $display("%b", po);
# 1  pi=13'b0001001111011;
#1 $display("%b", po);
# 1  pi=13'b0001001111100;
#1 $display("%b", po);
# 1  pi=13'b0001001111101;
#1 $display("%b", po);
# 1  pi=13'b0001001111110;
#1 $display("%b", po);
# 1  pi=13'b0001001111111;
#1 $display("%b", po);
# 1  pi=13'b0001010000000;
#1 $display("%b", po);
# 1  pi=13'b0001010000001;
#1 $display("%b", po);
# 1  pi=13'b0001010000010;
#1 $display("%b", po);
# 1  pi=13'b0001010000011;
#1 $display("%b", po);
# 1  pi=13'b0001010000100;
#1 $display("%b", po);
# 1  pi=13'b0001010000101;
#1 $display("%b", po);
# 1  pi=13'b0001010000110;
#1 $display("%b", po);
# 1  pi=13'b0001010000111;
#1 $display("%b", po);
# 1  pi=13'b0001010001000;
#1 $display("%b", po);
# 1  pi=13'b0001010001001;
#1 $display("%b", po);
# 1  pi=13'b0001010001010;
#1 $display("%b", po);
# 1  pi=13'b0001010001011;
#1 $display("%b", po);
# 1  pi=13'b0001010001100;
#1 $display("%b", po);
# 1  pi=13'b0001010001101;
#1 $display("%b", po);
# 1  pi=13'b0001010001110;
#1 $display("%b", po);
# 1  pi=13'b0001010001111;
#1 $display("%b", po);
# 1  pi=13'b0001010010000;
#1 $display("%b", po);
# 1  pi=13'b0001010010001;
#1 $display("%b", po);
# 1  pi=13'b0001010010010;
#1 $display("%b", po);
# 1  pi=13'b0001010010011;
#1 $display("%b", po);
# 1  pi=13'b0001010010100;
#1 $display("%b", po);
# 1  pi=13'b0001010010101;
#1 $display("%b", po);
# 1  pi=13'b0001010010110;
#1 $display("%b", po);
# 1  pi=13'b0001010010111;
#1 $display("%b", po);
# 1  pi=13'b0001010011000;
#1 $display("%b", po);
# 1  pi=13'b0001010011001;
#1 $display("%b", po);
# 1  pi=13'b0001010011010;
#1 $display("%b", po);
# 1  pi=13'b0001010011011;
#1 $display("%b", po);
# 1  pi=13'b0001010011100;
#1 $display("%b", po);
# 1  pi=13'b0001010011101;
#1 $display("%b", po);
# 1  pi=13'b0001010011110;
#1 $display("%b", po);
# 1  pi=13'b0001010011111;
#1 $display("%b", po);
# 1  pi=13'b0001010100000;
#1 $display("%b", po);
# 1  pi=13'b0001010100001;
#1 $display("%b", po);
# 1  pi=13'b0001010100010;
#1 $display("%b", po);
# 1  pi=13'b0001010100011;
#1 $display("%b", po);
# 1  pi=13'b0001010100100;
#1 $display("%b", po);
# 1  pi=13'b0001010100101;
#1 $display("%b", po);
# 1  pi=13'b0001010100110;
#1 $display("%b", po);
# 1  pi=13'b0001010100111;
#1 $display("%b", po);
# 1  pi=13'b0001010101000;
#1 $display("%b", po);
# 1  pi=13'b0001010101001;
#1 $display("%b", po);
# 1  pi=13'b0001010101010;
#1 $display("%b", po);
# 1  pi=13'b0001010101011;
#1 $display("%b", po);
# 1  pi=13'b0001010101100;
#1 $display("%b", po);
# 1  pi=13'b0001010101101;
#1 $display("%b", po);
# 1  pi=13'b0001010101110;
#1 $display("%b", po);
# 1  pi=13'b0001010101111;
#1 $display("%b", po);
# 1  pi=13'b0001010110000;
#1 $display("%b", po);
# 1  pi=13'b0001010110001;
#1 $display("%b", po);
# 1  pi=13'b0001010110010;
#1 $display("%b", po);
# 1  pi=13'b0001010110011;
#1 $display("%b", po);
# 1  pi=13'b0001010110100;
#1 $display("%b", po);
# 1  pi=13'b0001010110101;
#1 $display("%b", po);
# 1  pi=13'b0001010110110;
#1 $display("%b", po);
# 1  pi=13'b0001010110111;
#1 $display("%b", po);
# 1  pi=13'b0001010111000;
#1 $display("%b", po);
# 1  pi=13'b0001010111001;
#1 $display("%b", po);
# 1  pi=13'b0001010111010;
#1 $display("%b", po);
# 1  pi=13'b0001010111011;
#1 $display("%b", po);
# 1  pi=13'b0001010111100;
#1 $display("%b", po);
# 1  pi=13'b0001010111101;
#1 $display("%b", po);
# 1  pi=13'b0001010111110;
#1 $display("%b", po);
# 1  pi=13'b0001010111111;
#1 $display("%b", po);
# 1  pi=13'b0001011000000;
#1 $display("%b", po);
# 1  pi=13'b0001011000001;
#1 $display("%b", po);
# 1  pi=13'b0001011000010;
#1 $display("%b", po);
# 1  pi=13'b0001011000011;
#1 $display("%b", po);
# 1  pi=13'b0001011000100;
#1 $display("%b", po);
# 1  pi=13'b0001011000101;
#1 $display("%b", po);
# 1  pi=13'b0001011000110;
#1 $display("%b", po);
# 1  pi=13'b0001011000111;
#1 $display("%b", po);
# 1  pi=13'b0001011001000;
#1 $display("%b", po);
# 1  pi=13'b0001011001001;
#1 $display("%b", po);
# 1  pi=13'b0001011001010;
#1 $display("%b", po);
# 1  pi=13'b0001011001011;
#1 $display("%b", po);
# 1  pi=13'b0001011001100;
#1 $display("%b", po);
# 1  pi=13'b0001011001101;
#1 $display("%b", po);
# 1  pi=13'b0001011001110;
#1 $display("%b", po);
# 1  pi=13'b0001011001111;
#1 $display("%b", po);
# 1  pi=13'b0001011010000;
#1 $display("%b", po);
# 1  pi=13'b0001011010001;
#1 $display("%b", po);
# 1  pi=13'b0001011010010;
#1 $display("%b", po);
# 1  pi=13'b0001011010011;
#1 $display("%b", po);
# 1  pi=13'b0001011010100;
#1 $display("%b", po);
# 1  pi=13'b0001011010101;
#1 $display("%b", po);
# 1  pi=13'b0001011010110;
#1 $display("%b", po);
# 1  pi=13'b0001011010111;
#1 $display("%b", po);
# 1  pi=13'b0001011011000;
#1 $display("%b", po);
# 1  pi=13'b0001011011001;
#1 $display("%b", po);
# 1  pi=13'b0001011011010;
#1 $display("%b", po);
# 1  pi=13'b0001011011011;
#1 $display("%b", po);
# 1  pi=13'b0001011011100;
#1 $display("%b", po);
# 1  pi=13'b0001011011101;
#1 $display("%b", po);
# 1  pi=13'b0001011011110;
#1 $display("%b", po);
# 1  pi=13'b0001011011111;
#1 $display("%b", po);
# 1  pi=13'b0001011100000;
#1 $display("%b", po);
# 1  pi=13'b0001011100001;
#1 $display("%b", po);
# 1  pi=13'b0001011100010;
#1 $display("%b", po);
# 1  pi=13'b0001011100011;
#1 $display("%b", po);
# 1  pi=13'b0001011100100;
#1 $display("%b", po);
# 1  pi=13'b0001011100101;
#1 $display("%b", po);
# 1  pi=13'b0001011100110;
#1 $display("%b", po);
# 1  pi=13'b0001011100111;
#1 $display("%b", po);
# 1  pi=13'b0001011101000;
#1 $display("%b", po);
# 1  pi=13'b0001011101001;
#1 $display("%b", po);
# 1  pi=13'b0001011101010;
#1 $display("%b", po);
# 1  pi=13'b0001011101011;
#1 $display("%b", po);
# 1  pi=13'b0001011101100;
#1 $display("%b", po);
# 1  pi=13'b0001011101101;
#1 $display("%b", po);
# 1  pi=13'b0001011101110;
#1 $display("%b", po);
# 1  pi=13'b0001011101111;
#1 $display("%b", po);
# 1  pi=13'b0001011110000;
#1 $display("%b", po);
# 1  pi=13'b0001011110001;
#1 $display("%b", po);
# 1  pi=13'b0001011110010;
#1 $display("%b", po);
# 1  pi=13'b0001011110011;
#1 $display("%b", po);
# 1  pi=13'b0001011110100;
#1 $display("%b", po);
# 1  pi=13'b0001011110101;
#1 $display("%b", po);
# 1  pi=13'b0001011110110;
#1 $display("%b", po);
# 1  pi=13'b0001011110111;
#1 $display("%b", po);
# 1  pi=13'b0001011111000;
#1 $display("%b", po);
# 1  pi=13'b0001011111001;
#1 $display("%b", po);
# 1  pi=13'b0001011111010;
#1 $display("%b", po);
# 1  pi=13'b0001011111011;
#1 $display("%b", po);
# 1  pi=13'b0001011111100;
#1 $display("%b", po);
# 1  pi=13'b0001011111101;
#1 $display("%b", po);
# 1  pi=13'b0001011111110;
#1 $display("%b", po);
# 1  pi=13'b0001011111111;
#1 $display("%b", po);
# 1  pi=13'b0001100000000;
#1 $display("%b", po);
# 1  pi=13'b0001100000001;
#1 $display("%b", po);
# 1  pi=13'b0001100000010;
#1 $display("%b", po);
# 1  pi=13'b0001100000011;
#1 $display("%b", po);
# 1  pi=13'b0001100000100;
#1 $display("%b", po);
# 1  pi=13'b0001100000101;
#1 $display("%b", po);
# 1  pi=13'b0001100000110;
#1 $display("%b", po);
# 1  pi=13'b0001100000111;
#1 $display("%b", po);
# 1  pi=13'b0001100001000;
#1 $display("%b", po);
# 1  pi=13'b0001100001001;
#1 $display("%b", po);
# 1  pi=13'b0001100001010;
#1 $display("%b", po);
# 1  pi=13'b0001100001011;
#1 $display("%b", po);
# 1  pi=13'b0001100001100;
#1 $display("%b", po);
# 1  pi=13'b0001100001101;
#1 $display("%b", po);
# 1  pi=13'b0001100001110;
#1 $display("%b", po);
# 1  pi=13'b0001100001111;
#1 $display("%b", po);
# 1  pi=13'b0001100010000;
#1 $display("%b", po);
# 1  pi=13'b0001100010001;
#1 $display("%b", po);
# 1  pi=13'b0001100010010;
#1 $display("%b", po);
# 1  pi=13'b0001100010011;
#1 $display("%b", po);
# 1  pi=13'b0001100010100;
#1 $display("%b", po);
# 1  pi=13'b0001100010101;
#1 $display("%b", po);
# 1  pi=13'b0001100010110;
#1 $display("%b", po);
# 1  pi=13'b0001100010111;
#1 $display("%b", po);
# 1  pi=13'b0001100011000;
#1 $display("%b", po);
# 1  pi=13'b0001100011001;
#1 $display("%b", po);
# 1  pi=13'b0001100011010;
#1 $display("%b", po);
# 1  pi=13'b0001100011011;
#1 $display("%b", po);
# 1  pi=13'b0001100011100;
#1 $display("%b", po);
# 1  pi=13'b0001100011101;
#1 $display("%b", po);
# 1  pi=13'b0001100011110;
#1 $display("%b", po);
# 1  pi=13'b0001100011111;
#1 $display("%b", po);
# 1  pi=13'b0001100100000;
#1 $display("%b", po);
# 1  pi=13'b0001100100001;
#1 $display("%b", po);
# 1  pi=13'b0001100100010;
#1 $display("%b", po);
# 1  pi=13'b0001100100011;
#1 $display("%b", po);
# 1  pi=13'b0001100100100;
#1 $display("%b", po);
# 1  pi=13'b0001100100101;
#1 $display("%b", po);
# 1  pi=13'b0001100100110;
#1 $display("%b", po);
# 1  pi=13'b0001100100111;
#1 $display("%b", po);
# 1  pi=13'b0001100101000;
#1 $display("%b", po);
# 1  pi=13'b0001100101001;
#1 $display("%b", po);
# 1  pi=13'b0001100101010;
#1 $display("%b", po);
# 1  pi=13'b0001100101011;
#1 $display("%b", po);
# 1  pi=13'b0001100101100;
#1 $display("%b", po);
# 1  pi=13'b0001100101101;
#1 $display("%b", po);
# 1  pi=13'b0001100101110;
#1 $display("%b", po);
# 1  pi=13'b0001100101111;
#1 $display("%b", po);
# 1  pi=13'b0001100110000;
#1 $display("%b", po);
# 1  pi=13'b0001100110001;
#1 $display("%b", po);
# 1  pi=13'b0001100110010;
#1 $display("%b", po);
# 1  pi=13'b0001100110011;
#1 $display("%b", po);
# 1  pi=13'b0001100110100;
#1 $display("%b", po);
# 1  pi=13'b0001100110101;
#1 $display("%b", po);
# 1  pi=13'b0001100110110;
#1 $display("%b", po);
# 1  pi=13'b0001100110111;
#1 $display("%b", po);
# 1  pi=13'b0001100111000;
#1 $display("%b", po);
# 1  pi=13'b0001100111001;
#1 $display("%b", po);
# 1  pi=13'b0001100111010;
#1 $display("%b", po);
# 1  pi=13'b0001100111011;
#1 $display("%b", po);
# 1  pi=13'b0001100111100;
#1 $display("%b", po);
# 1  pi=13'b0001100111101;
#1 $display("%b", po);
# 1  pi=13'b0001100111110;
#1 $display("%b", po);
# 1  pi=13'b0001100111111;
#1 $display("%b", po);
# 1  pi=13'b0001101000000;
#1 $display("%b", po);
# 1  pi=13'b0001101000001;
#1 $display("%b", po);
# 1  pi=13'b0001101000010;
#1 $display("%b", po);
# 1  pi=13'b0001101000011;
#1 $display("%b", po);
# 1  pi=13'b0001101000100;
#1 $display("%b", po);
# 1  pi=13'b0001101000101;
#1 $display("%b", po);
# 1  pi=13'b0001101000110;
#1 $display("%b", po);
# 1  pi=13'b0001101000111;
#1 $display("%b", po);
# 1  pi=13'b0001101001000;
#1 $display("%b", po);
# 1  pi=13'b0001101001001;
#1 $display("%b", po);
# 1  pi=13'b0001101001010;
#1 $display("%b", po);
# 1  pi=13'b0001101001011;
#1 $display("%b", po);
# 1  pi=13'b0001101001100;
#1 $display("%b", po);
# 1  pi=13'b0001101001101;
#1 $display("%b", po);
# 1  pi=13'b0001101001110;
#1 $display("%b", po);
# 1  pi=13'b0001101001111;
#1 $display("%b", po);
# 1  pi=13'b0001101010000;
#1 $display("%b", po);
# 1  pi=13'b0001101010001;
#1 $display("%b", po);
# 1  pi=13'b0001101010010;
#1 $display("%b", po);
# 1  pi=13'b0001101010011;
#1 $display("%b", po);
# 1  pi=13'b0001101010100;
#1 $display("%b", po);
# 1  pi=13'b0001101010101;
#1 $display("%b", po);
# 1  pi=13'b0001101010110;
#1 $display("%b", po);
# 1  pi=13'b0001101010111;
#1 $display("%b", po);
# 1  pi=13'b0001101011000;
#1 $display("%b", po);
# 1  pi=13'b0001101011001;
#1 $display("%b", po);
# 1  pi=13'b0001101011010;
#1 $display("%b", po);
# 1  pi=13'b0001101011011;
#1 $display("%b", po);
# 1  pi=13'b0001101011100;
#1 $display("%b", po);
# 1  pi=13'b0001101011101;
#1 $display("%b", po);
# 1  pi=13'b0001101011110;
#1 $display("%b", po);
# 1  pi=13'b0001101011111;
#1 $display("%b", po);
# 1  pi=13'b0001101100000;
#1 $display("%b", po);
# 1  pi=13'b0001101100001;
#1 $display("%b", po);
# 1  pi=13'b0001101100010;
#1 $display("%b", po);
# 1  pi=13'b0001101100011;
#1 $display("%b", po);
# 1  pi=13'b0001101100100;
#1 $display("%b", po);
# 1  pi=13'b0001101100101;
#1 $display("%b", po);
# 1  pi=13'b0001101100110;
#1 $display("%b", po);
# 1  pi=13'b0001101100111;
#1 $display("%b", po);
# 1  pi=13'b0001101101000;
#1 $display("%b", po);
# 1  pi=13'b0001101101001;
#1 $display("%b", po);
# 1  pi=13'b0001101101010;
#1 $display("%b", po);
# 1  pi=13'b0001101101011;
#1 $display("%b", po);
# 1  pi=13'b0001101101100;
#1 $display("%b", po);
# 1  pi=13'b0001101101101;
#1 $display("%b", po);
# 1  pi=13'b0001101101110;
#1 $display("%b", po);
# 1  pi=13'b0001101101111;
#1 $display("%b", po);
# 1  pi=13'b0001101110000;
#1 $display("%b", po);
# 1  pi=13'b0001101110001;
#1 $display("%b", po);
# 1  pi=13'b0001101110010;
#1 $display("%b", po);
# 1  pi=13'b0001101110011;
#1 $display("%b", po);
# 1  pi=13'b0001101110100;
#1 $display("%b", po);
# 1  pi=13'b0001101110101;
#1 $display("%b", po);
# 1  pi=13'b0001101110110;
#1 $display("%b", po);
# 1  pi=13'b0001101110111;
#1 $display("%b", po);
# 1  pi=13'b0001101111000;
#1 $display("%b", po);
# 1  pi=13'b0001101111001;
#1 $display("%b", po);
# 1  pi=13'b0001101111010;
#1 $display("%b", po);
# 1  pi=13'b0001101111011;
#1 $display("%b", po);
# 1  pi=13'b0001101111100;
#1 $display("%b", po);
# 1  pi=13'b0001101111101;
#1 $display("%b", po);
# 1  pi=13'b0001101111110;
#1 $display("%b", po);
# 1  pi=13'b0001101111111;
#1 $display("%b", po);
# 1  pi=13'b0001110000000;
#1 $display("%b", po);
# 1  pi=13'b0001110000001;
#1 $display("%b", po);
# 1  pi=13'b0001110000010;
#1 $display("%b", po);
# 1  pi=13'b0001110000011;
#1 $display("%b", po);
# 1  pi=13'b0001110000100;
#1 $display("%b", po);
# 1  pi=13'b0001110000101;
#1 $display("%b", po);
# 1  pi=13'b0001110000110;
#1 $display("%b", po);
# 1  pi=13'b0001110000111;
#1 $display("%b", po);
# 1  pi=13'b0001110001000;
#1 $display("%b", po);
# 1  pi=13'b0001110001001;
#1 $display("%b", po);
# 1  pi=13'b0001110001010;
#1 $display("%b", po);
# 1  pi=13'b0001110001011;
#1 $display("%b", po);
# 1  pi=13'b0001110001100;
#1 $display("%b", po);
# 1  pi=13'b0001110001101;
#1 $display("%b", po);
# 1  pi=13'b0001110001110;
#1 $display("%b", po);
# 1  pi=13'b0001110001111;
#1 $display("%b", po);
# 1  pi=13'b0001110010000;
#1 $display("%b", po);
# 1  pi=13'b0001110010001;
#1 $display("%b", po);
# 1  pi=13'b0001110010010;
#1 $display("%b", po);
# 1  pi=13'b0001110010011;
#1 $display("%b", po);
# 1  pi=13'b0001110010100;
#1 $display("%b", po);
# 1  pi=13'b0001110010101;
#1 $display("%b", po);
# 1  pi=13'b0001110010110;
#1 $display("%b", po);
# 1  pi=13'b0001110010111;
#1 $display("%b", po);
# 1  pi=13'b0001110011000;
#1 $display("%b", po);
# 1  pi=13'b0001110011001;
#1 $display("%b", po);
# 1  pi=13'b0001110011010;
#1 $display("%b", po);
# 1  pi=13'b0001110011011;
#1 $display("%b", po);
# 1  pi=13'b0001110011100;
#1 $display("%b", po);
# 1  pi=13'b0001110011101;
#1 $display("%b", po);
# 1  pi=13'b0001110011110;
#1 $display("%b", po);
# 1  pi=13'b0001110011111;
#1 $display("%b", po);
# 1  pi=13'b0001110100000;
#1 $display("%b", po);
# 1  pi=13'b0001110100001;
#1 $display("%b", po);
# 1  pi=13'b0001110100010;
#1 $display("%b", po);
# 1  pi=13'b0001110100011;
#1 $display("%b", po);
# 1  pi=13'b0001110100100;
#1 $display("%b", po);
# 1  pi=13'b0001110100101;
#1 $display("%b", po);
# 1  pi=13'b0001110100110;
#1 $display("%b", po);
# 1  pi=13'b0001110100111;
#1 $display("%b", po);
# 1  pi=13'b0001110101000;
#1 $display("%b", po);
# 1  pi=13'b0001110101001;
#1 $display("%b", po);
# 1  pi=13'b0001110101010;
#1 $display("%b", po);
# 1  pi=13'b0001110101011;
#1 $display("%b", po);
# 1  pi=13'b0001110101100;
#1 $display("%b", po);
# 1  pi=13'b0001110101101;
#1 $display("%b", po);
# 1  pi=13'b0001110101110;
#1 $display("%b", po);
# 1  pi=13'b0001110101111;
#1 $display("%b", po);
# 1  pi=13'b0001110110000;
#1 $display("%b", po);
# 1  pi=13'b0001110110001;
#1 $display("%b", po);
# 1  pi=13'b0001110110010;
#1 $display("%b", po);
# 1  pi=13'b0001110110011;
#1 $display("%b", po);
# 1  pi=13'b0001110110100;
#1 $display("%b", po);
# 1  pi=13'b0001110110101;
#1 $display("%b", po);
# 1  pi=13'b0001110110110;
#1 $display("%b", po);
# 1  pi=13'b0001110110111;
#1 $display("%b", po);
# 1  pi=13'b0001110111000;
#1 $display("%b", po);
# 1  pi=13'b0001110111001;
#1 $display("%b", po);
# 1  pi=13'b0001110111010;
#1 $display("%b", po);
# 1  pi=13'b0001110111011;
#1 $display("%b", po);
# 1  pi=13'b0001110111100;
#1 $display("%b", po);
# 1  pi=13'b0001110111101;
#1 $display("%b", po);
# 1  pi=13'b0001110111110;
#1 $display("%b", po);
# 1  pi=13'b0001110111111;
#1 $display("%b", po);
# 1  pi=13'b0001111000000;
#1 $display("%b", po);
# 1  pi=13'b0001111000001;
#1 $display("%b", po);
# 1  pi=13'b0001111000010;
#1 $display("%b", po);
# 1  pi=13'b0001111000011;
#1 $display("%b", po);
# 1  pi=13'b0001111000100;
#1 $display("%b", po);
# 1  pi=13'b0001111000101;
#1 $display("%b", po);
# 1  pi=13'b0001111000110;
#1 $display("%b", po);
# 1  pi=13'b0001111000111;
#1 $display("%b", po);
# 1  pi=13'b0001111001000;
#1 $display("%b", po);
# 1  pi=13'b0001111001001;
#1 $display("%b", po);
# 1  pi=13'b0001111001010;
#1 $display("%b", po);
# 1  pi=13'b0001111001011;
#1 $display("%b", po);
# 1  pi=13'b0001111001100;
#1 $display("%b", po);
# 1  pi=13'b0001111001101;
#1 $display("%b", po);
# 1  pi=13'b0001111001110;
#1 $display("%b", po);
# 1  pi=13'b0001111001111;
#1 $display("%b", po);
# 1  pi=13'b0001111010000;
#1 $display("%b", po);
# 1  pi=13'b0001111010001;
#1 $display("%b", po);
# 1  pi=13'b0001111010010;
#1 $display("%b", po);
# 1  pi=13'b0001111010011;
#1 $display("%b", po);
# 1  pi=13'b0001111010100;
#1 $display("%b", po);
# 1  pi=13'b0001111010101;
#1 $display("%b", po);
# 1  pi=13'b0001111010110;
#1 $display("%b", po);
# 1  pi=13'b0001111010111;
#1 $display("%b", po);
# 1  pi=13'b0001111011000;
#1 $display("%b", po);
# 1  pi=13'b0001111011001;
#1 $display("%b", po);
# 1  pi=13'b0001111011010;
#1 $display("%b", po);
# 1  pi=13'b0001111011011;
#1 $display("%b", po);
# 1  pi=13'b0001111011100;
#1 $display("%b", po);
# 1  pi=13'b0001111011101;
#1 $display("%b", po);
# 1  pi=13'b0001111011110;
#1 $display("%b", po);
# 1  pi=13'b0001111011111;
#1 $display("%b", po);
# 1  pi=13'b0001111100000;
#1 $display("%b", po);
# 1  pi=13'b0001111100001;
#1 $display("%b", po);
# 1  pi=13'b0001111100010;
#1 $display("%b", po);
# 1  pi=13'b0001111100011;
#1 $display("%b", po);
# 1  pi=13'b0001111100100;
#1 $display("%b", po);
# 1  pi=13'b0001111100101;
#1 $display("%b", po);
# 1  pi=13'b0001111100110;
#1 $display("%b", po);
# 1  pi=13'b0001111100111;
#1 $display("%b", po);
# 1  pi=13'b0001111101000;
#1 $display("%b", po);
# 1  pi=13'b0001111101001;
#1 $display("%b", po);
# 1  pi=13'b0001111101010;
#1 $display("%b", po);
# 1  pi=13'b0001111101011;
#1 $display("%b", po);
# 1  pi=13'b0001111101100;
#1 $display("%b", po);
# 1  pi=13'b0001111101101;
#1 $display("%b", po);
# 1  pi=13'b0001111101110;
#1 $display("%b", po);
# 1  pi=13'b0001111101111;
#1 $display("%b", po);
# 1  pi=13'b0001111110000;
#1 $display("%b", po);
# 1  pi=13'b0001111110001;
#1 $display("%b", po);
# 1  pi=13'b0001111110010;
#1 $display("%b", po);
# 1  pi=13'b0001111110011;
#1 $display("%b", po);
# 1  pi=13'b0001111110100;
#1 $display("%b", po);
# 1  pi=13'b0001111110101;
#1 $display("%b", po);
# 1  pi=13'b0001111110110;
#1 $display("%b", po);
# 1  pi=13'b0001111110111;
#1 $display("%b", po);
# 1  pi=13'b0001111111000;
#1 $display("%b", po);
# 1  pi=13'b0001111111001;
#1 $display("%b", po);
# 1  pi=13'b0001111111010;
#1 $display("%b", po);
# 1  pi=13'b0001111111011;
#1 $display("%b", po);
# 1  pi=13'b0001111111100;
#1 $display("%b", po);
# 1  pi=13'b0001111111101;
#1 $display("%b", po);
# 1  pi=13'b0001111111110;
#1 $display("%b", po);
# 1  pi=13'b0001111111111;
#1 $display("%b", po);
# 1  pi=13'b0010000000000;
#1 $display("%b", po);
# 1  pi=13'b0010000000001;
#1 $display("%b", po);
# 1  pi=13'b0010000000010;
#1 $display("%b", po);
# 1  pi=13'b0010000000011;
#1 $display("%b", po);
# 1  pi=13'b0010000000100;
#1 $display("%b", po);
# 1  pi=13'b0010000000101;
#1 $display("%b", po);
# 1  pi=13'b0010000000110;
#1 $display("%b", po);
# 1  pi=13'b0010000000111;
#1 $display("%b", po);
# 1  pi=13'b0010000001000;
#1 $display("%b", po);
# 1  pi=13'b0010000001001;
#1 $display("%b", po);
# 1  pi=13'b0010000001010;
#1 $display("%b", po);
# 1  pi=13'b0010000001011;
#1 $display("%b", po);
# 1  pi=13'b0010000001100;
#1 $display("%b", po);
# 1  pi=13'b0010000001101;
#1 $display("%b", po);
# 1  pi=13'b0010000001110;
#1 $display("%b", po);
# 1  pi=13'b0010000001111;
#1 $display("%b", po);
# 1  pi=13'b0010000010000;
#1 $display("%b", po);
# 1  pi=13'b0010000010001;
#1 $display("%b", po);
# 1  pi=13'b0010000010010;
#1 $display("%b", po);
# 1  pi=13'b0010000010011;
#1 $display("%b", po);
# 1  pi=13'b0010000010100;
#1 $display("%b", po);
# 1  pi=13'b0010000010101;
#1 $display("%b", po);
# 1  pi=13'b0010000010110;
#1 $display("%b", po);
# 1  pi=13'b0010000010111;
#1 $display("%b", po);
# 1  pi=13'b0010000011000;
#1 $display("%b", po);
# 1  pi=13'b0010000011001;
#1 $display("%b", po);
# 1  pi=13'b0010000011010;
#1 $display("%b", po);
# 1  pi=13'b0010000011011;
#1 $display("%b", po);
# 1  pi=13'b0010000011100;
#1 $display("%b", po);
# 1  pi=13'b0010000011101;
#1 $display("%b", po);
# 1  pi=13'b0010000011110;
#1 $display("%b", po);
# 1  pi=13'b0010000011111;
#1 $display("%b", po);
# 1  pi=13'b0010000100000;
#1 $display("%b", po);
# 1  pi=13'b0010000100001;
#1 $display("%b", po);
# 1  pi=13'b0010000100010;
#1 $display("%b", po);
# 1  pi=13'b0010000100011;
#1 $display("%b", po);
# 1  pi=13'b0010000100100;
#1 $display("%b", po);
# 1  pi=13'b0010000100101;
#1 $display("%b", po);
# 1  pi=13'b0010000100110;
#1 $display("%b", po);
# 1  pi=13'b0010000100111;
#1 $display("%b", po);
# 1  pi=13'b0010000101000;
#1 $display("%b", po);
# 1  pi=13'b0010000101001;
#1 $display("%b", po);
# 1  pi=13'b0010000101010;
#1 $display("%b", po);
# 1  pi=13'b0010000101011;
#1 $display("%b", po);
# 1  pi=13'b0010000101100;
#1 $display("%b", po);
# 1  pi=13'b0010000101101;
#1 $display("%b", po);
# 1  pi=13'b0010000101110;
#1 $display("%b", po);
# 1  pi=13'b0010000101111;
#1 $display("%b", po);
# 1  pi=13'b0010000110000;
#1 $display("%b", po);
# 1  pi=13'b0010000110001;
#1 $display("%b", po);
# 1  pi=13'b0010000110010;
#1 $display("%b", po);
# 1  pi=13'b0010000110011;
#1 $display("%b", po);
# 1  pi=13'b0010000110100;
#1 $display("%b", po);
# 1  pi=13'b0010000110101;
#1 $display("%b", po);
# 1  pi=13'b0010000110110;
#1 $display("%b", po);
# 1  pi=13'b0010000110111;
#1 $display("%b", po);
# 1  pi=13'b0010000111000;
#1 $display("%b", po);
# 1  pi=13'b0010000111001;
#1 $display("%b", po);
# 1  pi=13'b0010000111010;
#1 $display("%b", po);
# 1  pi=13'b0010000111011;
#1 $display("%b", po);
# 1  pi=13'b0010000111100;
#1 $display("%b", po);
# 1  pi=13'b0010000111101;
#1 $display("%b", po);
# 1  pi=13'b0010000111110;
#1 $display("%b", po);
# 1  pi=13'b0010000111111;
#1 $display("%b", po);
# 1  pi=13'b0010001000000;
#1 $display("%b", po);
# 1  pi=13'b0010001000001;
#1 $display("%b", po);
# 1  pi=13'b0010001000010;
#1 $display("%b", po);
# 1  pi=13'b0010001000011;
#1 $display("%b", po);
# 1  pi=13'b0010001000100;
#1 $display("%b", po);
# 1  pi=13'b0010001000101;
#1 $display("%b", po);
# 1  pi=13'b0010001000110;
#1 $display("%b", po);
# 1  pi=13'b0010001000111;
#1 $display("%b", po);
# 1  pi=13'b0010001001000;
#1 $display("%b", po);
# 1  pi=13'b0010001001001;
#1 $display("%b", po);
# 1  pi=13'b0010001001010;
#1 $display("%b", po);
# 1  pi=13'b0010001001011;
#1 $display("%b", po);
# 1  pi=13'b0010001001100;
#1 $display("%b", po);
# 1  pi=13'b0010001001101;
#1 $display("%b", po);
# 1  pi=13'b0010001001110;
#1 $display("%b", po);
# 1  pi=13'b0010001001111;
#1 $display("%b", po);
# 1  pi=13'b0010001010000;
#1 $display("%b", po);
# 1  pi=13'b0010001010001;
#1 $display("%b", po);
# 1  pi=13'b0010001010010;
#1 $display("%b", po);
# 1  pi=13'b0010001010011;
#1 $display("%b", po);
# 1  pi=13'b0010001010100;
#1 $display("%b", po);
# 1  pi=13'b0010001010101;
#1 $display("%b", po);
# 1  pi=13'b0010001010110;
#1 $display("%b", po);
# 1  pi=13'b0010001010111;
#1 $display("%b", po);
# 1  pi=13'b0010001011000;
#1 $display("%b", po);
# 1  pi=13'b0010001011001;
#1 $display("%b", po);
# 1  pi=13'b0010001011010;
#1 $display("%b", po);
# 1  pi=13'b0010001011011;
#1 $display("%b", po);
# 1  pi=13'b0010001011100;
#1 $display("%b", po);
# 1  pi=13'b0010001011101;
#1 $display("%b", po);
# 1  pi=13'b0010001011110;
#1 $display("%b", po);
# 1  pi=13'b0010001011111;
#1 $display("%b", po);
# 1  pi=13'b0010001100000;
#1 $display("%b", po);
# 1  pi=13'b0010001100001;
#1 $display("%b", po);
# 1  pi=13'b0010001100010;
#1 $display("%b", po);
# 1  pi=13'b0010001100011;
#1 $display("%b", po);
# 1  pi=13'b0010001100100;
#1 $display("%b", po);
# 1  pi=13'b0010001100101;
#1 $display("%b", po);
# 1  pi=13'b0010001100110;
#1 $display("%b", po);
# 1  pi=13'b0010001100111;
#1 $display("%b", po);
# 1  pi=13'b0010001101000;
#1 $display("%b", po);
# 1  pi=13'b0010001101001;
#1 $display("%b", po);
# 1  pi=13'b0010001101010;
#1 $display("%b", po);
# 1  pi=13'b0010001101011;
#1 $display("%b", po);
# 1  pi=13'b0010001101100;
#1 $display("%b", po);
# 1  pi=13'b0010001101101;
#1 $display("%b", po);
# 1  pi=13'b0010001101110;
#1 $display("%b", po);
# 1  pi=13'b0010001101111;
#1 $display("%b", po);
# 1  pi=13'b0010001110000;
#1 $display("%b", po);
# 1  pi=13'b0010001110001;
#1 $display("%b", po);
# 1  pi=13'b0010001110010;
#1 $display("%b", po);
# 1  pi=13'b0010001110011;
#1 $display("%b", po);
# 1  pi=13'b0010001110100;
#1 $display("%b", po);
# 1  pi=13'b0010001110101;
#1 $display("%b", po);
# 1  pi=13'b0010001110110;
#1 $display("%b", po);
# 1  pi=13'b0010001110111;
#1 $display("%b", po);
# 1  pi=13'b0010001111000;
#1 $display("%b", po);
# 1  pi=13'b0010001111001;
#1 $display("%b", po);
# 1  pi=13'b0010001111010;
#1 $display("%b", po);
# 1  pi=13'b0010001111011;
#1 $display("%b", po);
# 1  pi=13'b0010001111100;
#1 $display("%b", po);
# 1  pi=13'b0010001111101;
#1 $display("%b", po);
# 1  pi=13'b0010001111110;
#1 $display("%b", po);
# 1  pi=13'b0010001111111;
#1 $display("%b", po);
# 1  pi=13'b0010010000000;
#1 $display("%b", po);
# 1  pi=13'b0010010000001;
#1 $display("%b", po);
# 1  pi=13'b0010010000010;
#1 $display("%b", po);
# 1  pi=13'b0010010000011;
#1 $display("%b", po);
# 1  pi=13'b0010010000100;
#1 $display("%b", po);
# 1  pi=13'b0010010000101;
#1 $display("%b", po);
# 1  pi=13'b0010010000110;
#1 $display("%b", po);
# 1  pi=13'b0010010000111;
#1 $display("%b", po);
# 1  pi=13'b0010010001000;
#1 $display("%b", po);
# 1  pi=13'b0010010001001;
#1 $display("%b", po);
# 1  pi=13'b0010010001010;
#1 $display("%b", po);
# 1  pi=13'b0010010001011;
#1 $display("%b", po);
# 1  pi=13'b0010010001100;
#1 $display("%b", po);
# 1  pi=13'b0010010001101;
#1 $display("%b", po);
# 1  pi=13'b0010010001110;
#1 $display("%b", po);
# 1  pi=13'b0010010001111;
#1 $display("%b", po);
# 1  pi=13'b0010010010000;
#1 $display("%b", po);
# 1  pi=13'b0010010010001;
#1 $display("%b", po);
# 1  pi=13'b0010010010010;
#1 $display("%b", po);
# 1  pi=13'b0010010010011;
#1 $display("%b", po);
# 1  pi=13'b0010010010100;
#1 $display("%b", po);
# 1  pi=13'b0010010010101;
#1 $display("%b", po);
# 1  pi=13'b0010010010110;
#1 $display("%b", po);
# 1  pi=13'b0010010010111;
#1 $display("%b", po);
# 1  pi=13'b0010010011000;
#1 $display("%b", po);
# 1  pi=13'b0010010011001;
#1 $display("%b", po);
# 1  pi=13'b0010010011010;
#1 $display("%b", po);
# 1  pi=13'b0010010011011;
#1 $display("%b", po);
# 1  pi=13'b0010010011100;
#1 $display("%b", po);
# 1  pi=13'b0010010011101;
#1 $display("%b", po);
# 1  pi=13'b0010010011110;
#1 $display("%b", po);
# 1  pi=13'b0010010011111;
#1 $display("%b", po);
# 1  pi=13'b0010010100000;
#1 $display("%b", po);
# 1  pi=13'b0010010100001;
#1 $display("%b", po);
# 1  pi=13'b0010010100010;
#1 $display("%b", po);
# 1  pi=13'b0010010100011;
#1 $display("%b", po);
# 1  pi=13'b0010010100100;
#1 $display("%b", po);
# 1  pi=13'b0010010100101;
#1 $display("%b", po);
# 1  pi=13'b0010010100110;
#1 $display("%b", po);
# 1  pi=13'b0010010100111;
#1 $display("%b", po);
# 1  pi=13'b0010010101000;
#1 $display("%b", po);
# 1  pi=13'b0010010101001;
#1 $display("%b", po);
# 1  pi=13'b0010010101010;
#1 $display("%b", po);
# 1  pi=13'b0010010101011;
#1 $display("%b", po);
# 1  pi=13'b0010010101100;
#1 $display("%b", po);
# 1  pi=13'b0010010101101;
#1 $display("%b", po);
# 1  pi=13'b0010010101110;
#1 $display("%b", po);
# 1  pi=13'b0010010101111;
#1 $display("%b", po);
# 1  pi=13'b0010010110000;
#1 $display("%b", po);
# 1  pi=13'b0010010110001;
#1 $display("%b", po);
# 1  pi=13'b0010010110010;
#1 $display("%b", po);
# 1  pi=13'b0010010110011;
#1 $display("%b", po);
# 1  pi=13'b0010010110100;
#1 $display("%b", po);
# 1  pi=13'b0010010110101;
#1 $display("%b", po);
# 1  pi=13'b0010010110110;
#1 $display("%b", po);
# 1  pi=13'b0010010110111;
#1 $display("%b", po);
# 1  pi=13'b0010010111000;
#1 $display("%b", po);
# 1  pi=13'b0010010111001;
#1 $display("%b", po);
# 1  pi=13'b0010010111010;
#1 $display("%b", po);
# 1  pi=13'b0010010111011;
#1 $display("%b", po);
# 1  pi=13'b0010010111100;
#1 $display("%b", po);
# 1  pi=13'b0010010111101;
#1 $display("%b", po);
# 1  pi=13'b0010010111110;
#1 $display("%b", po);
# 1  pi=13'b0010010111111;
#1 $display("%b", po);
# 1  pi=13'b0010011000000;
#1 $display("%b", po);
# 1  pi=13'b0010011000001;
#1 $display("%b", po);
# 1  pi=13'b0010011000010;
#1 $display("%b", po);
# 1  pi=13'b0010011000011;
#1 $display("%b", po);
# 1  pi=13'b0010011000100;
#1 $display("%b", po);
# 1  pi=13'b0010011000101;
#1 $display("%b", po);
# 1  pi=13'b0010011000110;
#1 $display("%b", po);
# 1  pi=13'b0010011000111;
#1 $display("%b", po);
# 1  pi=13'b0010011001000;
#1 $display("%b", po);
# 1  pi=13'b0010011001001;
#1 $display("%b", po);
# 1  pi=13'b0010011001010;
#1 $display("%b", po);
# 1  pi=13'b0010011001011;
#1 $display("%b", po);
# 1  pi=13'b0010011001100;
#1 $display("%b", po);
# 1  pi=13'b0010011001101;
#1 $display("%b", po);
# 1  pi=13'b0010011001110;
#1 $display("%b", po);
# 1  pi=13'b0010011001111;
#1 $display("%b", po);
# 1  pi=13'b0010011010000;
#1 $display("%b", po);
# 1  pi=13'b0010011010001;
#1 $display("%b", po);
# 1  pi=13'b0010011010010;
#1 $display("%b", po);
# 1  pi=13'b0010011010011;
#1 $display("%b", po);
# 1  pi=13'b0010011010100;
#1 $display("%b", po);
# 1  pi=13'b0010011010101;
#1 $display("%b", po);
# 1  pi=13'b0010011010110;
#1 $display("%b", po);
# 1  pi=13'b0010011010111;
#1 $display("%b", po);
# 1  pi=13'b0010011011000;
#1 $display("%b", po);
# 1  pi=13'b0010011011001;
#1 $display("%b", po);
# 1  pi=13'b0010011011010;
#1 $display("%b", po);
# 1  pi=13'b0010011011011;
#1 $display("%b", po);
# 1  pi=13'b0010011011100;
#1 $display("%b", po);
# 1  pi=13'b0010011011101;
#1 $display("%b", po);
# 1  pi=13'b0010011011110;
#1 $display("%b", po);
# 1  pi=13'b0010011011111;
#1 $display("%b", po);
# 1  pi=13'b0010011100000;
#1 $display("%b", po);
# 1  pi=13'b0010011100001;
#1 $display("%b", po);
# 1  pi=13'b0010011100010;
#1 $display("%b", po);
# 1  pi=13'b0010011100011;
#1 $display("%b", po);
# 1  pi=13'b0010011100100;
#1 $display("%b", po);
# 1  pi=13'b0010011100101;
#1 $display("%b", po);
# 1  pi=13'b0010011100110;
#1 $display("%b", po);
# 1  pi=13'b0010011100111;
#1 $display("%b", po);
# 1  pi=13'b0010011101000;
#1 $display("%b", po);
# 1  pi=13'b0010011101001;
#1 $display("%b", po);
# 1  pi=13'b0010011101010;
#1 $display("%b", po);
# 1  pi=13'b0010011101011;
#1 $display("%b", po);
# 1  pi=13'b0010011101100;
#1 $display("%b", po);
# 1  pi=13'b0010011101101;
#1 $display("%b", po);
# 1  pi=13'b0010011101110;
#1 $display("%b", po);
# 1  pi=13'b0010011101111;
#1 $display("%b", po);
# 1  pi=13'b0010011110000;
#1 $display("%b", po);
# 1  pi=13'b0010011110001;
#1 $display("%b", po);
# 1  pi=13'b0010011110010;
#1 $display("%b", po);
# 1  pi=13'b0010011110011;
#1 $display("%b", po);
# 1  pi=13'b0010011110100;
#1 $display("%b", po);
# 1  pi=13'b0010011110101;
#1 $display("%b", po);
# 1  pi=13'b0010011110110;
#1 $display("%b", po);
# 1  pi=13'b0010011110111;
#1 $display("%b", po);
# 1  pi=13'b0010011111000;
#1 $display("%b", po);
# 1  pi=13'b0010011111001;
#1 $display("%b", po);
# 1  pi=13'b0010011111010;
#1 $display("%b", po);
# 1  pi=13'b0010011111011;
#1 $display("%b", po);
# 1  pi=13'b0010011111100;
#1 $display("%b", po);
# 1  pi=13'b0010011111101;
#1 $display("%b", po);
# 1  pi=13'b0010011111110;
#1 $display("%b", po);
# 1  pi=13'b0010011111111;
#1 $display("%b", po);
# 1  pi=13'b0010100000000;
#1 $display("%b", po);
# 1  pi=13'b0010100000001;
#1 $display("%b", po);
# 1  pi=13'b0010100000010;
#1 $display("%b", po);
# 1  pi=13'b0010100000011;
#1 $display("%b", po);
# 1  pi=13'b0010100000100;
#1 $display("%b", po);
# 1  pi=13'b0010100000101;
#1 $display("%b", po);
# 1  pi=13'b0010100000110;
#1 $display("%b", po);
# 1  pi=13'b0010100000111;
#1 $display("%b", po);
# 1  pi=13'b0010100001000;
#1 $display("%b", po);
# 1  pi=13'b0010100001001;
#1 $display("%b", po);
# 1  pi=13'b0010100001010;
#1 $display("%b", po);
# 1  pi=13'b0010100001011;
#1 $display("%b", po);
# 1  pi=13'b0010100001100;
#1 $display("%b", po);
# 1  pi=13'b0010100001101;
#1 $display("%b", po);
# 1  pi=13'b0010100001110;
#1 $display("%b", po);
# 1  pi=13'b0010100001111;
#1 $display("%b", po);
# 1  pi=13'b0010100010000;
#1 $display("%b", po);
# 1  pi=13'b0010100010001;
#1 $display("%b", po);
# 1  pi=13'b0010100010010;
#1 $display("%b", po);
# 1  pi=13'b0010100010011;
#1 $display("%b", po);
# 1  pi=13'b0010100010100;
#1 $display("%b", po);
# 1  pi=13'b0010100010101;
#1 $display("%b", po);
# 1  pi=13'b0010100010110;
#1 $display("%b", po);
# 1  pi=13'b0010100010111;
#1 $display("%b", po);
# 1  pi=13'b0010100011000;
#1 $display("%b", po);
# 1  pi=13'b0010100011001;
#1 $display("%b", po);
# 1  pi=13'b0010100011010;
#1 $display("%b", po);
# 1  pi=13'b0010100011011;
#1 $display("%b", po);
# 1  pi=13'b0010100011100;
#1 $display("%b", po);
# 1  pi=13'b0010100011101;
#1 $display("%b", po);
# 1  pi=13'b0010100011110;
#1 $display("%b", po);
# 1  pi=13'b0010100011111;
#1 $display("%b", po);
# 1  pi=13'b0010100100000;
#1 $display("%b", po);
# 1  pi=13'b0010100100001;
#1 $display("%b", po);
# 1  pi=13'b0010100100010;
#1 $display("%b", po);
# 1  pi=13'b0010100100011;
#1 $display("%b", po);
# 1  pi=13'b0010100100100;
#1 $display("%b", po);
# 1  pi=13'b0010100100101;
#1 $display("%b", po);
# 1  pi=13'b0010100100110;
#1 $display("%b", po);
# 1  pi=13'b0010100100111;
#1 $display("%b", po);
# 1  pi=13'b0010100101000;
#1 $display("%b", po);
# 1  pi=13'b0010100101001;
#1 $display("%b", po);
# 1  pi=13'b0010100101010;
#1 $display("%b", po);
# 1  pi=13'b0010100101011;
#1 $display("%b", po);
# 1  pi=13'b0010100101100;
#1 $display("%b", po);
# 1  pi=13'b0010100101101;
#1 $display("%b", po);
# 1  pi=13'b0010100101110;
#1 $display("%b", po);
# 1  pi=13'b0010100101111;
#1 $display("%b", po);
# 1  pi=13'b0010100110000;
#1 $display("%b", po);
# 1  pi=13'b0010100110001;
#1 $display("%b", po);
# 1  pi=13'b0010100110010;
#1 $display("%b", po);
# 1  pi=13'b0010100110011;
#1 $display("%b", po);
# 1  pi=13'b0010100110100;
#1 $display("%b", po);
# 1  pi=13'b0010100110101;
#1 $display("%b", po);
# 1  pi=13'b0010100110110;
#1 $display("%b", po);
# 1  pi=13'b0010100110111;
#1 $display("%b", po);
# 1  pi=13'b0010100111000;
#1 $display("%b", po);
# 1  pi=13'b0010100111001;
#1 $display("%b", po);
# 1  pi=13'b0010100111010;
#1 $display("%b", po);
# 1  pi=13'b0010100111011;
#1 $display("%b", po);
# 1  pi=13'b0010100111100;
#1 $display("%b", po);
# 1  pi=13'b0010100111101;
#1 $display("%b", po);
# 1  pi=13'b0010100111110;
#1 $display("%b", po);
# 1  pi=13'b0010100111111;
#1 $display("%b", po);
# 1  pi=13'b0010101000000;
#1 $display("%b", po);
# 1  pi=13'b0010101000001;
#1 $display("%b", po);
# 1  pi=13'b0010101000010;
#1 $display("%b", po);
# 1  pi=13'b0010101000011;
#1 $display("%b", po);
# 1  pi=13'b0010101000100;
#1 $display("%b", po);
# 1  pi=13'b0010101000101;
#1 $display("%b", po);
# 1  pi=13'b0010101000110;
#1 $display("%b", po);
# 1  pi=13'b0010101000111;
#1 $display("%b", po);
# 1  pi=13'b0010101001000;
#1 $display("%b", po);
# 1  pi=13'b0010101001001;
#1 $display("%b", po);
# 1  pi=13'b0010101001010;
#1 $display("%b", po);
# 1  pi=13'b0010101001011;
#1 $display("%b", po);
# 1  pi=13'b0010101001100;
#1 $display("%b", po);
# 1  pi=13'b0010101001101;
#1 $display("%b", po);
# 1  pi=13'b0010101001110;
#1 $display("%b", po);
# 1  pi=13'b0010101001111;
#1 $display("%b", po);
# 1  pi=13'b0010101010000;
#1 $display("%b", po);
# 1  pi=13'b0010101010001;
#1 $display("%b", po);
# 1  pi=13'b0010101010010;
#1 $display("%b", po);
# 1  pi=13'b0010101010011;
#1 $display("%b", po);
# 1  pi=13'b0010101010100;
#1 $display("%b", po);
# 1  pi=13'b0010101010101;
#1 $display("%b", po);
# 1  pi=13'b0010101010110;
#1 $display("%b", po);
# 1  pi=13'b0010101010111;
#1 $display("%b", po);
# 1  pi=13'b0010101011000;
#1 $display("%b", po);
# 1  pi=13'b0010101011001;
#1 $display("%b", po);
# 1  pi=13'b0010101011010;
#1 $display("%b", po);
# 1  pi=13'b0010101011011;
#1 $display("%b", po);
# 1  pi=13'b0010101011100;
#1 $display("%b", po);
# 1  pi=13'b0010101011101;
#1 $display("%b", po);
# 1  pi=13'b0010101011110;
#1 $display("%b", po);
# 1  pi=13'b0010101011111;
#1 $display("%b", po);
# 1  pi=13'b0010101100000;
#1 $display("%b", po);
# 1  pi=13'b0010101100001;
#1 $display("%b", po);
# 1  pi=13'b0010101100010;
#1 $display("%b", po);
# 1  pi=13'b0010101100011;
#1 $display("%b", po);
# 1  pi=13'b0010101100100;
#1 $display("%b", po);
# 1  pi=13'b0010101100101;
#1 $display("%b", po);
# 1  pi=13'b0010101100110;
#1 $display("%b", po);
# 1  pi=13'b0010101100111;
#1 $display("%b", po);
# 1  pi=13'b0010101101000;
#1 $display("%b", po);
# 1  pi=13'b0010101101001;
#1 $display("%b", po);
# 1  pi=13'b0010101101010;
#1 $display("%b", po);
# 1  pi=13'b0010101101011;
#1 $display("%b", po);
# 1  pi=13'b0010101101100;
#1 $display("%b", po);
# 1  pi=13'b0010101101101;
#1 $display("%b", po);
# 1  pi=13'b0010101101110;
#1 $display("%b", po);
# 1  pi=13'b0010101101111;
#1 $display("%b", po);
# 1  pi=13'b0010101110000;
#1 $display("%b", po);
# 1  pi=13'b0010101110001;
#1 $display("%b", po);
# 1  pi=13'b0010101110010;
#1 $display("%b", po);
# 1  pi=13'b0010101110011;
#1 $display("%b", po);
# 1  pi=13'b0010101110100;
#1 $display("%b", po);
# 1  pi=13'b0010101110101;
#1 $display("%b", po);
# 1  pi=13'b0010101110110;
#1 $display("%b", po);
# 1  pi=13'b0010101110111;
#1 $display("%b", po);
# 1  pi=13'b0010101111000;
#1 $display("%b", po);
# 1  pi=13'b0010101111001;
#1 $display("%b", po);
# 1  pi=13'b0010101111010;
#1 $display("%b", po);
# 1  pi=13'b0010101111011;
#1 $display("%b", po);
# 1  pi=13'b0010101111100;
#1 $display("%b", po);
# 1  pi=13'b0010101111101;
#1 $display("%b", po);
# 1  pi=13'b0010101111110;
#1 $display("%b", po);
# 1  pi=13'b0010101111111;
#1 $display("%b", po);
# 1  pi=13'b0010110000000;
#1 $display("%b", po);
# 1  pi=13'b0010110000001;
#1 $display("%b", po);
# 1  pi=13'b0010110000010;
#1 $display("%b", po);
# 1  pi=13'b0010110000011;
#1 $display("%b", po);
# 1  pi=13'b0010110000100;
#1 $display("%b", po);
# 1  pi=13'b0010110000101;
#1 $display("%b", po);
# 1  pi=13'b0010110000110;
#1 $display("%b", po);
# 1  pi=13'b0010110000111;
#1 $display("%b", po);
# 1  pi=13'b0010110001000;
#1 $display("%b", po);
# 1  pi=13'b0010110001001;
#1 $display("%b", po);
# 1  pi=13'b0010110001010;
#1 $display("%b", po);
# 1  pi=13'b0010110001011;
#1 $display("%b", po);
# 1  pi=13'b0010110001100;
#1 $display("%b", po);
# 1  pi=13'b0010110001101;
#1 $display("%b", po);
# 1  pi=13'b0010110001110;
#1 $display("%b", po);
# 1  pi=13'b0010110001111;
#1 $display("%b", po);
# 1  pi=13'b0010110010000;
#1 $display("%b", po);
# 1  pi=13'b0010110010001;
#1 $display("%b", po);
# 1  pi=13'b0010110010010;
#1 $display("%b", po);
# 1  pi=13'b0010110010011;
#1 $display("%b", po);
# 1  pi=13'b0010110010100;
#1 $display("%b", po);
# 1  pi=13'b0010110010101;
#1 $display("%b", po);
# 1  pi=13'b0010110010110;
#1 $display("%b", po);
# 1  pi=13'b0010110010111;
#1 $display("%b", po);
# 1  pi=13'b0010110011000;
#1 $display("%b", po);
# 1  pi=13'b0010110011001;
#1 $display("%b", po);
# 1  pi=13'b0010110011010;
#1 $display("%b", po);
# 1  pi=13'b0010110011011;
#1 $display("%b", po);
# 1  pi=13'b0010110011100;
#1 $display("%b", po);
# 1  pi=13'b0010110011101;
#1 $display("%b", po);
# 1  pi=13'b0010110011110;
#1 $display("%b", po);
# 1  pi=13'b0010110011111;
#1 $display("%b", po);
# 1  pi=13'b0010110100000;
#1 $display("%b", po);
# 1  pi=13'b0010110100001;
#1 $display("%b", po);
# 1  pi=13'b0010110100010;
#1 $display("%b", po);
# 1  pi=13'b0010110100011;
#1 $display("%b", po);
# 1  pi=13'b0010110100100;
#1 $display("%b", po);
# 1  pi=13'b0010110100101;
#1 $display("%b", po);
# 1  pi=13'b0010110100110;
#1 $display("%b", po);
# 1  pi=13'b0010110100111;
#1 $display("%b", po);
# 1  pi=13'b0010110101000;
#1 $display("%b", po);
# 1  pi=13'b0010110101001;
#1 $display("%b", po);
# 1  pi=13'b0010110101010;
#1 $display("%b", po);
# 1  pi=13'b0010110101011;
#1 $display("%b", po);
# 1  pi=13'b0010110101100;
#1 $display("%b", po);
# 1  pi=13'b0010110101101;
#1 $display("%b", po);
# 1  pi=13'b0010110101110;
#1 $display("%b", po);
# 1  pi=13'b0010110101111;
#1 $display("%b", po);
# 1  pi=13'b0010110110000;
#1 $display("%b", po);
# 1  pi=13'b0010110110001;
#1 $display("%b", po);
# 1  pi=13'b0010110110010;
#1 $display("%b", po);
# 1  pi=13'b0010110110011;
#1 $display("%b", po);
# 1  pi=13'b0010110110100;
#1 $display("%b", po);
# 1  pi=13'b0010110110101;
#1 $display("%b", po);
# 1  pi=13'b0010110110110;
#1 $display("%b", po);
# 1  pi=13'b0010110110111;
#1 $display("%b", po);
# 1  pi=13'b0010110111000;
#1 $display("%b", po);
# 1  pi=13'b0010110111001;
#1 $display("%b", po);
# 1  pi=13'b0010110111010;
#1 $display("%b", po);
# 1  pi=13'b0010110111011;
#1 $display("%b", po);
# 1  pi=13'b0010110111100;
#1 $display("%b", po);
# 1  pi=13'b0010110111101;
#1 $display("%b", po);
# 1  pi=13'b0010110111110;
#1 $display("%b", po);
# 1  pi=13'b0010110111111;
#1 $display("%b", po);
# 1  pi=13'b0010111000000;
#1 $display("%b", po);
# 1  pi=13'b0010111000001;
#1 $display("%b", po);
# 1  pi=13'b0010111000010;
#1 $display("%b", po);
# 1  pi=13'b0010111000011;
#1 $display("%b", po);
# 1  pi=13'b0010111000100;
#1 $display("%b", po);
# 1  pi=13'b0010111000101;
#1 $display("%b", po);
# 1  pi=13'b0010111000110;
#1 $display("%b", po);
# 1  pi=13'b0010111000111;
#1 $display("%b", po);
# 1  pi=13'b0010111001000;
#1 $display("%b", po);
# 1  pi=13'b0010111001001;
#1 $display("%b", po);
# 1  pi=13'b0010111001010;
#1 $display("%b", po);
# 1  pi=13'b0010111001011;
#1 $display("%b", po);
# 1  pi=13'b0010111001100;
#1 $display("%b", po);
# 1  pi=13'b0010111001101;
#1 $display("%b", po);
# 1  pi=13'b0010111001110;
#1 $display("%b", po);
# 1  pi=13'b0010111001111;
#1 $display("%b", po);
# 1  pi=13'b0010111010000;
#1 $display("%b", po);
# 1  pi=13'b0010111010001;
#1 $display("%b", po);
# 1  pi=13'b0010111010010;
#1 $display("%b", po);
# 1  pi=13'b0010111010011;
#1 $display("%b", po);
# 1  pi=13'b0010111010100;
#1 $display("%b", po);
# 1  pi=13'b0010111010101;
#1 $display("%b", po);
# 1  pi=13'b0010111010110;
#1 $display("%b", po);
# 1  pi=13'b0010111010111;
#1 $display("%b", po);
# 1  pi=13'b0010111011000;
#1 $display("%b", po);
# 1  pi=13'b0010111011001;
#1 $display("%b", po);
# 1  pi=13'b0010111011010;
#1 $display("%b", po);
# 1  pi=13'b0010111011011;
#1 $display("%b", po);
# 1  pi=13'b0010111011100;
#1 $display("%b", po);
# 1  pi=13'b0010111011101;
#1 $display("%b", po);
# 1  pi=13'b0010111011110;
#1 $display("%b", po);
# 1  pi=13'b0010111011111;
#1 $display("%b", po);
# 1  pi=13'b0010111100000;
#1 $display("%b", po);
# 1  pi=13'b0010111100001;
#1 $display("%b", po);
# 1  pi=13'b0010111100010;
#1 $display("%b", po);
# 1  pi=13'b0010111100011;
#1 $display("%b", po);
# 1  pi=13'b0010111100100;
#1 $display("%b", po);
# 1  pi=13'b0010111100101;
#1 $display("%b", po);
# 1  pi=13'b0010111100110;
#1 $display("%b", po);
# 1  pi=13'b0010111100111;
#1 $display("%b", po);
# 1  pi=13'b0010111101000;
#1 $display("%b", po);
# 1  pi=13'b0010111101001;
#1 $display("%b", po);
# 1  pi=13'b0010111101010;
#1 $display("%b", po);
# 1  pi=13'b0010111101011;
#1 $display("%b", po);
# 1  pi=13'b0010111101100;
#1 $display("%b", po);
# 1  pi=13'b0010111101101;
#1 $display("%b", po);
# 1  pi=13'b0010111101110;
#1 $display("%b", po);
# 1  pi=13'b0010111101111;
#1 $display("%b", po);
# 1  pi=13'b0010111110000;
#1 $display("%b", po);
# 1  pi=13'b0010111110001;
#1 $display("%b", po);
# 1  pi=13'b0010111110010;
#1 $display("%b", po);
# 1  pi=13'b0010111110011;
#1 $display("%b", po);
# 1  pi=13'b0010111110100;
#1 $display("%b", po);
# 1  pi=13'b0010111110101;
#1 $display("%b", po);
# 1  pi=13'b0010111110110;
#1 $display("%b", po);
# 1  pi=13'b0010111110111;
#1 $display("%b", po);
# 1  pi=13'b0010111111000;
#1 $display("%b", po);
# 1  pi=13'b0010111111001;
#1 $display("%b", po);
# 1  pi=13'b0010111111010;
#1 $display("%b", po);
# 1  pi=13'b0010111111011;
#1 $display("%b", po);
# 1  pi=13'b0010111111100;
#1 $display("%b", po);
# 1  pi=13'b0010111111101;
#1 $display("%b", po);
# 1  pi=13'b0010111111110;
#1 $display("%b", po);
# 1  pi=13'b0010111111111;
#1 $display("%b", po);
# 1  pi=13'b0011000000000;
#1 $display("%b", po);
# 1  pi=13'b0011000000001;
#1 $display("%b", po);
# 1  pi=13'b0011000000010;
#1 $display("%b", po);
# 1  pi=13'b0011000000011;
#1 $display("%b", po);
# 1  pi=13'b0011000000100;
#1 $display("%b", po);
# 1  pi=13'b0011000000101;
#1 $display("%b", po);
# 1  pi=13'b0011000000110;
#1 $display("%b", po);
# 1  pi=13'b0011000000111;
#1 $display("%b", po);
# 1  pi=13'b0011000001000;
#1 $display("%b", po);
# 1  pi=13'b0011000001001;
#1 $display("%b", po);
# 1  pi=13'b0011000001010;
#1 $display("%b", po);
# 1  pi=13'b0011000001011;
#1 $display("%b", po);
# 1  pi=13'b0011000001100;
#1 $display("%b", po);
# 1  pi=13'b0011000001101;
#1 $display("%b", po);
# 1  pi=13'b0011000001110;
#1 $display("%b", po);
# 1  pi=13'b0011000001111;
#1 $display("%b", po);
# 1  pi=13'b0011000010000;
#1 $display("%b", po);
# 1  pi=13'b0011000010001;
#1 $display("%b", po);
# 1  pi=13'b0011000010010;
#1 $display("%b", po);
# 1  pi=13'b0011000010011;
#1 $display("%b", po);
# 1  pi=13'b0011000010100;
#1 $display("%b", po);
# 1  pi=13'b0011000010101;
#1 $display("%b", po);
# 1  pi=13'b0011000010110;
#1 $display("%b", po);
# 1  pi=13'b0011000010111;
#1 $display("%b", po);
# 1  pi=13'b0011000011000;
#1 $display("%b", po);
# 1  pi=13'b0011000011001;
#1 $display("%b", po);
# 1  pi=13'b0011000011010;
#1 $display("%b", po);
# 1  pi=13'b0011000011011;
#1 $display("%b", po);
# 1  pi=13'b0011000011100;
#1 $display("%b", po);
# 1  pi=13'b0011000011101;
#1 $display("%b", po);
# 1  pi=13'b0011000011110;
#1 $display("%b", po);
# 1  pi=13'b0011000011111;
#1 $display("%b", po);
# 1  pi=13'b0011000100000;
#1 $display("%b", po);
# 1  pi=13'b0011000100001;
#1 $display("%b", po);
# 1  pi=13'b0011000100010;
#1 $display("%b", po);
# 1  pi=13'b0011000100011;
#1 $display("%b", po);
# 1  pi=13'b0011000100100;
#1 $display("%b", po);
# 1  pi=13'b0011000100101;
#1 $display("%b", po);
# 1  pi=13'b0011000100110;
#1 $display("%b", po);
# 1  pi=13'b0011000100111;
#1 $display("%b", po);
# 1  pi=13'b0011000101000;
#1 $display("%b", po);
# 1  pi=13'b0011000101001;
#1 $display("%b", po);
# 1  pi=13'b0011000101010;
#1 $display("%b", po);
# 1  pi=13'b0011000101011;
#1 $display("%b", po);
# 1  pi=13'b0011000101100;
#1 $display("%b", po);
# 1  pi=13'b0011000101101;
#1 $display("%b", po);
# 1  pi=13'b0011000101110;
#1 $display("%b", po);
# 1  pi=13'b0011000101111;
#1 $display("%b", po);
# 1  pi=13'b0011000110000;
#1 $display("%b", po);
# 1  pi=13'b0011000110001;
#1 $display("%b", po);
# 1  pi=13'b0011000110010;
#1 $display("%b", po);
# 1  pi=13'b0011000110011;
#1 $display("%b", po);
# 1  pi=13'b0011000110100;
#1 $display("%b", po);
# 1  pi=13'b0011000110101;
#1 $display("%b", po);
# 1  pi=13'b0011000110110;
#1 $display("%b", po);
# 1  pi=13'b0011000110111;
#1 $display("%b", po);
# 1  pi=13'b0011000111000;
#1 $display("%b", po);
# 1  pi=13'b0011000111001;
#1 $display("%b", po);
# 1  pi=13'b0011000111010;
#1 $display("%b", po);
# 1  pi=13'b0011000111011;
#1 $display("%b", po);
# 1  pi=13'b0011000111100;
#1 $display("%b", po);
# 1  pi=13'b0011000111101;
#1 $display("%b", po);
# 1  pi=13'b0011000111110;
#1 $display("%b", po);
# 1  pi=13'b0011000111111;
#1 $display("%b", po);
# 1  pi=13'b0011001000000;
#1 $display("%b", po);
# 1  pi=13'b0011001000001;
#1 $display("%b", po);
# 1  pi=13'b0011001000010;
#1 $display("%b", po);
# 1  pi=13'b0011001000011;
#1 $display("%b", po);
# 1  pi=13'b0011001000100;
#1 $display("%b", po);
# 1  pi=13'b0011001000101;
#1 $display("%b", po);
# 1  pi=13'b0011001000110;
#1 $display("%b", po);
# 1  pi=13'b0011001000111;
#1 $display("%b", po);
# 1  pi=13'b0011001001000;
#1 $display("%b", po);
# 1  pi=13'b0011001001001;
#1 $display("%b", po);
# 1  pi=13'b0011001001010;
#1 $display("%b", po);
# 1  pi=13'b0011001001011;
#1 $display("%b", po);
# 1  pi=13'b0011001001100;
#1 $display("%b", po);
# 1  pi=13'b0011001001101;
#1 $display("%b", po);
# 1  pi=13'b0011001001110;
#1 $display("%b", po);
# 1  pi=13'b0011001001111;
#1 $display("%b", po);
# 1  pi=13'b0011001010000;
#1 $display("%b", po);
# 1  pi=13'b0011001010001;
#1 $display("%b", po);
# 1  pi=13'b0011001010010;
#1 $display("%b", po);
# 1  pi=13'b0011001010011;
#1 $display("%b", po);
# 1  pi=13'b0011001010100;
#1 $display("%b", po);
# 1  pi=13'b0011001010101;
#1 $display("%b", po);
# 1  pi=13'b0011001010110;
#1 $display("%b", po);
# 1  pi=13'b0011001010111;
#1 $display("%b", po);
# 1  pi=13'b0011001011000;
#1 $display("%b", po);
# 1  pi=13'b0011001011001;
#1 $display("%b", po);
# 1  pi=13'b0011001011010;
#1 $display("%b", po);
# 1  pi=13'b0011001011011;
#1 $display("%b", po);
# 1  pi=13'b0011001011100;
#1 $display("%b", po);
# 1  pi=13'b0011001011101;
#1 $display("%b", po);
# 1  pi=13'b0011001011110;
#1 $display("%b", po);
# 1  pi=13'b0011001011111;
#1 $display("%b", po);
# 1  pi=13'b0011001100000;
#1 $display("%b", po);
# 1  pi=13'b0011001100001;
#1 $display("%b", po);
# 1  pi=13'b0011001100010;
#1 $display("%b", po);
# 1  pi=13'b0011001100011;
#1 $display("%b", po);
# 1  pi=13'b0011001100100;
#1 $display("%b", po);
# 1  pi=13'b0011001100101;
#1 $display("%b", po);
# 1  pi=13'b0011001100110;
#1 $display("%b", po);
# 1  pi=13'b0011001100111;
#1 $display("%b", po);
# 1  pi=13'b0011001101000;
#1 $display("%b", po);
# 1  pi=13'b0011001101001;
#1 $display("%b", po);
# 1  pi=13'b0011001101010;
#1 $display("%b", po);
# 1  pi=13'b0011001101011;
#1 $display("%b", po);
# 1  pi=13'b0011001101100;
#1 $display("%b", po);
# 1  pi=13'b0011001101101;
#1 $display("%b", po);
# 1  pi=13'b0011001101110;
#1 $display("%b", po);
# 1  pi=13'b0011001101111;
#1 $display("%b", po);
# 1  pi=13'b0011001110000;
#1 $display("%b", po);
# 1  pi=13'b0011001110001;
#1 $display("%b", po);
# 1  pi=13'b0011001110010;
#1 $display("%b", po);
# 1  pi=13'b0011001110011;
#1 $display("%b", po);
# 1  pi=13'b0011001110100;
#1 $display("%b", po);
# 1  pi=13'b0011001110101;
#1 $display("%b", po);
# 1  pi=13'b0011001110110;
#1 $display("%b", po);
# 1  pi=13'b0011001110111;
#1 $display("%b", po);
# 1  pi=13'b0011001111000;
#1 $display("%b", po);
# 1  pi=13'b0011001111001;
#1 $display("%b", po);
# 1  pi=13'b0011001111010;
#1 $display("%b", po);
# 1  pi=13'b0011001111011;
#1 $display("%b", po);
# 1  pi=13'b0011001111100;
#1 $display("%b", po);
# 1  pi=13'b0011001111101;
#1 $display("%b", po);
# 1  pi=13'b0011001111110;
#1 $display("%b", po);
# 1  pi=13'b0011001111111;
#1 $display("%b", po);
# 1  pi=13'b0011010000000;
#1 $display("%b", po);
# 1  pi=13'b0011010000001;
#1 $display("%b", po);
# 1  pi=13'b0011010000010;
#1 $display("%b", po);
# 1  pi=13'b0011010000011;
#1 $display("%b", po);
# 1  pi=13'b0011010000100;
#1 $display("%b", po);
# 1  pi=13'b0011010000101;
#1 $display("%b", po);
# 1  pi=13'b0011010000110;
#1 $display("%b", po);
# 1  pi=13'b0011010000111;
#1 $display("%b", po);
# 1  pi=13'b0011010001000;
#1 $display("%b", po);
# 1  pi=13'b0011010001001;
#1 $display("%b", po);
# 1  pi=13'b0011010001010;
#1 $display("%b", po);
# 1  pi=13'b0011010001011;
#1 $display("%b", po);
# 1  pi=13'b0011010001100;
#1 $display("%b", po);
# 1  pi=13'b0011010001101;
#1 $display("%b", po);
# 1  pi=13'b0011010001110;
#1 $display("%b", po);
# 1  pi=13'b0011010001111;
#1 $display("%b", po);
# 1  pi=13'b0011010010000;
#1 $display("%b", po);
# 1  pi=13'b0011010010001;
#1 $display("%b", po);
# 1  pi=13'b0011010010010;
#1 $display("%b", po);
# 1  pi=13'b0011010010011;
#1 $display("%b", po);
# 1  pi=13'b0011010010100;
#1 $display("%b", po);
# 1  pi=13'b0011010010101;
#1 $display("%b", po);
# 1  pi=13'b0011010010110;
#1 $display("%b", po);
# 1  pi=13'b0011010010111;
#1 $display("%b", po);
# 1  pi=13'b0011010011000;
#1 $display("%b", po);
# 1  pi=13'b0011010011001;
#1 $display("%b", po);
# 1  pi=13'b0011010011010;
#1 $display("%b", po);
# 1  pi=13'b0011010011011;
#1 $display("%b", po);
# 1  pi=13'b0011010011100;
#1 $display("%b", po);
# 1  pi=13'b0011010011101;
#1 $display("%b", po);
# 1  pi=13'b0011010011110;
#1 $display("%b", po);
# 1  pi=13'b0011010011111;
#1 $display("%b", po);
# 1  pi=13'b0011010100000;
#1 $display("%b", po);
# 1  pi=13'b0011010100001;
#1 $display("%b", po);
# 1  pi=13'b0011010100010;
#1 $display("%b", po);
# 1  pi=13'b0011010100011;
#1 $display("%b", po);
# 1  pi=13'b0011010100100;
#1 $display("%b", po);
# 1  pi=13'b0011010100101;
#1 $display("%b", po);
# 1  pi=13'b0011010100110;
#1 $display("%b", po);
# 1  pi=13'b0011010100111;
#1 $display("%b", po);
# 1  pi=13'b0011010101000;
#1 $display("%b", po);
# 1  pi=13'b0011010101001;
#1 $display("%b", po);
# 1  pi=13'b0011010101010;
#1 $display("%b", po);
# 1  pi=13'b0011010101011;
#1 $display("%b", po);
# 1  pi=13'b0011010101100;
#1 $display("%b", po);
# 1  pi=13'b0011010101101;
#1 $display("%b", po);
# 1  pi=13'b0011010101110;
#1 $display("%b", po);
# 1  pi=13'b0011010101111;
#1 $display("%b", po);
# 1  pi=13'b0011010110000;
#1 $display("%b", po);
# 1  pi=13'b0011010110001;
#1 $display("%b", po);
# 1  pi=13'b0011010110010;
#1 $display("%b", po);
# 1  pi=13'b0011010110011;
#1 $display("%b", po);
# 1  pi=13'b0011010110100;
#1 $display("%b", po);
# 1  pi=13'b0011010110101;
#1 $display("%b", po);
# 1  pi=13'b0011010110110;
#1 $display("%b", po);
# 1  pi=13'b0011010110111;
#1 $display("%b", po);
# 1  pi=13'b0011010111000;
#1 $display("%b", po);
# 1  pi=13'b0011010111001;
#1 $display("%b", po);
# 1  pi=13'b0011010111010;
#1 $display("%b", po);
# 1  pi=13'b0011010111011;
#1 $display("%b", po);
# 1  pi=13'b0011010111100;
#1 $display("%b", po);
# 1  pi=13'b0011010111101;
#1 $display("%b", po);
# 1  pi=13'b0011010111110;
#1 $display("%b", po);
# 1  pi=13'b0011010111111;
#1 $display("%b", po);
# 1  pi=13'b0011011000000;
#1 $display("%b", po);
# 1  pi=13'b0011011000001;
#1 $display("%b", po);
# 1  pi=13'b0011011000010;
#1 $display("%b", po);
# 1  pi=13'b0011011000011;
#1 $display("%b", po);
# 1  pi=13'b0011011000100;
#1 $display("%b", po);
# 1  pi=13'b0011011000101;
#1 $display("%b", po);
# 1  pi=13'b0011011000110;
#1 $display("%b", po);
# 1  pi=13'b0011011000111;
#1 $display("%b", po);
# 1  pi=13'b0011011001000;
#1 $display("%b", po);
# 1  pi=13'b0011011001001;
#1 $display("%b", po);
# 1  pi=13'b0011011001010;
#1 $display("%b", po);
# 1  pi=13'b0011011001011;
#1 $display("%b", po);
# 1  pi=13'b0011011001100;
#1 $display("%b", po);
# 1  pi=13'b0011011001101;
#1 $display("%b", po);
# 1  pi=13'b0011011001110;
#1 $display("%b", po);
# 1  pi=13'b0011011001111;
#1 $display("%b", po);
# 1  pi=13'b0011011010000;
#1 $display("%b", po);
# 1  pi=13'b0011011010001;
#1 $display("%b", po);
# 1  pi=13'b0011011010010;
#1 $display("%b", po);
# 1  pi=13'b0011011010011;
#1 $display("%b", po);
# 1  pi=13'b0011011010100;
#1 $display("%b", po);
# 1  pi=13'b0011011010101;
#1 $display("%b", po);
# 1  pi=13'b0011011010110;
#1 $display("%b", po);
# 1  pi=13'b0011011010111;
#1 $display("%b", po);
# 1  pi=13'b0011011011000;
#1 $display("%b", po);
# 1  pi=13'b0011011011001;
#1 $display("%b", po);
# 1  pi=13'b0011011011010;
#1 $display("%b", po);
# 1  pi=13'b0011011011011;
#1 $display("%b", po);
# 1  pi=13'b0011011011100;
#1 $display("%b", po);
# 1  pi=13'b0011011011101;
#1 $display("%b", po);
# 1  pi=13'b0011011011110;
#1 $display("%b", po);
# 1  pi=13'b0011011011111;
#1 $display("%b", po);
# 1  pi=13'b0011011100000;
#1 $display("%b", po);
# 1  pi=13'b0011011100001;
#1 $display("%b", po);
# 1  pi=13'b0011011100010;
#1 $display("%b", po);
# 1  pi=13'b0011011100011;
#1 $display("%b", po);
# 1  pi=13'b0011011100100;
#1 $display("%b", po);
# 1  pi=13'b0011011100101;
#1 $display("%b", po);
# 1  pi=13'b0011011100110;
#1 $display("%b", po);
# 1  pi=13'b0011011100111;
#1 $display("%b", po);
# 1  pi=13'b0011011101000;
#1 $display("%b", po);
# 1  pi=13'b0011011101001;
#1 $display("%b", po);
# 1  pi=13'b0011011101010;
#1 $display("%b", po);
# 1  pi=13'b0011011101011;
#1 $display("%b", po);
# 1  pi=13'b0011011101100;
#1 $display("%b", po);
# 1  pi=13'b0011011101101;
#1 $display("%b", po);
# 1  pi=13'b0011011101110;
#1 $display("%b", po);
# 1  pi=13'b0011011101111;
#1 $display("%b", po);
# 1  pi=13'b0011011110000;
#1 $display("%b", po);
# 1  pi=13'b0011011110001;
#1 $display("%b", po);
# 1  pi=13'b0011011110010;
#1 $display("%b", po);
# 1  pi=13'b0011011110011;
#1 $display("%b", po);
# 1  pi=13'b0011011110100;
#1 $display("%b", po);
# 1  pi=13'b0011011110101;
#1 $display("%b", po);
# 1  pi=13'b0011011110110;
#1 $display("%b", po);
# 1  pi=13'b0011011110111;
#1 $display("%b", po);
# 1  pi=13'b0011011111000;
#1 $display("%b", po);
# 1  pi=13'b0011011111001;
#1 $display("%b", po);
# 1  pi=13'b0011011111010;
#1 $display("%b", po);
# 1  pi=13'b0011011111011;
#1 $display("%b", po);
# 1  pi=13'b0011011111100;
#1 $display("%b", po);
# 1  pi=13'b0011011111101;
#1 $display("%b", po);
# 1  pi=13'b0011011111110;
#1 $display("%b", po);
# 1  pi=13'b0011011111111;
#1 $display("%b", po);
# 1  pi=13'b0011100000000;
#1 $display("%b", po);
# 1  pi=13'b0011100000001;
#1 $display("%b", po);
# 1  pi=13'b0011100000010;
#1 $display("%b", po);
# 1  pi=13'b0011100000011;
#1 $display("%b", po);
# 1  pi=13'b0011100000100;
#1 $display("%b", po);
# 1  pi=13'b0011100000101;
#1 $display("%b", po);
# 1  pi=13'b0011100000110;
#1 $display("%b", po);
# 1  pi=13'b0011100000111;
#1 $display("%b", po);
# 1  pi=13'b0011100001000;
#1 $display("%b", po);
# 1  pi=13'b0011100001001;
#1 $display("%b", po);
# 1  pi=13'b0011100001010;
#1 $display("%b", po);
# 1  pi=13'b0011100001011;
#1 $display("%b", po);
# 1  pi=13'b0011100001100;
#1 $display("%b", po);
# 1  pi=13'b0011100001101;
#1 $display("%b", po);
# 1  pi=13'b0011100001110;
#1 $display("%b", po);
# 1  pi=13'b0011100001111;
#1 $display("%b", po);
# 1  pi=13'b0011100010000;
#1 $display("%b", po);
# 1  pi=13'b0011100010001;
#1 $display("%b", po);
# 1  pi=13'b0011100010010;
#1 $display("%b", po);
# 1  pi=13'b0011100010011;
#1 $display("%b", po);
# 1  pi=13'b0011100010100;
#1 $display("%b", po);
# 1  pi=13'b0011100010101;
#1 $display("%b", po);
# 1  pi=13'b0011100010110;
#1 $display("%b", po);
# 1  pi=13'b0011100010111;
#1 $display("%b", po);
# 1  pi=13'b0011100011000;
#1 $display("%b", po);
# 1  pi=13'b0011100011001;
#1 $display("%b", po);
# 1  pi=13'b0011100011010;
#1 $display("%b", po);
# 1  pi=13'b0011100011011;
#1 $display("%b", po);
# 1  pi=13'b0011100011100;
#1 $display("%b", po);
# 1  pi=13'b0011100011101;
#1 $display("%b", po);
# 1  pi=13'b0011100011110;
#1 $display("%b", po);
# 1  pi=13'b0011100011111;
#1 $display("%b", po);
# 1  pi=13'b0011100100000;
#1 $display("%b", po);
# 1  pi=13'b0011100100001;
#1 $display("%b", po);
# 1  pi=13'b0011100100010;
#1 $display("%b", po);
# 1  pi=13'b0011100100011;
#1 $display("%b", po);
# 1  pi=13'b0011100100100;
#1 $display("%b", po);
# 1  pi=13'b0011100100101;
#1 $display("%b", po);
# 1  pi=13'b0011100100110;
#1 $display("%b", po);
# 1  pi=13'b0011100100111;
#1 $display("%b", po);
# 1  pi=13'b0011100101000;
#1 $display("%b", po);
# 1  pi=13'b0011100101001;
#1 $display("%b", po);
# 1  pi=13'b0011100101010;
#1 $display("%b", po);
# 1  pi=13'b0011100101011;
#1 $display("%b", po);
# 1  pi=13'b0011100101100;
#1 $display("%b", po);
# 1  pi=13'b0011100101101;
#1 $display("%b", po);
# 1  pi=13'b0011100101110;
#1 $display("%b", po);
# 1  pi=13'b0011100101111;
#1 $display("%b", po);
# 1  pi=13'b0011100110000;
#1 $display("%b", po);
# 1  pi=13'b0011100110001;
#1 $display("%b", po);
# 1  pi=13'b0011100110010;
#1 $display("%b", po);
# 1  pi=13'b0011100110011;
#1 $display("%b", po);
# 1  pi=13'b0011100110100;
#1 $display("%b", po);
# 1  pi=13'b0011100110101;
#1 $display("%b", po);
# 1  pi=13'b0011100110110;
#1 $display("%b", po);
# 1  pi=13'b0011100110111;
#1 $display("%b", po);
# 1  pi=13'b0011100111000;
#1 $display("%b", po);
# 1  pi=13'b0011100111001;
#1 $display("%b", po);
# 1  pi=13'b0011100111010;
#1 $display("%b", po);
# 1  pi=13'b0011100111011;
#1 $display("%b", po);
# 1  pi=13'b0011100111100;
#1 $display("%b", po);
# 1  pi=13'b0011100111101;
#1 $display("%b", po);
# 1  pi=13'b0011100111110;
#1 $display("%b", po);
# 1  pi=13'b0011100111111;
#1 $display("%b", po);
# 1  pi=13'b0011101000000;
#1 $display("%b", po);
# 1  pi=13'b0011101000001;
#1 $display("%b", po);
# 1  pi=13'b0011101000010;
#1 $display("%b", po);
# 1  pi=13'b0011101000011;
#1 $display("%b", po);
# 1  pi=13'b0011101000100;
#1 $display("%b", po);
# 1  pi=13'b0011101000101;
#1 $display("%b", po);
# 1  pi=13'b0011101000110;
#1 $display("%b", po);
# 1  pi=13'b0011101000111;
#1 $display("%b", po);
# 1  pi=13'b0011101001000;
#1 $display("%b", po);
# 1  pi=13'b0011101001001;
#1 $display("%b", po);
# 1  pi=13'b0011101001010;
#1 $display("%b", po);
# 1  pi=13'b0011101001011;
#1 $display("%b", po);
# 1  pi=13'b0011101001100;
#1 $display("%b", po);
# 1  pi=13'b0011101001101;
#1 $display("%b", po);
# 1  pi=13'b0011101001110;
#1 $display("%b", po);
# 1  pi=13'b0011101001111;
#1 $display("%b", po);
# 1  pi=13'b0011101010000;
#1 $display("%b", po);
# 1  pi=13'b0011101010001;
#1 $display("%b", po);
# 1  pi=13'b0011101010010;
#1 $display("%b", po);
# 1  pi=13'b0011101010011;
#1 $display("%b", po);
# 1  pi=13'b0011101010100;
#1 $display("%b", po);
# 1  pi=13'b0011101010101;
#1 $display("%b", po);
# 1  pi=13'b0011101010110;
#1 $display("%b", po);
# 1  pi=13'b0011101010111;
#1 $display("%b", po);
# 1  pi=13'b0011101011000;
#1 $display("%b", po);
# 1  pi=13'b0011101011001;
#1 $display("%b", po);
# 1  pi=13'b0011101011010;
#1 $display("%b", po);
# 1  pi=13'b0011101011011;
#1 $display("%b", po);
# 1  pi=13'b0011101011100;
#1 $display("%b", po);
# 1  pi=13'b0011101011101;
#1 $display("%b", po);
# 1  pi=13'b0011101011110;
#1 $display("%b", po);
# 1  pi=13'b0011101011111;
#1 $display("%b", po);
# 1  pi=13'b0011101100000;
#1 $display("%b", po);
# 1  pi=13'b0011101100001;
#1 $display("%b", po);
# 1  pi=13'b0011101100010;
#1 $display("%b", po);
# 1  pi=13'b0011101100011;
#1 $display("%b", po);
# 1  pi=13'b0011101100100;
#1 $display("%b", po);
# 1  pi=13'b0011101100101;
#1 $display("%b", po);
# 1  pi=13'b0011101100110;
#1 $display("%b", po);
# 1  pi=13'b0011101100111;
#1 $display("%b", po);
# 1  pi=13'b0011101101000;
#1 $display("%b", po);
# 1  pi=13'b0011101101001;
#1 $display("%b", po);
# 1  pi=13'b0011101101010;
#1 $display("%b", po);
# 1  pi=13'b0011101101011;
#1 $display("%b", po);
# 1  pi=13'b0011101101100;
#1 $display("%b", po);
# 1  pi=13'b0011101101101;
#1 $display("%b", po);
# 1  pi=13'b0011101101110;
#1 $display("%b", po);
# 1  pi=13'b0011101101111;
#1 $display("%b", po);
# 1  pi=13'b0011101110000;
#1 $display("%b", po);
# 1  pi=13'b0011101110001;
#1 $display("%b", po);
# 1  pi=13'b0011101110010;
#1 $display("%b", po);
# 1  pi=13'b0011101110011;
#1 $display("%b", po);
# 1  pi=13'b0011101110100;
#1 $display("%b", po);
# 1  pi=13'b0011101110101;
#1 $display("%b", po);
# 1  pi=13'b0011101110110;
#1 $display("%b", po);
# 1  pi=13'b0011101110111;
#1 $display("%b", po);
# 1  pi=13'b0011101111000;
#1 $display("%b", po);
# 1  pi=13'b0011101111001;
#1 $display("%b", po);
# 1  pi=13'b0011101111010;
#1 $display("%b", po);
# 1  pi=13'b0011101111011;
#1 $display("%b", po);
# 1  pi=13'b0011101111100;
#1 $display("%b", po);
# 1  pi=13'b0011101111101;
#1 $display("%b", po);
# 1  pi=13'b0011101111110;
#1 $display("%b", po);
# 1  pi=13'b0011101111111;
#1 $display("%b", po);
# 1  pi=13'b0011110000000;
#1 $display("%b", po);
# 1  pi=13'b0011110000001;
#1 $display("%b", po);
# 1  pi=13'b0011110000010;
#1 $display("%b", po);
# 1  pi=13'b0011110000011;
#1 $display("%b", po);
# 1  pi=13'b0011110000100;
#1 $display("%b", po);
# 1  pi=13'b0011110000101;
#1 $display("%b", po);
# 1  pi=13'b0011110000110;
#1 $display("%b", po);
# 1  pi=13'b0011110000111;
#1 $display("%b", po);
# 1  pi=13'b0011110001000;
#1 $display("%b", po);
# 1  pi=13'b0011110001001;
#1 $display("%b", po);
# 1  pi=13'b0011110001010;
#1 $display("%b", po);
# 1  pi=13'b0011110001011;
#1 $display("%b", po);
# 1  pi=13'b0011110001100;
#1 $display("%b", po);
# 1  pi=13'b0011110001101;
#1 $display("%b", po);
# 1  pi=13'b0011110001110;
#1 $display("%b", po);
# 1  pi=13'b0011110001111;
#1 $display("%b", po);
# 1  pi=13'b0011110010000;
#1 $display("%b", po);
# 1  pi=13'b0011110010001;
#1 $display("%b", po);
# 1  pi=13'b0011110010010;
#1 $display("%b", po);
# 1  pi=13'b0011110010011;
#1 $display("%b", po);
# 1  pi=13'b0011110010100;
#1 $display("%b", po);
# 1  pi=13'b0011110010101;
#1 $display("%b", po);
# 1  pi=13'b0011110010110;
#1 $display("%b", po);
# 1  pi=13'b0011110010111;
#1 $display("%b", po);
# 1  pi=13'b0011110011000;
#1 $display("%b", po);
# 1  pi=13'b0011110011001;
#1 $display("%b", po);
# 1  pi=13'b0011110011010;
#1 $display("%b", po);
# 1  pi=13'b0011110011011;
#1 $display("%b", po);
# 1  pi=13'b0011110011100;
#1 $display("%b", po);
# 1  pi=13'b0011110011101;
#1 $display("%b", po);
# 1  pi=13'b0011110011110;
#1 $display("%b", po);
# 1  pi=13'b0011110011111;
#1 $display("%b", po);
# 1  pi=13'b0011110100000;
#1 $display("%b", po);
# 1  pi=13'b0011110100001;
#1 $display("%b", po);
# 1  pi=13'b0011110100010;
#1 $display("%b", po);
# 1  pi=13'b0011110100011;
#1 $display("%b", po);
# 1  pi=13'b0011110100100;
#1 $display("%b", po);
# 1  pi=13'b0011110100101;
#1 $display("%b", po);
# 1  pi=13'b0011110100110;
#1 $display("%b", po);
# 1  pi=13'b0011110100111;
#1 $display("%b", po);
# 1  pi=13'b0011110101000;
#1 $display("%b", po);
# 1  pi=13'b0011110101001;
#1 $display("%b", po);
# 1  pi=13'b0011110101010;
#1 $display("%b", po);
# 1  pi=13'b0011110101011;
#1 $display("%b", po);
# 1  pi=13'b0011110101100;
#1 $display("%b", po);
# 1  pi=13'b0011110101101;
#1 $display("%b", po);
# 1  pi=13'b0011110101110;
#1 $display("%b", po);
# 1  pi=13'b0011110101111;
#1 $display("%b", po);
# 1  pi=13'b0011110110000;
#1 $display("%b", po);
# 1  pi=13'b0011110110001;
#1 $display("%b", po);
# 1  pi=13'b0011110110010;
#1 $display("%b", po);
# 1  pi=13'b0011110110011;
#1 $display("%b", po);
# 1  pi=13'b0011110110100;
#1 $display("%b", po);
# 1  pi=13'b0011110110101;
#1 $display("%b", po);
# 1  pi=13'b0011110110110;
#1 $display("%b", po);
# 1  pi=13'b0011110110111;
#1 $display("%b", po);
# 1  pi=13'b0011110111000;
#1 $display("%b", po);
# 1  pi=13'b0011110111001;
#1 $display("%b", po);
# 1  pi=13'b0011110111010;
#1 $display("%b", po);
# 1  pi=13'b0011110111011;
#1 $display("%b", po);
# 1  pi=13'b0011110111100;
#1 $display("%b", po);
# 1  pi=13'b0011110111101;
#1 $display("%b", po);
# 1  pi=13'b0011110111110;
#1 $display("%b", po);
# 1  pi=13'b0011110111111;
#1 $display("%b", po);
# 1  pi=13'b0011111000000;
#1 $display("%b", po);
# 1  pi=13'b0011111000001;
#1 $display("%b", po);
# 1  pi=13'b0011111000010;
#1 $display("%b", po);
# 1  pi=13'b0011111000011;
#1 $display("%b", po);
# 1  pi=13'b0011111000100;
#1 $display("%b", po);
# 1  pi=13'b0011111000101;
#1 $display("%b", po);
# 1  pi=13'b0011111000110;
#1 $display("%b", po);
# 1  pi=13'b0011111000111;
#1 $display("%b", po);
# 1  pi=13'b0011111001000;
#1 $display("%b", po);
# 1  pi=13'b0011111001001;
#1 $display("%b", po);
# 1  pi=13'b0011111001010;
#1 $display("%b", po);
# 1  pi=13'b0011111001011;
#1 $display("%b", po);
# 1  pi=13'b0011111001100;
#1 $display("%b", po);
# 1  pi=13'b0011111001101;
#1 $display("%b", po);
# 1  pi=13'b0011111001110;
#1 $display("%b", po);
# 1  pi=13'b0011111001111;
#1 $display("%b", po);
# 1  pi=13'b0011111010000;
#1 $display("%b", po);
# 1  pi=13'b0011111010001;
#1 $display("%b", po);
# 1  pi=13'b0011111010010;
#1 $display("%b", po);
# 1  pi=13'b0011111010011;
#1 $display("%b", po);
# 1  pi=13'b0011111010100;
#1 $display("%b", po);
# 1  pi=13'b0011111010101;
#1 $display("%b", po);
# 1  pi=13'b0011111010110;
#1 $display("%b", po);
# 1  pi=13'b0011111010111;
#1 $display("%b", po);
# 1  pi=13'b0011111011000;
#1 $display("%b", po);
# 1  pi=13'b0011111011001;
#1 $display("%b", po);
# 1  pi=13'b0011111011010;
#1 $display("%b", po);
# 1  pi=13'b0011111011011;
#1 $display("%b", po);
# 1  pi=13'b0011111011100;
#1 $display("%b", po);
# 1  pi=13'b0011111011101;
#1 $display("%b", po);
# 1  pi=13'b0011111011110;
#1 $display("%b", po);
# 1  pi=13'b0011111011111;
#1 $display("%b", po);
# 1  pi=13'b0011111100000;
#1 $display("%b", po);
# 1  pi=13'b0011111100001;
#1 $display("%b", po);
# 1  pi=13'b0011111100010;
#1 $display("%b", po);
# 1  pi=13'b0011111100011;
#1 $display("%b", po);
# 1  pi=13'b0011111100100;
#1 $display("%b", po);
# 1  pi=13'b0011111100101;
#1 $display("%b", po);
# 1  pi=13'b0011111100110;
#1 $display("%b", po);
# 1  pi=13'b0011111100111;
#1 $display("%b", po);
# 1  pi=13'b0011111101000;
#1 $display("%b", po);
# 1  pi=13'b0011111101001;
#1 $display("%b", po);
# 1  pi=13'b0011111101010;
#1 $display("%b", po);
# 1  pi=13'b0011111101011;
#1 $display("%b", po);
# 1  pi=13'b0011111101100;
#1 $display("%b", po);
# 1  pi=13'b0011111101101;
#1 $display("%b", po);
# 1  pi=13'b0011111101110;
#1 $display("%b", po);
# 1  pi=13'b0011111101111;
#1 $display("%b", po);
# 1  pi=13'b0011111110000;
#1 $display("%b", po);
# 1  pi=13'b0011111110001;
#1 $display("%b", po);
# 1  pi=13'b0011111110010;
#1 $display("%b", po);
# 1  pi=13'b0011111110011;
#1 $display("%b", po);
# 1  pi=13'b0011111110100;
#1 $display("%b", po);
# 1  pi=13'b0011111110101;
#1 $display("%b", po);
# 1  pi=13'b0011111110110;
#1 $display("%b", po);
# 1  pi=13'b0011111110111;
#1 $display("%b", po);
# 1  pi=13'b0011111111000;
#1 $display("%b", po);
# 1  pi=13'b0011111111001;
#1 $display("%b", po);
# 1  pi=13'b0011111111010;
#1 $display("%b", po);
# 1  pi=13'b0011111111011;
#1 $display("%b", po);
# 1  pi=13'b0011111111100;
#1 $display("%b", po);
# 1  pi=13'b0011111111101;
#1 $display("%b", po);
# 1  pi=13'b0011111111110;
#1 $display("%b", po);
# 1  pi=13'b0011111111111;
#1 $display("%b", po);
# 1  pi=13'b0100000000000;
#1 $display("%b", po);
# 1  pi=13'b0100000000001;
#1 $display("%b", po);
# 1  pi=13'b0100000000010;
#1 $display("%b", po);
# 1  pi=13'b0100000000011;
#1 $display("%b", po);
# 1  pi=13'b0100000000100;
#1 $display("%b", po);
# 1  pi=13'b0100000000101;
#1 $display("%b", po);
# 1  pi=13'b0100000000110;
#1 $display("%b", po);
# 1  pi=13'b0100000000111;
#1 $display("%b", po);
# 1  pi=13'b0100000001000;
#1 $display("%b", po);
# 1  pi=13'b0100000001001;
#1 $display("%b", po);
# 1  pi=13'b0100000001010;
#1 $display("%b", po);
# 1  pi=13'b0100000001011;
#1 $display("%b", po);
# 1  pi=13'b0100000001100;
#1 $display("%b", po);
# 1  pi=13'b0100000001101;
#1 $display("%b", po);
# 1  pi=13'b0100000001110;
#1 $display("%b", po);
# 1  pi=13'b0100000001111;
#1 $display("%b", po);
# 1  pi=13'b0100000010000;
#1 $display("%b", po);
# 1  pi=13'b0100000010001;
#1 $display("%b", po);
# 1  pi=13'b0100000010010;
#1 $display("%b", po);
# 1  pi=13'b0100000010011;
#1 $display("%b", po);
# 1  pi=13'b0100000010100;
#1 $display("%b", po);
# 1  pi=13'b0100000010101;
#1 $display("%b", po);
# 1  pi=13'b0100000010110;
#1 $display("%b", po);
# 1  pi=13'b0100000010111;
#1 $display("%b", po);
# 1  pi=13'b0100000011000;
#1 $display("%b", po);
# 1  pi=13'b0100000011001;
#1 $display("%b", po);
# 1  pi=13'b0100000011010;
#1 $display("%b", po);
# 1  pi=13'b0100000011011;
#1 $display("%b", po);
# 1  pi=13'b0100000011100;
#1 $display("%b", po);
# 1  pi=13'b0100000011101;
#1 $display("%b", po);
# 1  pi=13'b0100000011110;
#1 $display("%b", po);
# 1  pi=13'b0100000011111;
#1 $display("%b", po);
# 1  pi=13'b0100000100000;
#1 $display("%b", po);
# 1  pi=13'b0100000100001;
#1 $display("%b", po);
# 1  pi=13'b0100000100010;
#1 $display("%b", po);
# 1  pi=13'b0100000100011;
#1 $display("%b", po);
# 1  pi=13'b0100000100100;
#1 $display("%b", po);
# 1  pi=13'b0100000100101;
#1 $display("%b", po);
# 1  pi=13'b0100000100110;
#1 $display("%b", po);
# 1  pi=13'b0100000100111;
#1 $display("%b", po);
# 1  pi=13'b0100000101000;
#1 $display("%b", po);
# 1  pi=13'b0100000101001;
#1 $display("%b", po);
# 1  pi=13'b0100000101010;
#1 $display("%b", po);
# 1  pi=13'b0100000101011;
#1 $display("%b", po);
# 1  pi=13'b0100000101100;
#1 $display("%b", po);
# 1  pi=13'b0100000101101;
#1 $display("%b", po);
# 1  pi=13'b0100000101110;
#1 $display("%b", po);
# 1  pi=13'b0100000101111;
#1 $display("%b", po);
# 1  pi=13'b0100000110000;
#1 $display("%b", po);
# 1  pi=13'b0100000110001;
#1 $display("%b", po);
# 1  pi=13'b0100000110010;
#1 $display("%b", po);
# 1  pi=13'b0100000110011;
#1 $display("%b", po);
# 1  pi=13'b0100000110100;
#1 $display("%b", po);
# 1  pi=13'b0100000110101;
#1 $display("%b", po);
# 1  pi=13'b0100000110110;
#1 $display("%b", po);
# 1  pi=13'b0100000110111;
#1 $display("%b", po);
# 1  pi=13'b0100000111000;
#1 $display("%b", po);
# 1  pi=13'b0100000111001;
#1 $display("%b", po);
# 1  pi=13'b0100000111010;
#1 $display("%b", po);
# 1  pi=13'b0100000111011;
#1 $display("%b", po);
# 1  pi=13'b0100000111100;
#1 $display("%b", po);
# 1  pi=13'b0100000111101;
#1 $display("%b", po);
# 1  pi=13'b0100000111110;
#1 $display("%b", po);
# 1  pi=13'b0100000111111;
#1 $display("%b", po);
# 1  pi=13'b0100001000000;
#1 $display("%b", po);
# 1  pi=13'b0100001000001;
#1 $display("%b", po);
# 1  pi=13'b0100001000010;
#1 $display("%b", po);
# 1  pi=13'b0100001000011;
#1 $display("%b", po);
# 1  pi=13'b0100001000100;
#1 $display("%b", po);
# 1  pi=13'b0100001000101;
#1 $display("%b", po);
# 1  pi=13'b0100001000110;
#1 $display("%b", po);
# 1  pi=13'b0100001000111;
#1 $display("%b", po);
# 1  pi=13'b0100001001000;
#1 $display("%b", po);
# 1  pi=13'b0100001001001;
#1 $display("%b", po);
# 1  pi=13'b0100001001010;
#1 $display("%b", po);
# 1  pi=13'b0100001001011;
#1 $display("%b", po);
# 1  pi=13'b0100001001100;
#1 $display("%b", po);
# 1  pi=13'b0100001001101;
#1 $display("%b", po);
# 1  pi=13'b0100001001110;
#1 $display("%b", po);
# 1  pi=13'b0100001001111;
#1 $display("%b", po);
# 1  pi=13'b0100001010000;
#1 $display("%b", po);
# 1  pi=13'b0100001010001;
#1 $display("%b", po);
# 1  pi=13'b0100001010010;
#1 $display("%b", po);
# 1  pi=13'b0100001010011;
#1 $display("%b", po);
# 1  pi=13'b0100001010100;
#1 $display("%b", po);
# 1  pi=13'b0100001010101;
#1 $display("%b", po);
# 1  pi=13'b0100001010110;
#1 $display("%b", po);
# 1  pi=13'b0100001010111;
#1 $display("%b", po);
# 1  pi=13'b0100001011000;
#1 $display("%b", po);
# 1  pi=13'b0100001011001;
#1 $display("%b", po);
# 1  pi=13'b0100001011010;
#1 $display("%b", po);
# 1  pi=13'b0100001011011;
#1 $display("%b", po);
# 1  pi=13'b0100001011100;
#1 $display("%b", po);
# 1  pi=13'b0100001011101;
#1 $display("%b", po);
# 1  pi=13'b0100001011110;
#1 $display("%b", po);
# 1  pi=13'b0100001011111;
#1 $display("%b", po);
# 1  pi=13'b0100001100000;
#1 $display("%b", po);
# 1  pi=13'b0100001100001;
#1 $display("%b", po);
# 1  pi=13'b0100001100010;
#1 $display("%b", po);
# 1  pi=13'b0100001100011;
#1 $display("%b", po);
# 1  pi=13'b0100001100100;
#1 $display("%b", po);
# 1  pi=13'b0100001100101;
#1 $display("%b", po);
# 1  pi=13'b0100001100110;
#1 $display("%b", po);
# 1  pi=13'b0100001100111;
#1 $display("%b", po);
# 1  pi=13'b0100001101000;
#1 $display("%b", po);
# 1  pi=13'b0100001101001;
#1 $display("%b", po);
# 1  pi=13'b0100001101010;
#1 $display("%b", po);
# 1  pi=13'b0100001101011;
#1 $display("%b", po);
# 1  pi=13'b0100001101100;
#1 $display("%b", po);
# 1  pi=13'b0100001101101;
#1 $display("%b", po);
# 1  pi=13'b0100001101110;
#1 $display("%b", po);
# 1  pi=13'b0100001101111;
#1 $display("%b", po);
# 1  pi=13'b0100001110000;
#1 $display("%b", po);
# 1  pi=13'b0100001110001;
#1 $display("%b", po);
# 1  pi=13'b0100001110010;
#1 $display("%b", po);
# 1  pi=13'b0100001110011;
#1 $display("%b", po);
# 1  pi=13'b0100001110100;
#1 $display("%b", po);
# 1  pi=13'b0100001110101;
#1 $display("%b", po);
# 1  pi=13'b0100001110110;
#1 $display("%b", po);
# 1  pi=13'b0100001110111;
#1 $display("%b", po);
# 1  pi=13'b0100001111000;
#1 $display("%b", po);
# 1  pi=13'b0100001111001;
#1 $display("%b", po);
# 1  pi=13'b0100001111010;
#1 $display("%b", po);
# 1  pi=13'b0100001111011;
#1 $display("%b", po);
# 1  pi=13'b0100001111100;
#1 $display("%b", po);
# 1  pi=13'b0100001111101;
#1 $display("%b", po);
# 1  pi=13'b0100001111110;
#1 $display("%b", po);
# 1  pi=13'b0100001111111;
#1 $display("%b", po);
# 1  pi=13'b0100010000000;
#1 $display("%b", po);
# 1  pi=13'b0100010000001;
#1 $display("%b", po);
# 1  pi=13'b0100010000010;
#1 $display("%b", po);
# 1  pi=13'b0100010000011;
#1 $display("%b", po);
# 1  pi=13'b0100010000100;
#1 $display("%b", po);
# 1  pi=13'b0100010000101;
#1 $display("%b", po);
# 1  pi=13'b0100010000110;
#1 $display("%b", po);
# 1  pi=13'b0100010000111;
#1 $display("%b", po);
# 1  pi=13'b0100010001000;
#1 $display("%b", po);
# 1  pi=13'b0100010001001;
#1 $display("%b", po);
# 1  pi=13'b0100010001010;
#1 $display("%b", po);
# 1  pi=13'b0100010001011;
#1 $display("%b", po);
# 1  pi=13'b0100010001100;
#1 $display("%b", po);
# 1  pi=13'b0100010001101;
#1 $display("%b", po);
# 1  pi=13'b0100010001110;
#1 $display("%b", po);
# 1  pi=13'b0100010001111;
#1 $display("%b", po);
# 1  pi=13'b0100010010000;
#1 $display("%b", po);
# 1  pi=13'b0100010010001;
#1 $display("%b", po);
# 1  pi=13'b0100010010010;
#1 $display("%b", po);
# 1  pi=13'b0100010010011;
#1 $display("%b", po);
# 1  pi=13'b0100010010100;
#1 $display("%b", po);
# 1  pi=13'b0100010010101;
#1 $display("%b", po);
# 1  pi=13'b0100010010110;
#1 $display("%b", po);
# 1  pi=13'b0100010010111;
#1 $display("%b", po);
# 1  pi=13'b0100010011000;
#1 $display("%b", po);
# 1  pi=13'b0100010011001;
#1 $display("%b", po);
# 1  pi=13'b0100010011010;
#1 $display("%b", po);
# 1  pi=13'b0100010011011;
#1 $display("%b", po);
# 1  pi=13'b0100010011100;
#1 $display("%b", po);
# 1  pi=13'b0100010011101;
#1 $display("%b", po);
# 1  pi=13'b0100010011110;
#1 $display("%b", po);
# 1  pi=13'b0100010011111;
#1 $display("%b", po);
# 1  pi=13'b0100010100000;
#1 $display("%b", po);
# 1  pi=13'b0100010100001;
#1 $display("%b", po);
# 1  pi=13'b0100010100010;
#1 $display("%b", po);
# 1  pi=13'b0100010100011;
#1 $display("%b", po);
# 1  pi=13'b0100010100100;
#1 $display("%b", po);
# 1  pi=13'b0100010100101;
#1 $display("%b", po);
# 1  pi=13'b0100010100110;
#1 $display("%b", po);
# 1  pi=13'b0100010100111;
#1 $display("%b", po);
# 1  pi=13'b0100010101000;
#1 $display("%b", po);
# 1  pi=13'b0100010101001;
#1 $display("%b", po);
# 1  pi=13'b0100010101010;
#1 $display("%b", po);
# 1  pi=13'b0100010101011;
#1 $display("%b", po);
# 1  pi=13'b0100010101100;
#1 $display("%b", po);
# 1  pi=13'b0100010101101;
#1 $display("%b", po);
# 1  pi=13'b0100010101110;
#1 $display("%b", po);
# 1  pi=13'b0100010101111;
#1 $display("%b", po);
# 1  pi=13'b0100010110000;
#1 $display("%b", po);
# 1  pi=13'b0100010110001;
#1 $display("%b", po);
# 1  pi=13'b0100010110010;
#1 $display("%b", po);
# 1  pi=13'b0100010110011;
#1 $display("%b", po);
# 1  pi=13'b0100010110100;
#1 $display("%b", po);
# 1  pi=13'b0100010110101;
#1 $display("%b", po);
# 1  pi=13'b0100010110110;
#1 $display("%b", po);
# 1  pi=13'b0100010110111;
#1 $display("%b", po);
# 1  pi=13'b0100010111000;
#1 $display("%b", po);
# 1  pi=13'b0100010111001;
#1 $display("%b", po);
# 1  pi=13'b0100010111010;
#1 $display("%b", po);
# 1  pi=13'b0100010111011;
#1 $display("%b", po);
# 1  pi=13'b0100010111100;
#1 $display("%b", po);
# 1  pi=13'b0100010111101;
#1 $display("%b", po);
# 1  pi=13'b0100010111110;
#1 $display("%b", po);
# 1  pi=13'b0100010111111;
#1 $display("%b", po);
# 1  pi=13'b0100011000000;
#1 $display("%b", po);
# 1  pi=13'b0100011000001;
#1 $display("%b", po);
# 1  pi=13'b0100011000010;
#1 $display("%b", po);
# 1  pi=13'b0100011000011;
#1 $display("%b", po);
# 1  pi=13'b0100011000100;
#1 $display("%b", po);
# 1  pi=13'b0100011000101;
#1 $display("%b", po);
# 1  pi=13'b0100011000110;
#1 $display("%b", po);
# 1  pi=13'b0100011000111;
#1 $display("%b", po);
# 1  pi=13'b0100011001000;
#1 $display("%b", po);
# 1  pi=13'b0100011001001;
#1 $display("%b", po);
# 1  pi=13'b0100011001010;
#1 $display("%b", po);
# 1  pi=13'b0100011001011;
#1 $display("%b", po);
# 1  pi=13'b0100011001100;
#1 $display("%b", po);
# 1  pi=13'b0100011001101;
#1 $display("%b", po);
# 1  pi=13'b0100011001110;
#1 $display("%b", po);
# 1  pi=13'b0100011001111;
#1 $display("%b", po);
# 1  pi=13'b0100011010000;
#1 $display("%b", po);
# 1  pi=13'b0100011010001;
#1 $display("%b", po);
# 1  pi=13'b0100011010010;
#1 $display("%b", po);
# 1  pi=13'b0100011010011;
#1 $display("%b", po);
# 1  pi=13'b0100011010100;
#1 $display("%b", po);
# 1  pi=13'b0100011010101;
#1 $display("%b", po);
# 1  pi=13'b0100011010110;
#1 $display("%b", po);
# 1  pi=13'b0100011010111;
#1 $display("%b", po);
# 1  pi=13'b0100011011000;
#1 $display("%b", po);
# 1  pi=13'b0100011011001;
#1 $display("%b", po);
# 1  pi=13'b0100011011010;
#1 $display("%b", po);
# 1  pi=13'b0100011011011;
#1 $display("%b", po);
# 1  pi=13'b0100011011100;
#1 $display("%b", po);
# 1  pi=13'b0100011011101;
#1 $display("%b", po);
# 1  pi=13'b0100011011110;
#1 $display("%b", po);
# 1  pi=13'b0100011011111;
#1 $display("%b", po);
# 1  pi=13'b0100011100000;
#1 $display("%b", po);
# 1  pi=13'b0100011100001;
#1 $display("%b", po);
# 1  pi=13'b0100011100010;
#1 $display("%b", po);
# 1  pi=13'b0100011100011;
#1 $display("%b", po);
# 1  pi=13'b0100011100100;
#1 $display("%b", po);
# 1  pi=13'b0100011100101;
#1 $display("%b", po);
# 1  pi=13'b0100011100110;
#1 $display("%b", po);
# 1  pi=13'b0100011100111;
#1 $display("%b", po);
# 1  pi=13'b0100011101000;
#1 $display("%b", po);
# 1  pi=13'b0100011101001;
#1 $display("%b", po);
# 1  pi=13'b0100011101010;
#1 $display("%b", po);
# 1  pi=13'b0100011101011;
#1 $display("%b", po);
# 1  pi=13'b0100011101100;
#1 $display("%b", po);
# 1  pi=13'b0100011101101;
#1 $display("%b", po);
# 1  pi=13'b0100011101110;
#1 $display("%b", po);
# 1  pi=13'b0100011101111;
#1 $display("%b", po);
# 1  pi=13'b0100011110000;
#1 $display("%b", po);
# 1  pi=13'b0100011110001;
#1 $display("%b", po);
# 1  pi=13'b0100011110010;
#1 $display("%b", po);
# 1  pi=13'b0100011110011;
#1 $display("%b", po);
# 1  pi=13'b0100011110100;
#1 $display("%b", po);
# 1  pi=13'b0100011110101;
#1 $display("%b", po);
# 1  pi=13'b0100011110110;
#1 $display("%b", po);
# 1  pi=13'b0100011110111;
#1 $display("%b", po);
# 1  pi=13'b0100011111000;
#1 $display("%b", po);
# 1  pi=13'b0100011111001;
#1 $display("%b", po);
# 1  pi=13'b0100011111010;
#1 $display("%b", po);
# 1  pi=13'b0100011111011;
#1 $display("%b", po);
# 1  pi=13'b0100011111100;
#1 $display("%b", po);
# 1  pi=13'b0100011111101;
#1 $display("%b", po);
# 1  pi=13'b0100011111110;
#1 $display("%b", po);
# 1  pi=13'b0100011111111;
#1 $display("%b", po);
# 1  pi=13'b0100100000000;
#1 $display("%b", po);
# 1  pi=13'b0100100000001;
#1 $display("%b", po);
# 1  pi=13'b0100100000010;
#1 $display("%b", po);
# 1  pi=13'b0100100000011;
#1 $display("%b", po);
# 1  pi=13'b0100100000100;
#1 $display("%b", po);
# 1  pi=13'b0100100000101;
#1 $display("%b", po);
# 1  pi=13'b0100100000110;
#1 $display("%b", po);
# 1  pi=13'b0100100000111;
#1 $display("%b", po);
# 1  pi=13'b0100100001000;
#1 $display("%b", po);
# 1  pi=13'b0100100001001;
#1 $display("%b", po);
# 1  pi=13'b0100100001010;
#1 $display("%b", po);
# 1  pi=13'b0100100001011;
#1 $display("%b", po);
# 1  pi=13'b0100100001100;
#1 $display("%b", po);
# 1  pi=13'b0100100001101;
#1 $display("%b", po);
# 1  pi=13'b0100100001110;
#1 $display("%b", po);
# 1  pi=13'b0100100001111;
#1 $display("%b", po);
# 1  pi=13'b0100100010000;
#1 $display("%b", po);
# 1  pi=13'b0100100010001;
#1 $display("%b", po);
# 1  pi=13'b0100100010010;
#1 $display("%b", po);
# 1  pi=13'b0100100010011;
#1 $display("%b", po);
# 1  pi=13'b0100100010100;
#1 $display("%b", po);
# 1  pi=13'b0100100010101;
#1 $display("%b", po);
# 1  pi=13'b0100100010110;
#1 $display("%b", po);
# 1  pi=13'b0100100010111;
#1 $display("%b", po);
# 1  pi=13'b0100100011000;
#1 $display("%b", po);
# 1  pi=13'b0100100011001;
#1 $display("%b", po);
# 1  pi=13'b0100100011010;
#1 $display("%b", po);
# 1  pi=13'b0100100011011;
#1 $display("%b", po);
# 1  pi=13'b0100100011100;
#1 $display("%b", po);
# 1  pi=13'b0100100011101;
#1 $display("%b", po);
# 1  pi=13'b0100100011110;
#1 $display("%b", po);
# 1  pi=13'b0100100011111;
#1 $display("%b", po);
# 1  pi=13'b0100100100000;
#1 $display("%b", po);
# 1  pi=13'b0100100100001;
#1 $display("%b", po);
# 1  pi=13'b0100100100010;
#1 $display("%b", po);
# 1  pi=13'b0100100100011;
#1 $display("%b", po);
# 1  pi=13'b0100100100100;
#1 $display("%b", po);
# 1  pi=13'b0100100100101;
#1 $display("%b", po);
# 1  pi=13'b0100100100110;
#1 $display("%b", po);
# 1  pi=13'b0100100100111;
#1 $display("%b", po);
# 1  pi=13'b0100100101000;
#1 $display("%b", po);
# 1  pi=13'b0100100101001;
#1 $display("%b", po);
# 1  pi=13'b0100100101010;
#1 $display("%b", po);
# 1  pi=13'b0100100101011;
#1 $display("%b", po);
# 1  pi=13'b0100100101100;
#1 $display("%b", po);
# 1  pi=13'b0100100101101;
#1 $display("%b", po);
# 1  pi=13'b0100100101110;
#1 $display("%b", po);
# 1  pi=13'b0100100101111;
#1 $display("%b", po);
# 1  pi=13'b0100100110000;
#1 $display("%b", po);
# 1  pi=13'b0100100110001;
#1 $display("%b", po);
# 1  pi=13'b0100100110010;
#1 $display("%b", po);
# 1  pi=13'b0100100110011;
#1 $display("%b", po);
# 1  pi=13'b0100100110100;
#1 $display("%b", po);
# 1  pi=13'b0100100110101;
#1 $display("%b", po);
# 1  pi=13'b0100100110110;
#1 $display("%b", po);
# 1  pi=13'b0100100110111;
#1 $display("%b", po);
# 1  pi=13'b0100100111000;
#1 $display("%b", po);
# 1  pi=13'b0100100111001;
#1 $display("%b", po);
# 1  pi=13'b0100100111010;
#1 $display("%b", po);
# 1  pi=13'b0100100111011;
#1 $display("%b", po);
# 1  pi=13'b0100100111100;
#1 $display("%b", po);
# 1  pi=13'b0100100111101;
#1 $display("%b", po);
# 1  pi=13'b0100100111110;
#1 $display("%b", po);
# 1  pi=13'b0100100111111;
#1 $display("%b", po);
# 1  pi=13'b0100101000000;
#1 $display("%b", po);
# 1  pi=13'b0100101000001;
#1 $display("%b", po);
# 1  pi=13'b0100101000010;
#1 $display("%b", po);
# 1  pi=13'b0100101000011;
#1 $display("%b", po);
# 1  pi=13'b0100101000100;
#1 $display("%b", po);
# 1  pi=13'b0100101000101;
#1 $display("%b", po);
# 1  pi=13'b0100101000110;
#1 $display("%b", po);
# 1  pi=13'b0100101000111;
#1 $display("%b", po);
# 1  pi=13'b0100101001000;
#1 $display("%b", po);
# 1  pi=13'b0100101001001;
#1 $display("%b", po);
# 1  pi=13'b0100101001010;
#1 $display("%b", po);
# 1  pi=13'b0100101001011;
#1 $display("%b", po);
# 1  pi=13'b0100101001100;
#1 $display("%b", po);
# 1  pi=13'b0100101001101;
#1 $display("%b", po);
# 1  pi=13'b0100101001110;
#1 $display("%b", po);
# 1  pi=13'b0100101001111;
#1 $display("%b", po);
# 1  pi=13'b0100101010000;
#1 $display("%b", po);
# 1  pi=13'b0100101010001;
#1 $display("%b", po);
# 1  pi=13'b0100101010010;
#1 $display("%b", po);
# 1  pi=13'b0100101010011;
#1 $display("%b", po);
# 1  pi=13'b0100101010100;
#1 $display("%b", po);
# 1  pi=13'b0100101010101;
#1 $display("%b", po);
# 1  pi=13'b0100101010110;
#1 $display("%b", po);
# 1  pi=13'b0100101010111;
#1 $display("%b", po);
# 1  pi=13'b0100101011000;
#1 $display("%b", po);
# 1  pi=13'b0100101011001;
#1 $display("%b", po);
# 1  pi=13'b0100101011010;
#1 $display("%b", po);
# 1  pi=13'b0100101011011;
#1 $display("%b", po);
# 1  pi=13'b0100101011100;
#1 $display("%b", po);
# 1  pi=13'b0100101011101;
#1 $display("%b", po);
# 1  pi=13'b0100101011110;
#1 $display("%b", po);
# 1  pi=13'b0100101011111;
#1 $display("%b", po);
# 1  pi=13'b0100101100000;
#1 $display("%b", po);
# 1  pi=13'b0100101100001;
#1 $display("%b", po);
# 1  pi=13'b0100101100010;
#1 $display("%b", po);
# 1  pi=13'b0100101100011;
#1 $display("%b", po);
# 1  pi=13'b0100101100100;
#1 $display("%b", po);
# 1  pi=13'b0100101100101;
#1 $display("%b", po);
# 1  pi=13'b0100101100110;
#1 $display("%b", po);
# 1  pi=13'b0100101100111;
#1 $display("%b", po);
# 1  pi=13'b0100101101000;
#1 $display("%b", po);
# 1  pi=13'b0100101101001;
#1 $display("%b", po);
# 1  pi=13'b0100101101010;
#1 $display("%b", po);
# 1  pi=13'b0100101101011;
#1 $display("%b", po);
# 1  pi=13'b0100101101100;
#1 $display("%b", po);
# 1  pi=13'b0100101101101;
#1 $display("%b", po);
# 1  pi=13'b0100101101110;
#1 $display("%b", po);
# 1  pi=13'b0100101101111;
#1 $display("%b", po);
# 1  pi=13'b0100101110000;
#1 $display("%b", po);
# 1  pi=13'b0100101110001;
#1 $display("%b", po);
# 1  pi=13'b0100101110010;
#1 $display("%b", po);
# 1  pi=13'b0100101110011;
#1 $display("%b", po);
# 1  pi=13'b0100101110100;
#1 $display("%b", po);
# 1  pi=13'b0100101110101;
#1 $display("%b", po);
# 1  pi=13'b0100101110110;
#1 $display("%b", po);
# 1  pi=13'b0100101110111;
#1 $display("%b", po);
# 1  pi=13'b0100101111000;
#1 $display("%b", po);
# 1  pi=13'b0100101111001;
#1 $display("%b", po);
# 1  pi=13'b0100101111010;
#1 $display("%b", po);
# 1  pi=13'b0100101111011;
#1 $display("%b", po);
# 1  pi=13'b0100101111100;
#1 $display("%b", po);
# 1  pi=13'b0100101111101;
#1 $display("%b", po);
# 1  pi=13'b0100101111110;
#1 $display("%b", po);
# 1  pi=13'b0100101111111;
#1 $display("%b", po);
# 1  pi=13'b0100110000000;
#1 $display("%b", po);
# 1  pi=13'b0100110000001;
#1 $display("%b", po);
# 1  pi=13'b0100110000010;
#1 $display("%b", po);
# 1  pi=13'b0100110000011;
#1 $display("%b", po);
# 1  pi=13'b0100110000100;
#1 $display("%b", po);
# 1  pi=13'b0100110000101;
#1 $display("%b", po);
# 1  pi=13'b0100110000110;
#1 $display("%b", po);
# 1  pi=13'b0100110000111;
#1 $display("%b", po);
# 1  pi=13'b0100110001000;
#1 $display("%b", po);
# 1  pi=13'b0100110001001;
#1 $display("%b", po);
# 1  pi=13'b0100110001010;
#1 $display("%b", po);
# 1  pi=13'b0100110001011;
#1 $display("%b", po);
# 1  pi=13'b0100110001100;
#1 $display("%b", po);
# 1  pi=13'b0100110001101;
#1 $display("%b", po);
# 1  pi=13'b0100110001110;
#1 $display("%b", po);
# 1  pi=13'b0100110001111;
#1 $display("%b", po);
# 1  pi=13'b0100110010000;
#1 $display("%b", po);
# 1  pi=13'b0100110010001;
#1 $display("%b", po);
# 1  pi=13'b0100110010010;
#1 $display("%b", po);
# 1  pi=13'b0100110010011;
#1 $display("%b", po);
# 1  pi=13'b0100110010100;
#1 $display("%b", po);
# 1  pi=13'b0100110010101;
#1 $display("%b", po);
# 1  pi=13'b0100110010110;
#1 $display("%b", po);
# 1  pi=13'b0100110010111;
#1 $display("%b", po);
# 1  pi=13'b0100110011000;
#1 $display("%b", po);
# 1  pi=13'b0100110011001;
#1 $display("%b", po);
# 1  pi=13'b0100110011010;
#1 $display("%b", po);
# 1  pi=13'b0100110011011;
#1 $display("%b", po);
# 1  pi=13'b0100110011100;
#1 $display("%b", po);
# 1  pi=13'b0100110011101;
#1 $display("%b", po);
# 1  pi=13'b0100110011110;
#1 $display("%b", po);
# 1  pi=13'b0100110011111;
#1 $display("%b", po);
# 1  pi=13'b0100110100000;
#1 $display("%b", po);
# 1  pi=13'b0100110100001;
#1 $display("%b", po);
# 1  pi=13'b0100110100010;
#1 $display("%b", po);
# 1  pi=13'b0100110100011;
#1 $display("%b", po);
# 1  pi=13'b0100110100100;
#1 $display("%b", po);
# 1  pi=13'b0100110100101;
#1 $display("%b", po);
# 1  pi=13'b0100110100110;
#1 $display("%b", po);
# 1  pi=13'b0100110100111;
#1 $display("%b", po);
# 1  pi=13'b0100110101000;
#1 $display("%b", po);
# 1  pi=13'b0100110101001;
#1 $display("%b", po);
# 1  pi=13'b0100110101010;
#1 $display("%b", po);
# 1  pi=13'b0100110101011;
#1 $display("%b", po);
# 1  pi=13'b0100110101100;
#1 $display("%b", po);
# 1  pi=13'b0100110101101;
#1 $display("%b", po);
# 1  pi=13'b0100110101110;
#1 $display("%b", po);
# 1  pi=13'b0100110101111;
#1 $display("%b", po);
# 1  pi=13'b0100110110000;
#1 $display("%b", po);
# 1  pi=13'b0100110110001;
#1 $display("%b", po);
# 1  pi=13'b0100110110010;
#1 $display("%b", po);
# 1  pi=13'b0100110110011;
#1 $display("%b", po);
# 1  pi=13'b0100110110100;
#1 $display("%b", po);
# 1  pi=13'b0100110110101;
#1 $display("%b", po);
# 1  pi=13'b0100110110110;
#1 $display("%b", po);
# 1  pi=13'b0100110110111;
#1 $display("%b", po);
# 1  pi=13'b0100110111000;
#1 $display("%b", po);
# 1  pi=13'b0100110111001;
#1 $display("%b", po);
# 1  pi=13'b0100110111010;
#1 $display("%b", po);
# 1  pi=13'b0100110111011;
#1 $display("%b", po);
# 1  pi=13'b0100110111100;
#1 $display("%b", po);
# 1  pi=13'b0100110111101;
#1 $display("%b", po);
# 1  pi=13'b0100110111110;
#1 $display("%b", po);
# 1  pi=13'b0100110111111;
#1 $display("%b", po);
# 1  pi=13'b0100111000000;
#1 $display("%b", po);
# 1  pi=13'b0100111000001;
#1 $display("%b", po);
# 1  pi=13'b0100111000010;
#1 $display("%b", po);
# 1  pi=13'b0100111000011;
#1 $display("%b", po);
# 1  pi=13'b0100111000100;
#1 $display("%b", po);
# 1  pi=13'b0100111000101;
#1 $display("%b", po);
# 1  pi=13'b0100111000110;
#1 $display("%b", po);
# 1  pi=13'b0100111000111;
#1 $display("%b", po);
# 1  pi=13'b0100111001000;
#1 $display("%b", po);
# 1  pi=13'b0100111001001;
#1 $display("%b", po);
# 1  pi=13'b0100111001010;
#1 $display("%b", po);
# 1  pi=13'b0100111001011;
#1 $display("%b", po);
# 1  pi=13'b0100111001100;
#1 $display("%b", po);
# 1  pi=13'b0100111001101;
#1 $display("%b", po);
# 1  pi=13'b0100111001110;
#1 $display("%b", po);
# 1  pi=13'b0100111001111;
#1 $display("%b", po);
# 1  pi=13'b0100111010000;
#1 $display("%b", po);
# 1  pi=13'b0100111010001;
#1 $display("%b", po);
# 1  pi=13'b0100111010010;
#1 $display("%b", po);
# 1  pi=13'b0100111010011;
#1 $display("%b", po);
# 1  pi=13'b0100111010100;
#1 $display("%b", po);
# 1  pi=13'b0100111010101;
#1 $display("%b", po);
# 1  pi=13'b0100111010110;
#1 $display("%b", po);
# 1  pi=13'b0100111010111;
#1 $display("%b", po);
# 1  pi=13'b0100111011000;
#1 $display("%b", po);
# 1  pi=13'b0100111011001;
#1 $display("%b", po);
# 1  pi=13'b0100111011010;
#1 $display("%b", po);
# 1  pi=13'b0100111011011;
#1 $display("%b", po);
# 1  pi=13'b0100111011100;
#1 $display("%b", po);
# 1  pi=13'b0100111011101;
#1 $display("%b", po);
# 1  pi=13'b0100111011110;
#1 $display("%b", po);
# 1  pi=13'b0100111011111;
#1 $display("%b", po);
# 1  pi=13'b0100111100000;
#1 $display("%b", po);
# 1  pi=13'b0100111100001;
#1 $display("%b", po);
# 1  pi=13'b0100111100010;
#1 $display("%b", po);
# 1  pi=13'b0100111100011;
#1 $display("%b", po);
# 1  pi=13'b0100111100100;
#1 $display("%b", po);
# 1  pi=13'b0100111100101;
#1 $display("%b", po);
# 1  pi=13'b0100111100110;
#1 $display("%b", po);
# 1  pi=13'b0100111100111;
#1 $display("%b", po);
# 1  pi=13'b0100111101000;
#1 $display("%b", po);
# 1  pi=13'b0100111101001;
#1 $display("%b", po);
# 1  pi=13'b0100111101010;
#1 $display("%b", po);
# 1  pi=13'b0100111101011;
#1 $display("%b", po);
# 1  pi=13'b0100111101100;
#1 $display("%b", po);
# 1  pi=13'b0100111101101;
#1 $display("%b", po);
# 1  pi=13'b0100111101110;
#1 $display("%b", po);
# 1  pi=13'b0100111101111;
#1 $display("%b", po);
# 1  pi=13'b0100111110000;
#1 $display("%b", po);
# 1  pi=13'b0100111110001;
#1 $display("%b", po);
# 1  pi=13'b0100111110010;
#1 $display("%b", po);
# 1  pi=13'b0100111110011;
#1 $display("%b", po);
# 1  pi=13'b0100111110100;
#1 $display("%b", po);
# 1  pi=13'b0100111110101;
#1 $display("%b", po);
# 1  pi=13'b0100111110110;
#1 $display("%b", po);
# 1  pi=13'b0100111110111;
#1 $display("%b", po);
# 1  pi=13'b0100111111000;
#1 $display("%b", po);
# 1  pi=13'b0100111111001;
#1 $display("%b", po);
# 1  pi=13'b0100111111010;
#1 $display("%b", po);
# 1  pi=13'b0100111111011;
#1 $display("%b", po);
# 1  pi=13'b0100111111100;
#1 $display("%b", po);
# 1  pi=13'b0100111111101;
#1 $display("%b", po);
# 1  pi=13'b0100111111110;
#1 $display("%b", po);
# 1  pi=13'b0100111111111;
#1 $display("%b", po);
# 1  pi=13'b0101000000000;
#1 $display("%b", po);
# 1  pi=13'b0101000000001;
#1 $display("%b", po);
# 1  pi=13'b0101000000010;
#1 $display("%b", po);
# 1  pi=13'b0101000000011;
#1 $display("%b", po);
# 1  pi=13'b0101000000100;
#1 $display("%b", po);
# 1  pi=13'b0101000000101;
#1 $display("%b", po);
# 1  pi=13'b0101000000110;
#1 $display("%b", po);
# 1  pi=13'b0101000000111;
#1 $display("%b", po);
# 1  pi=13'b0101000001000;
#1 $display("%b", po);
# 1  pi=13'b0101000001001;
#1 $display("%b", po);
# 1  pi=13'b0101000001010;
#1 $display("%b", po);
# 1  pi=13'b0101000001011;
#1 $display("%b", po);
# 1  pi=13'b0101000001100;
#1 $display("%b", po);
# 1  pi=13'b0101000001101;
#1 $display("%b", po);
# 1  pi=13'b0101000001110;
#1 $display("%b", po);
# 1  pi=13'b0101000001111;
#1 $display("%b", po);
# 1  pi=13'b0101000010000;
#1 $display("%b", po);
# 1  pi=13'b0101000010001;
#1 $display("%b", po);
# 1  pi=13'b0101000010010;
#1 $display("%b", po);
# 1  pi=13'b0101000010011;
#1 $display("%b", po);
# 1  pi=13'b0101000010100;
#1 $display("%b", po);
# 1  pi=13'b0101000010101;
#1 $display("%b", po);
# 1  pi=13'b0101000010110;
#1 $display("%b", po);
# 1  pi=13'b0101000010111;
#1 $display("%b", po);
# 1  pi=13'b0101000011000;
#1 $display("%b", po);
# 1  pi=13'b0101000011001;
#1 $display("%b", po);
# 1  pi=13'b0101000011010;
#1 $display("%b", po);
# 1  pi=13'b0101000011011;
#1 $display("%b", po);
# 1  pi=13'b0101000011100;
#1 $display("%b", po);
# 1  pi=13'b0101000011101;
#1 $display("%b", po);
# 1  pi=13'b0101000011110;
#1 $display("%b", po);
# 1  pi=13'b0101000011111;
#1 $display("%b", po);
# 1  pi=13'b0101000100000;
#1 $display("%b", po);
# 1  pi=13'b0101000100001;
#1 $display("%b", po);
# 1  pi=13'b0101000100010;
#1 $display("%b", po);
# 1  pi=13'b0101000100011;
#1 $display("%b", po);
# 1  pi=13'b0101000100100;
#1 $display("%b", po);
# 1  pi=13'b0101000100101;
#1 $display("%b", po);
# 1  pi=13'b0101000100110;
#1 $display("%b", po);
# 1  pi=13'b0101000100111;
#1 $display("%b", po);
# 1  pi=13'b0101000101000;
#1 $display("%b", po);
# 1  pi=13'b0101000101001;
#1 $display("%b", po);
# 1  pi=13'b0101000101010;
#1 $display("%b", po);
# 1  pi=13'b0101000101011;
#1 $display("%b", po);
# 1  pi=13'b0101000101100;
#1 $display("%b", po);
# 1  pi=13'b0101000101101;
#1 $display("%b", po);
# 1  pi=13'b0101000101110;
#1 $display("%b", po);
# 1  pi=13'b0101000101111;
#1 $display("%b", po);
# 1  pi=13'b0101000110000;
#1 $display("%b", po);
# 1  pi=13'b0101000110001;
#1 $display("%b", po);
# 1  pi=13'b0101000110010;
#1 $display("%b", po);
# 1  pi=13'b0101000110011;
#1 $display("%b", po);
# 1  pi=13'b0101000110100;
#1 $display("%b", po);
# 1  pi=13'b0101000110101;
#1 $display("%b", po);
# 1  pi=13'b0101000110110;
#1 $display("%b", po);
# 1  pi=13'b0101000110111;
#1 $display("%b", po);
# 1  pi=13'b0101000111000;
#1 $display("%b", po);
# 1  pi=13'b0101000111001;
#1 $display("%b", po);
# 1  pi=13'b0101000111010;
#1 $display("%b", po);
# 1  pi=13'b0101000111011;
#1 $display("%b", po);
# 1  pi=13'b0101000111100;
#1 $display("%b", po);
# 1  pi=13'b0101000111101;
#1 $display("%b", po);
# 1  pi=13'b0101000111110;
#1 $display("%b", po);
# 1  pi=13'b0101000111111;
#1 $display("%b", po);
# 1  pi=13'b0101001000000;
#1 $display("%b", po);
# 1  pi=13'b0101001000001;
#1 $display("%b", po);
# 1  pi=13'b0101001000010;
#1 $display("%b", po);
# 1  pi=13'b0101001000011;
#1 $display("%b", po);
# 1  pi=13'b0101001000100;
#1 $display("%b", po);
# 1  pi=13'b0101001000101;
#1 $display("%b", po);
# 1  pi=13'b0101001000110;
#1 $display("%b", po);
# 1  pi=13'b0101001000111;
#1 $display("%b", po);
# 1  pi=13'b0101001001000;
#1 $display("%b", po);
# 1  pi=13'b0101001001001;
#1 $display("%b", po);
# 1  pi=13'b0101001001010;
#1 $display("%b", po);
# 1  pi=13'b0101001001011;
#1 $display("%b", po);
# 1  pi=13'b0101001001100;
#1 $display("%b", po);
# 1  pi=13'b0101001001101;
#1 $display("%b", po);
# 1  pi=13'b0101001001110;
#1 $display("%b", po);
# 1  pi=13'b0101001001111;
#1 $display("%b", po);
# 1  pi=13'b0101001010000;
#1 $display("%b", po);
# 1  pi=13'b0101001010001;
#1 $display("%b", po);
# 1  pi=13'b0101001010010;
#1 $display("%b", po);
# 1  pi=13'b0101001010011;
#1 $display("%b", po);
# 1  pi=13'b0101001010100;
#1 $display("%b", po);
# 1  pi=13'b0101001010101;
#1 $display("%b", po);
# 1  pi=13'b0101001010110;
#1 $display("%b", po);
# 1  pi=13'b0101001010111;
#1 $display("%b", po);
# 1  pi=13'b0101001011000;
#1 $display("%b", po);
# 1  pi=13'b0101001011001;
#1 $display("%b", po);
# 1  pi=13'b0101001011010;
#1 $display("%b", po);
# 1  pi=13'b0101001011011;
#1 $display("%b", po);
# 1  pi=13'b0101001011100;
#1 $display("%b", po);
# 1  pi=13'b0101001011101;
#1 $display("%b", po);
# 1  pi=13'b0101001011110;
#1 $display("%b", po);
# 1  pi=13'b0101001011111;
#1 $display("%b", po);
# 1  pi=13'b0101001100000;
#1 $display("%b", po);
# 1  pi=13'b0101001100001;
#1 $display("%b", po);
# 1  pi=13'b0101001100010;
#1 $display("%b", po);
# 1  pi=13'b0101001100011;
#1 $display("%b", po);
# 1  pi=13'b0101001100100;
#1 $display("%b", po);
# 1  pi=13'b0101001100101;
#1 $display("%b", po);
# 1  pi=13'b0101001100110;
#1 $display("%b", po);
# 1  pi=13'b0101001100111;
#1 $display("%b", po);
# 1  pi=13'b0101001101000;
#1 $display("%b", po);
# 1  pi=13'b0101001101001;
#1 $display("%b", po);
# 1  pi=13'b0101001101010;
#1 $display("%b", po);
# 1  pi=13'b0101001101011;
#1 $display("%b", po);
# 1  pi=13'b0101001101100;
#1 $display("%b", po);
# 1  pi=13'b0101001101101;
#1 $display("%b", po);
# 1  pi=13'b0101001101110;
#1 $display("%b", po);
# 1  pi=13'b0101001101111;
#1 $display("%b", po);
# 1  pi=13'b0101001110000;
#1 $display("%b", po);
# 1  pi=13'b0101001110001;
#1 $display("%b", po);
# 1  pi=13'b0101001110010;
#1 $display("%b", po);
# 1  pi=13'b0101001110011;
#1 $display("%b", po);
# 1  pi=13'b0101001110100;
#1 $display("%b", po);
# 1  pi=13'b0101001110101;
#1 $display("%b", po);
# 1  pi=13'b0101001110110;
#1 $display("%b", po);
# 1  pi=13'b0101001110111;
#1 $display("%b", po);
# 1  pi=13'b0101001111000;
#1 $display("%b", po);
# 1  pi=13'b0101001111001;
#1 $display("%b", po);
# 1  pi=13'b0101001111010;
#1 $display("%b", po);
# 1  pi=13'b0101001111011;
#1 $display("%b", po);
# 1  pi=13'b0101001111100;
#1 $display("%b", po);
# 1  pi=13'b0101001111101;
#1 $display("%b", po);
# 1  pi=13'b0101001111110;
#1 $display("%b", po);
# 1  pi=13'b0101001111111;
#1 $display("%b", po);
# 1  pi=13'b0101010000000;
#1 $display("%b", po);
# 1  pi=13'b0101010000001;
#1 $display("%b", po);
# 1  pi=13'b0101010000010;
#1 $display("%b", po);
# 1  pi=13'b0101010000011;
#1 $display("%b", po);
# 1  pi=13'b0101010000100;
#1 $display("%b", po);
# 1  pi=13'b0101010000101;
#1 $display("%b", po);
# 1  pi=13'b0101010000110;
#1 $display("%b", po);
# 1  pi=13'b0101010000111;
#1 $display("%b", po);
# 1  pi=13'b0101010001000;
#1 $display("%b", po);
# 1  pi=13'b0101010001001;
#1 $display("%b", po);
# 1  pi=13'b0101010001010;
#1 $display("%b", po);
# 1  pi=13'b0101010001011;
#1 $display("%b", po);
# 1  pi=13'b0101010001100;
#1 $display("%b", po);
# 1  pi=13'b0101010001101;
#1 $display("%b", po);
# 1  pi=13'b0101010001110;
#1 $display("%b", po);
# 1  pi=13'b0101010001111;
#1 $display("%b", po);
# 1  pi=13'b0101010010000;
#1 $display("%b", po);
# 1  pi=13'b0101010010001;
#1 $display("%b", po);
# 1  pi=13'b0101010010010;
#1 $display("%b", po);
# 1  pi=13'b0101010010011;
#1 $display("%b", po);
# 1  pi=13'b0101010010100;
#1 $display("%b", po);
# 1  pi=13'b0101010010101;
#1 $display("%b", po);
# 1  pi=13'b0101010010110;
#1 $display("%b", po);
# 1  pi=13'b0101010010111;
#1 $display("%b", po);
# 1  pi=13'b0101010011000;
#1 $display("%b", po);
# 1  pi=13'b0101010011001;
#1 $display("%b", po);
# 1  pi=13'b0101010011010;
#1 $display("%b", po);
# 1  pi=13'b0101010011011;
#1 $display("%b", po);
# 1  pi=13'b0101010011100;
#1 $display("%b", po);
# 1  pi=13'b0101010011101;
#1 $display("%b", po);
# 1  pi=13'b0101010011110;
#1 $display("%b", po);
# 1  pi=13'b0101010011111;
#1 $display("%b", po);
# 1  pi=13'b0101010100000;
#1 $display("%b", po);
# 1  pi=13'b0101010100001;
#1 $display("%b", po);
# 1  pi=13'b0101010100010;
#1 $display("%b", po);
# 1  pi=13'b0101010100011;
#1 $display("%b", po);
# 1  pi=13'b0101010100100;
#1 $display("%b", po);
# 1  pi=13'b0101010100101;
#1 $display("%b", po);
# 1  pi=13'b0101010100110;
#1 $display("%b", po);
# 1  pi=13'b0101010100111;
#1 $display("%b", po);
# 1  pi=13'b0101010101000;
#1 $display("%b", po);
# 1  pi=13'b0101010101001;
#1 $display("%b", po);
# 1  pi=13'b0101010101010;
#1 $display("%b", po);
# 1  pi=13'b0101010101011;
#1 $display("%b", po);
# 1  pi=13'b0101010101100;
#1 $display("%b", po);
# 1  pi=13'b0101010101101;
#1 $display("%b", po);
# 1  pi=13'b0101010101110;
#1 $display("%b", po);
# 1  pi=13'b0101010101111;
#1 $display("%b", po);
# 1  pi=13'b0101010110000;
#1 $display("%b", po);
# 1  pi=13'b0101010110001;
#1 $display("%b", po);
# 1  pi=13'b0101010110010;
#1 $display("%b", po);
# 1  pi=13'b0101010110011;
#1 $display("%b", po);
# 1  pi=13'b0101010110100;
#1 $display("%b", po);
# 1  pi=13'b0101010110101;
#1 $display("%b", po);
# 1  pi=13'b0101010110110;
#1 $display("%b", po);
# 1  pi=13'b0101010110111;
#1 $display("%b", po);
# 1  pi=13'b0101010111000;
#1 $display("%b", po);
# 1  pi=13'b0101010111001;
#1 $display("%b", po);
# 1  pi=13'b0101010111010;
#1 $display("%b", po);
# 1  pi=13'b0101010111011;
#1 $display("%b", po);
# 1  pi=13'b0101010111100;
#1 $display("%b", po);
# 1  pi=13'b0101010111101;
#1 $display("%b", po);
# 1  pi=13'b0101010111110;
#1 $display("%b", po);
# 1  pi=13'b0101010111111;
#1 $display("%b", po);
# 1  pi=13'b0101011000000;
#1 $display("%b", po);
# 1  pi=13'b0101011000001;
#1 $display("%b", po);
# 1  pi=13'b0101011000010;
#1 $display("%b", po);
# 1  pi=13'b0101011000011;
#1 $display("%b", po);
# 1  pi=13'b0101011000100;
#1 $display("%b", po);
# 1  pi=13'b0101011000101;
#1 $display("%b", po);
# 1  pi=13'b0101011000110;
#1 $display("%b", po);
# 1  pi=13'b0101011000111;
#1 $display("%b", po);
# 1  pi=13'b0101011001000;
#1 $display("%b", po);
# 1  pi=13'b0101011001001;
#1 $display("%b", po);
# 1  pi=13'b0101011001010;
#1 $display("%b", po);
# 1  pi=13'b0101011001011;
#1 $display("%b", po);
# 1  pi=13'b0101011001100;
#1 $display("%b", po);
# 1  pi=13'b0101011001101;
#1 $display("%b", po);
# 1  pi=13'b0101011001110;
#1 $display("%b", po);
# 1  pi=13'b0101011001111;
#1 $display("%b", po);
# 1  pi=13'b0101011010000;
#1 $display("%b", po);
# 1  pi=13'b0101011010001;
#1 $display("%b", po);
# 1  pi=13'b0101011010010;
#1 $display("%b", po);
# 1  pi=13'b0101011010011;
#1 $display("%b", po);
# 1  pi=13'b0101011010100;
#1 $display("%b", po);
# 1  pi=13'b0101011010101;
#1 $display("%b", po);
# 1  pi=13'b0101011010110;
#1 $display("%b", po);
# 1  pi=13'b0101011010111;
#1 $display("%b", po);
# 1  pi=13'b0101011011000;
#1 $display("%b", po);
# 1  pi=13'b0101011011001;
#1 $display("%b", po);
# 1  pi=13'b0101011011010;
#1 $display("%b", po);
# 1  pi=13'b0101011011011;
#1 $display("%b", po);
# 1  pi=13'b0101011011100;
#1 $display("%b", po);
# 1  pi=13'b0101011011101;
#1 $display("%b", po);
# 1  pi=13'b0101011011110;
#1 $display("%b", po);
# 1  pi=13'b0101011011111;
#1 $display("%b", po);
# 1  pi=13'b0101011100000;
#1 $display("%b", po);
# 1  pi=13'b0101011100001;
#1 $display("%b", po);
# 1  pi=13'b0101011100010;
#1 $display("%b", po);
# 1  pi=13'b0101011100011;
#1 $display("%b", po);
# 1  pi=13'b0101011100100;
#1 $display("%b", po);
# 1  pi=13'b0101011100101;
#1 $display("%b", po);
# 1  pi=13'b0101011100110;
#1 $display("%b", po);
# 1  pi=13'b0101011100111;
#1 $display("%b", po);
# 1  pi=13'b0101011101000;
#1 $display("%b", po);
# 1  pi=13'b0101011101001;
#1 $display("%b", po);
# 1  pi=13'b0101011101010;
#1 $display("%b", po);
# 1  pi=13'b0101011101011;
#1 $display("%b", po);
# 1  pi=13'b0101011101100;
#1 $display("%b", po);
# 1  pi=13'b0101011101101;
#1 $display("%b", po);
# 1  pi=13'b0101011101110;
#1 $display("%b", po);
# 1  pi=13'b0101011101111;
#1 $display("%b", po);
# 1  pi=13'b0101011110000;
#1 $display("%b", po);
# 1  pi=13'b0101011110001;
#1 $display("%b", po);
# 1  pi=13'b0101011110010;
#1 $display("%b", po);
# 1  pi=13'b0101011110011;
#1 $display("%b", po);
# 1  pi=13'b0101011110100;
#1 $display("%b", po);
# 1  pi=13'b0101011110101;
#1 $display("%b", po);
# 1  pi=13'b0101011110110;
#1 $display("%b", po);
# 1  pi=13'b0101011110111;
#1 $display("%b", po);
# 1  pi=13'b0101011111000;
#1 $display("%b", po);
# 1  pi=13'b0101011111001;
#1 $display("%b", po);
# 1  pi=13'b0101011111010;
#1 $display("%b", po);
# 1  pi=13'b0101011111011;
#1 $display("%b", po);
# 1  pi=13'b0101011111100;
#1 $display("%b", po);
# 1  pi=13'b0101011111101;
#1 $display("%b", po);
# 1  pi=13'b0101011111110;
#1 $display("%b", po);
# 1  pi=13'b0101011111111;
#1 $display("%b", po);
# 1  pi=13'b0101100000000;
#1 $display("%b", po);
# 1  pi=13'b0101100000001;
#1 $display("%b", po);
# 1  pi=13'b0101100000010;
#1 $display("%b", po);
# 1  pi=13'b0101100000011;
#1 $display("%b", po);
# 1  pi=13'b0101100000100;
#1 $display("%b", po);
# 1  pi=13'b0101100000101;
#1 $display("%b", po);
# 1  pi=13'b0101100000110;
#1 $display("%b", po);
# 1  pi=13'b0101100000111;
#1 $display("%b", po);
# 1  pi=13'b0101100001000;
#1 $display("%b", po);
# 1  pi=13'b0101100001001;
#1 $display("%b", po);
# 1  pi=13'b0101100001010;
#1 $display("%b", po);
# 1  pi=13'b0101100001011;
#1 $display("%b", po);
# 1  pi=13'b0101100001100;
#1 $display("%b", po);
# 1  pi=13'b0101100001101;
#1 $display("%b", po);
# 1  pi=13'b0101100001110;
#1 $display("%b", po);
# 1  pi=13'b0101100001111;
#1 $display("%b", po);
# 1  pi=13'b0101100010000;
#1 $display("%b", po);
# 1  pi=13'b0101100010001;
#1 $display("%b", po);
# 1  pi=13'b0101100010010;
#1 $display("%b", po);
# 1  pi=13'b0101100010011;
#1 $display("%b", po);
# 1  pi=13'b0101100010100;
#1 $display("%b", po);
# 1  pi=13'b0101100010101;
#1 $display("%b", po);
# 1  pi=13'b0101100010110;
#1 $display("%b", po);
# 1  pi=13'b0101100010111;
#1 $display("%b", po);
# 1  pi=13'b0101100011000;
#1 $display("%b", po);
# 1  pi=13'b0101100011001;
#1 $display("%b", po);
# 1  pi=13'b0101100011010;
#1 $display("%b", po);
# 1  pi=13'b0101100011011;
#1 $display("%b", po);
# 1  pi=13'b0101100011100;
#1 $display("%b", po);
# 1  pi=13'b0101100011101;
#1 $display("%b", po);
# 1  pi=13'b0101100011110;
#1 $display("%b", po);
# 1  pi=13'b0101100011111;
#1 $display("%b", po);
# 1  pi=13'b0101100100000;
#1 $display("%b", po);
# 1  pi=13'b0101100100001;
#1 $display("%b", po);
# 1  pi=13'b0101100100010;
#1 $display("%b", po);
# 1  pi=13'b0101100100011;
#1 $display("%b", po);
# 1  pi=13'b0101100100100;
#1 $display("%b", po);
# 1  pi=13'b0101100100101;
#1 $display("%b", po);
# 1  pi=13'b0101100100110;
#1 $display("%b", po);
# 1  pi=13'b0101100100111;
#1 $display("%b", po);
# 1  pi=13'b0101100101000;
#1 $display("%b", po);
# 1  pi=13'b0101100101001;
#1 $display("%b", po);
# 1  pi=13'b0101100101010;
#1 $display("%b", po);
# 1  pi=13'b0101100101011;
#1 $display("%b", po);
# 1  pi=13'b0101100101100;
#1 $display("%b", po);
# 1  pi=13'b0101100101101;
#1 $display("%b", po);
# 1  pi=13'b0101100101110;
#1 $display("%b", po);
# 1  pi=13'b0101100101111;
#1 $display("%b", po);
# 1  pi=13'b0101100110000;
#1 $display("%b", po);
# 1  pi=13'b0101100110001;
#1 $display("%b", po);
# 1  pi=13'b0101100110010;
#1 $display("%b", po);
# 1  pi=13'b0101100110011;
#1 $display("%b", po);
# 1  pi=13'b0101100110100;
#1 $display("%b", po);
# 1  pi=13'b0101100110101;
#1 $display("%b", po);
# 1  pi=13'b0101100110110;
#1 $display("%b", po);
# 1  pi=13'b0101100110111;
#1 $display("%b", po);
# 1  pi=13'b0101100111000;
#1 $display("%b", po);
# 1  pi=13'b0101100111001;
#1 $display("%b", po);
# 1  pi=13'b0101100111010;
#1 $display("%b", po);
# 1  pi=13'b0101100111011;
#1 $display("%b", po);
# 1  pi=13'b0101100111100;
#1 $display("%b", po);
# 1  pi=13'b0101100111101;
#1 $display("%b", po);
# 1  pi=13'b0101100111110;
#1 $display("%b", po);
# 1  pi=13'b0101100111111;
#1 $display("%b", po);
# 1  pi=13'b0101101000000;
#1 $display("%b", po);
# 1  pi=13'b0101101000001;
#1 $display("%b", po);
# 1  pi=13'b0101101000010;
#1 $display("%b", po);
# 1  pi=13'b0101101000011;
#1 $display("%b", po);
# 1  pi=13'b0101101000100;
#1 $display("%b", po);
# 1  pi=13'b0101101000101;
#1 $display("%b", po);
# 1  pi=13'b0101101000110;
#1 $display("%b", po);
# 1  pi=13'b0101101000111;
#1 $display("%b", po);
# 1  pi=13'b0101101001000;
#1 $display("%b", po);
# 1  pi=13'b0101101001001;
#1 $display("%b", po);
# 1  pi=13'b0101101001010;
#1 $display("%b", po);
# 1  pi=13'b0101101001011;
#1 $display("%b", po);
# 1  pi=13'b0101101001100;
#1 $display("%b", po);
# 1  pi=13'b0101101001101;
#1 $display("%b", po);
# 1  pi=13'b0101101001110;
#1 $display("%b", po);
# 1  pi=13'b0101101001111;
#1 $display("%b", po);
# 1  pi=13'b0101101010000;
#1 $display("%b", po);
# 1  pi=13'b0101101010001;
#1 $display("%b", po);
# 1  pi=13'b0101101010010;
#1 $display("%b", po);
# 1  pi=13'b0101101010011;
#1 $display("%b", po);
# 1  pi=13'b0101101010100;
#1 $display("%b", po);
# 1  pi=13'b0101101010101;
#1 $display("%b", po);
# 1  pi=13'b0101101010110;
#1 $display("%b", po);
# 1  pi=13'b0101101010111;
#1 $display("%b", po);
# 1  pi=13'b0101101011000;
#1 $display("%b", po);
# 1  pi=13'b0101101011001;
#1 $display("%b", po);
# 1  pi=13'b0101101011010;
#1 $display("%b", po);
# 1  pi=13'b0101101011011;
#1 $display("%b", po);
# 1  pi=13'b0101101011100;
#1 $display("%b", po);
# 1  pi=13'b0101101011101;
#1 $display("%b", po);
# 1  pi=13'b0101101011110;
#1 $display("%b", po);
# 1  pi=13'b0101101011111;
#1 $display("%b", po);
# 1  pi=13'b0101101100000;
#1 $display("%b", po);
# 1  pi=13'b0101101100001;
#1 $display("%b", po);
# 1  pi=13'b0101101100010;
#1 $display("%b", po);
# 1  pi=13'b0101101100011;
#1 $display("%b", po);
# 1  pi=13'b0101101100100;
#1 $display("%b", po);
# 1  pi=13'b0101101100101;
#1 $display("%b", po);
# 1  pi=13'b0101101100110;
#1 $display("%b", po);
# 1  pi=13'b0101101100111;
#1 $display("%b", po);
# 1  pi=13'b0101101101000;
#1 $display("%b", po);
# 1  pi=13'b0101101101001;
#1 $display("%b", po);
# 1  pi=13'b0101101101010;
#1 $display("%b", po);
# 1  pi=13'b0101101101011;
#1 $display("%b", po);
# 1  pi=13'b0101101101100;
#1 $display("%b", po);
# 1  pi=13'b0101101101101;
#1 $display("%b", po);
# 1  pi=13'b0101101101110;
#1 $display("%b", po);
# 1  pi=13'b0101101101111;
#1 $display("%b", po);
# 1  pi=13'b0101101110000;
#1 $display("%b", po);
# 1  pi=13'b0101101110001;
#1 $display("%b", po);
# 1  pi=13'b0101101110010;
#1 $display("%b", po);
# 1  pi=13'b0101101110011;
#1 $display("%b", po);
# 1  pi=13'b0101101110100;
#1 $display("%b", po);
# 1  pi=13'b0101101110101;
#1 $display("%b", po);
# 1  pi=13'b0101101110110;
#1 $display("%b", po);
# 1  pi=13'b0101101110111;
#1 $display("%b", po);
# 1  pi=13'b0101101111000;
#1 $display("%b", po);
# 1  pi=13'b0101101111001;
#1 $display("%b", po);
# 1  pi=13'b0101101111010;
#1 $display("%b", po);
# 1  pi=13'b0101101111011;
#1 $display("%b", po);
# 1  pi=13'b0101101111100;
#1 $display("%b", po);
# 1  pi=13'b0101101111101;
#1 $display("%b", po);
# 1  pi=13'b0101101111110;
#1 $display("%b", po);
# 1  pi=13'b0101101111111;
#1 $display("%b", po);
# 1  pi=13'b0101110000000;
#1 $display("%b", po);
# 1  pi=13'b0101110000001;
#1 $display("%b", po);
# 1  pi=13'b0101110000010;
#1 $display("%b", po);
# 1  pi=13'b0101110000011;
#1 $display("%b", po);
# 1  pi=13'b0101110000100;
#1 $display("%b", po);
# 1  pi=13'b0101110000101;
#1 $display("%b", po);
# 1  pi=13'b0101110000110;
#1 $display("%b", po);
# 1  pi=13'b0101110000111;
#1 $display("%b", po);
# 1  pi=13'b0101110001000;
#1 $display("%b", po);
# 1  pi=13'b0101110001001;
#1 $display("%b", po);
# 1  pi=13'b0101110001010;
#1 $display("%b", po);
# 1  pi=13'b0101110001011;
#1 $display("%b", po);
# 1  pi=13'b0101110001100;
#1 $display("%b", po);
# 1  pi=13'b0101110001101;
#1 $display("%b", po);
# 1  pi=13'b0101110001110;
#1 $display("%b", po);
# 1  pi=13'b0101110001111;
#1 $display("%b", po);
# 1  pi=13'b0101110010000;
#1 $display("%b", po);
# 1  pi=13'b0101110010001;
#1 $display("%b", po);
# 1  pi=13'b0101110010010;
#1 $display("%b", po);
# 1  pi=13'b0101110010011;
#1 $display("%b", po);
# 1  pi=13'b0101110010100;
#1 $display("%b", po);
# 1  pi=13'b0101110010101;
#1 $display("%b", po);
# 1  pi=13'b0101110010110;
#1 $display("%b", po);
# 1  pi=13'b0101110010111;
#1 $display("%b", po);
# 1  pi=13'b0101110011000;
#1 $display("%b", po);
# 1  pi=13'b0101110011001;
#1 $display("%b", po);
# 1  pi=13'b0101110011010;
#1 $display("%b", po);
# 1  pi=13'b0101110011011;
#1 $display("%b", po);
# 1  pi=13'b0101110011100;
#1 $display("%b", po);
# 1  pi=13'b0101110011101;
#1 $display("%b", po);
# 1  pi=13'b0101110011110;
#1 $display("%b", po);
# 1  pi=13'b0101110011111;
#1 $display("%b", po);
# 1  pi=13'b0101110100000;
#1 $display("%b", po);
# 1  pi=13'b0101110100001;
#1 $display("%b", po);
# 1  pi=13'b0101110100010;
#1 $display("%b", po);
# 1  pi=13'b0101110100011;
#1 $display("%b", po);
# 1  pi=13'b0101110100100;
#1 $display("%b", po);
# 1  pi=13'b0101110100101;
#1 $display("%b", po);
# 1  pi=13'b0101110100110;
#1 $display("%b", po);
# 1  pi=13'b0101110100111;
#1 $display("%b", po);
# 1  pi=13'b0101110101000;
#1 $display("%b", po);
# 1  pi=13'b0101110101001;
#1 $display("%b", po);
# 1  pi=13'b0101110101010;
#1 $display("%b", po);
# 1  pi=13'b0101110101011;
#1 $display("%b", po);
# 1  pi=13'b0101110101100;
#1 $display("%b", po);
# 1  pi=13'b0101110101101;
#1 $display("%b", po);
# 1  pi=13'b0101110101110;
#1 $display("%b", po);
# 1  pi=13'b0101110101111;
#1 $display("%b", po);
# 1  pi=13'b0101110110000;
#1 $display("%b", po);
# 1  pi=13'b0101110110001;
#1 $display("%b", po);
# 1  pi=13'b0101110110010;
#1 $display("%b", po);
# 1  pi=13'b0101110110011;
#1 $display("%b", po);
# 1  pi=13'b0101110110100;
#1 $display("%b", po);
# 1  pi=13'b0101110110101;
#1 $display("%b", po);
# 1  pi=13'b0101110110110;
#1 $display("%b", po);
# 1  pi=13'b0101110110111;
#1 $display("%b", po);
# 1  pi=13'b0101110111000;
#1 $display("%b", po);
# 1  pi=13'b0101110111001;
#1 $display("%b", po);
# 1  pi=13'b0101110111010;
#1 $display("%b", po);
# 1  pi=13'b0101110111011;
#1 $display("%b", po);
# 1  pi=13'b0101110111100;
#1 $display("%b", po);
# 1  pi=13'b0101110111101;
#1 $display("%b", po);
# 1  pi=13'b0101110111110;
#1 $display("%b", po);
# 1  pi=13'b0101110111111;
#1 $display("%b", po);
# 1  pi=13'b0101111000000;
#1 $display("%b", po);
# 1  pi=13'b0101111000001;
#1 $display("%b", po);
# 1  pi=13'b0101111000010;
#1 $display("%b", po);
# 1  pi=13'b0101111000011;
#1 $display("%b", po);
# 1  pi=13'b0101111000100;
#1 $display("%b", po);
# 1  pi=13'b0101111000101;
#1 $display("%b", po);
# 1  pi=13'b0101111000110;
#1 $display("%b", po);
# 1  pi=13'b0101111000111;
#1 $display("%b", po);
# 1  pi=13'b0101111001000;
#1 $display("%b", po);
# 1  pi=13'b0101111001001;
#1 $display("%b", po);
# 1  pi=13'b0101111001010;
#1 $display("%b", po);
# 1  pi=13'b0101111001011;
#1 $display("%b", po);
# 1  pi=13'b0101111001100;
#1 $display("%b", po);
# 1  pi=13'b0101111001101;
#1 $display("%b", po);
# 1  pi=13'b0101111001110;
#1 $display("%b", po);
# 1  pi=13'b0101111001111;
#1 $display("%b", po);
# 1  pi=13'b0101111010000;
#1 $display("%b", po);
# 1  pi=13'b0101111010001;
#1 $display("%b", po);
# 1  pi=13'b0101111010010;
#1 $display("%b", po);
# 1  pi=13'b0101111010011;
#1 $display("%b", po);
# 1  pi=13'b0101111010100;
#1 $display("%b", po);
# 1  pi=13'b0101111010101;
#1 $display("%b", po);
# 1  pi=13'b0101111010110;
#1 $display("%b", po);
# 1  pi=13'b0101111010111;
#1 $display("%b", po);
# 1  pi=13'b0101111011000;
#1 $display("%b", po);
# 1  pi=13'b0101111011001;
#1 $display("%b", po);
# 1  pi=13'b0101111011010;
#1 $display("%b", po);
# 1  pi=13'b0101111011011;
#1 $display("%b", po);
# 1  pi=13'b0101111011100;
#1 $display("%b", po);
# 1  pi=13'b0101111011101;
#1 $display("%b", po);
# 1  pi=13'b0101111011110;
#1 $display("%b", po);
# 1  pi=13'b0101111011111;
#1 $display("%b", po);
# 1  pi=13'b0101111100000;
#1 $display("%b", po);
# 1  pi=13'b0101111100001;
#1 $display("%b", po);
# 1  pi=13'b0101111100010;
#1 $display("%b", po);
# 1  pi=13'b0101111100011;
#1 $display("%b", po);
# 1  pi=13'b0101111100100;
#1 $display("%b", po);
# 1  pi=13'b0101111100101;
#1 $display("%b", po);
# 1  pi=13'b0101111100110;
#1 $display("%b", po);
# 1  pi=13'b0101111100111;
#1 $display("%b", po);
# 1  pi=13'b0101111101000;
#1 $display("%b", po);
# 1  pi=13'b0101111101001;
#1 $display("%b", po);
# 1  pi=13'b0101111101010;
#1 $display("%b", po);
# 1  pi=13'b0101111101011;
#1 $display("%b", po);
# 1  pi=13'b0101111101100;
#1 $display("%b", po);
# 1  pi=13'b0101111101101;
#1 $display("%b", po);
# 1  pi=13'b0101111101110;
#1 $display("%b", po);
# 1  pi=13'b0101111101111;
#1 $display("%b", po);
# 1  pi=13'b0101111110000;
#1 $display("%b", po);
# 1  pi=13'b0101111110001;
#1 $display("%b", po);
# 1  pi=13'b0101111110010;
#1 $display("%b", po);
# 1  pi=13'b0101111110011;
#1 $display("%b", po);
# 1  pi=13'b0101111110100;
#1 $display("%b", po);
# 1  pi=13'b0101111110101;
#1 $display("%b", po);
# 1  pi=13'b0101111110110;
#1 $display("%b", po);
# 1  pi=13'b0101111110111;
#1 $display("%b", po);
# 1  pi=13'b0101111111000;
#1 $display("%b", po);
# 1  pi=13'b0101111111001;
#1 $display("%b", po);
# 1  pi=13'b0101111111010;
#1 $display("%b", po);
# 1  pi=13'b0101111111011;
#1 $display("%b", po);
# 1  pi=13'b0101111111100;
#1 $display("%b", po);
# 1  pi=13'b0101111111101;
#1 $display("%b", po);
# 1  pi=13'b0101111111110;
#1 $display("%b", po);
# 1  pi=13'b0101111111111;
#1 $display("%b", po);
# 1  pi=13'b0110000000000;
#1 $display("%b", po);
# 1  pi=13'b0110000000001;
#1 $display("%b", po);
# 1  pi=13'b0110000000010;
#1 $display("%b", po);
# 1  pi=13'b0110000000011;
#1 $display("%b", po);
# 1  pi=13'b0110000000100;
#1 $display("%b", po);
# 1  pi=13'b0110000000101;
#1 $display("%b", po);
# 1  pi=13'b0110000000110;
#1 $display("%b", po);
# 1  pi=13'b0110000000111;
#1 $display("%b", po);
# 1  pi=13'b0110000001000;
#1 $display("%b", po);
# 1  pi=13'b0110000001001;
#1 $display("%b", po);
# 1  pi=13'b0110000001010;
#1 $display("%b", po);
# 1  pi=13'b0110000001011;
#1 $display("%b", po);
# 1  pi=13'b0110000001100;
#1 $display("%b", po);
# 1  pi=13'b0110000001101;
#1 $display("%b", po);
# 1  pi=13'b0110000001110;
#1 $display("%b", po);
# 1  pi=13'b0110000001111;
#1 $display("%b", po);
# 1  pi=13'b0110000010000;
#1 $display("%b", po);
# 1  pi=13'b0110000010001;
#1 $display("%b", po);
# 1  pi=13'b0110000010010;
#1 $display("%b", po);
# 1  pi=13'b0110000010011;
#1 $display("%b", po);
# 1  pi=13'b0110000010100;
#1 $display("%b", po);
# 1  pi=13'b0110000010101;
#1 $display("%b", po);
# 1  pi=13'b0110000010110;
#1 $display("%b", po);
# 1  pi=13'b0110000010111;
#1 $display("%b", po);
# 1  pi=13'b0110000011000;
#1 $display("%b", po);
# 1  pi=13'b0110000011001;
#1 $display("%b", po);
# 1  pi=13'b0110000011010;
#1 $display("%b", po);
# 1  pi=13'b0110000011011;
#1 $display("%b", po);
# 1  pi=13'b0110000011100;
#1 $display("%b", po);
# 1  pi=13'b0110000011101;
#1 $display("%b", po);
# 1  pi=13'b0110000011110;
#1 $display("%b", po);
# 1  pi=13'b0110000011111;
#1 $display("%b", po);
# 1  pi=13'b0110000100000;
#1 $display("%b", po);
# 1  pi=13'b0110000100001;
#1 $display("%b", po);
# 1  pi=13'b0110000100010;
#1 $display("%b", po);
# 1  pi=13'b0110000100011;
#1 $display("%b", po);
# 1  pi=13'b0110000100100;
#1 $display("%b", po);
# 1  pi=13'b0110000100101;
#1 $display("%b", po);
# 1  pi=13'b0110000100110;
#1 $display("%b", po);
# 1  pi=13'b0110000100111;
#1 $display("%b", po);
# 1  pi=13'b0110000101000;
#1 $display("%b", po);
# 1  pi=13'b0110000101001;
#1 $display("%b", po);
# 1  pi=13'b0110000101010;
#1 $display("%b", po);
# 1  pi=13'b0110000101011;
#1 $display("%b", po);
# 1  pi=13'b0110000101100;
#1 $display("%b", po);
# 1  pi=13'b0110000101101;
#1 $display("%b", po);
# 1  pi=13'b0110000101110;
#1 $display("%b", po);
# 1  pi=13'b0110000101111;
#1 $display("%b", po);
# 1  pi=13'b0110000110000;
#1 $display("%b", po);
# 1  pi=13'b0110000110001;
#1 $display("%b", po);
# 1  pi=13'b0110000110010;
#1 $display("%b", po);
# 1  pi=13'b0110000110011;
#1 $display("%b", po);
# 1  pi=13'b0110000110100;
#1 $display("%b", po);
# 1  pi=13'b0110000110101;
#1 $display("%b", po);
# 1  pi=13'b0110000110110;
#1 $display("%b", po);
# 1  pi=13'b0110000110111;
#1 $display("%b", po);
# 1  pi=13'b0110000111000;
#1 $display("%b", po);
# 1  pi=13'b0110000111001;
#1 $display("%b", po);
# 1  pi=13'b0110000111010;
#1 $display("%b", po);
# 1  pi=13'b0110000111011;
#1 $display("%b", po);
# 1  pi=13'b0110000111100;
#1 $display("%b", po);
# 1  pi=13'b0110000111101;
#1 $display("%b", po);
# 1  pi=13'b0110000111110;
#1 $display("%b", po);
# 1  pi=13'b0110000111111;
#1 $display("%b", po);
# 1  pi=13'b0110001000000;
#1 $display("%b", po);
# 1  pi=13'b0110001000001;
#1 $display("%b", po);
# 1  pi=13'b0110001000010;
#1 $display("%b", po);
# 1  pi=13'b0110001000011;
#1 $display("%b", po);
# 1  pi=13'b0110001000100;
#1 $display("%b", po);
# 1  pi=13'b0110001000101;
#1 $display("%b", po);
# 1  pi=13'b0110001000110;
#1 $display("%b", po);
# 1  pi=13'b0110001000111;
#1 $display("%b", po);
# 1  pi=13'b0110001001000;
#1 $display("%b", po);
# 1  pi=13'b0110001001001;
#1 $display("%b", po);
# 1  pi=13'b0110001001010;
#1 $display("%b", po);
# 1  pi=13'b0110001001011;
#1 $display("%b", po);
# 1  pi=13'b0110001001100;
#1 $display("%b", po);
# 1  pi=13'b0110001001101;
#1 $display("%b", po);
# 1  pi=13'b0110001001110;
#1 $display("%b", po);
# 1  pi=13'b0110001001111;
#1 $display("%b", po);
# 1  pi=13'b0110001010000;
#1 $display("%b", po);
# 1  pi=13'b0110001010001;
#1 $display("%b", po);
# 1  pi=13'b0110001010010;
#1 $display("%b", po);
# 1  pi=13'b0110001010011;
#1 $display("%b", po);
# 1  pi=13'b0110001010100;
#1 $display("%b", po);
# 1  pi=13'b0110001010101;
#1 $display("%b", po);
# 1  pi=13'b0110001010110;
#1 $display("%b", po);
# 1  pi=13'b0110001010111;
#1 $display("%b", po);
# 1  pi=13'b0110001011000;
#1 $display("%b", po);
# 1  pi=13'b0110001011001;
#1 $display("%b", po);
# 1  pi=13'b0110001011010;
#1 $display("%b", po);
# 1  pi=13'b0110001011011;
#1 $display("%b", po);
# 1  pi=13'b0110001011100;
#1 $display("%b", po);
# 1  pi=13'b0110001011101;
#1 $display("%b", po);
# 1  pi=13'b0110001011110;
#1 $display("%b", po);
# 1  pi=13'b0110001011111;
#1 $display("%b", po);
# 1  pi=13'b0110001100000;
#1 $display("%b", po);
# 1  pi=13'b0110001100001;
#1 $display("%b", po);
# 1  pi=13'b0110001100010;
#1 $display("%b", po);
# 1  pi=13'b0110001100011;
#1 $display("%b", po);
# 1  pi=13'b0110001100100;
#1 $display("%b", po);
# 1  pi=13'b0110001100101;
#1 $display("%b", po);
# 1  pi=13'b0110001100110;
#1 $display("%b", po);
# 1  pi=13'b0110001100111;
#1 $display("%b", po);
# 1  pi=13'b0110001101000;
#1 $display("%b", po);
# 1  pi=13'b0110001101001;
#1 $display("%b", po);
# 1  pi=13'b0110001101010;
#1 $display("%b", po);
# 1  pi=13'b0110001101011;
#1 $display("%b", po);
# 1  pi=13'b0110001101100;
#1 $display("%b", po);
# 1  pi=13'b0110001101101;
#1 $display("%b", po);
# 1  pi=13'b0110001101110;
#1 $display("%b", po);
# 1  pi=13'b0110001101111;
#1 $display("%b", po);
# 1  pi=13'b0110001110000;
#1 $display("%b", po);
# 1  pi=13'b0110001110001;
#1 $display("%b", po);
# 1  pi=13'b0110001110010;
#1 $display("%b", po);
# 1  pi=13'b0110001110011;
#1 $display("%b", po);
# 1  pi=13'b0110001110100;
#1 $display("%b", po);
# 1  pi=13'b0110001110101;
#1 $display("%b", po);
# 1  pi=13'b0110001110110;
#1 $display("%b", po);
# 1  pi=13'b0110001110111;
#1 $display("%b", po);
# 1  pi=13'b0110001111000;
#1 $display("%b", po);
# 1  pi=13'b0110001111001;
#1 $display("%b", po);
# 1  pi=13'b0110001111010;
#1 $display("%b", po);
# 1  pi=13'b0110001111011;
#1 $display("%b", po);
# 1  pi=13'b0110001111100;
#1 $display("%b", po);
# 1  pi=13'b0110001111101;
#1 $display("%b", po);
# 1  pi=13'b0110001111110;
#1 $display("%b", po);
# 1  pi=13'b0110001111111;
#1 $display("%b", po);
# 1  pi=13'b0110010000000;
#1 $display("%b", po);
# 1  pi=13'b0110010000001;
#1 $display("%b", po);
# 1  pi=13'b0110010000010;
#1 $display("%b", po);
# 1  pi=13'b0110010000011;
#1 $display("%b", po);
# 1  pi=13'b0110010000100;
#1 $display("%b", po);
# 1  pi=13'b0110010000101;
#1 $display("%b", po);
# 1  pi=13'b0110010000110;
#1 $display("%b", po);
# 1  pi=13'b0110010000111;
#1 $display("%b", po);
# 1  pi=13'b0110010001000;
#1 $display("%b", po);
# 1  pi=13'b0110010001001;
#1 $display("%b", po);
# 1  pi=13'b0110010001010;
#1 $display("%b", po);
# 1  pi=13'b0110010001011;
#1 $display("%b", po);
# 1  pi=13'b0110010001100;
#1 $display("%b", po);
# 1  pi=13'b0110010001101;
#1 $display("%b", po);
# 1  pi=13'b0110010001110;
#1 $display("%b", po);
# 1  pi=13'b0110010001111;
#1 $display("%b", po);
# 1  pi=13'b0110010010000;
#1 $display("%b", po);
# 1  pi=13'b0110010010001;
#1 $display("%b", po);
# 1  pi=13'b0110010010010;
#1 $display("%b", po);
# 1  pi=13'b0110010010011;
#1 $display("%b", po);
# 1  pi=13'b0110010010100;
#1 $display("%b", po);
# 1  pi=13'b0110010010101;
#1 $display("%b", po);
# 1  pi=13'b0110010010110;
#1 $display("%b", po);
# 1  pi=13'b0110010010111;
#1 $display("%b", po);
# 1  pi=13'b0110010011000;
#1 $display("%b", po);
# 1  pi=13'b0110010011001;
#1 $display("%b", po);
# 1  pi=13'b0110010011010;
#1 $display("%b", po);
# 1  pi=13'b0110010011011;
#1 $display("%b", po);
# 1  pi=13'b0110010011100;
#1 $display("%b", po);
# 1  pi=13'b0110010011101;
#1 $display("%b", po);
# 1  pi=13'b0110010011110;
#1 $display("%b", po);
# 1  pi=13'b0110010011111;
#1 $display("%b", po);
# 1  pi=13'b0110010100000;
#1 $display("%b", po);
# 1  pi=13'b0110010100001;
#1 $display("%b", po);
# 1  pi=13'b0110010100010;
#1 $display("%b", po);
# 1  pi=13'b0110010100011;
#1 $display("%b", po);
# 1  pi=13'b0110010100100;
#1 $display("%b", po);
# 1  pi=13'b0110010100101;
#1 $display("%b", po);
# 1  pi=13'b0110010100110;
#1 $display("%b", po);
# 1  pi=13'b0110010100111;
#1 $display("%b", po);
# 1  pi=13'b0110010101000;
#1 $display("%b", po);
# 1  pi=13'b0110010101001;
#1 $display("%b", po);
# 1  pi=13'b0110010101010;
#1 $display("%b", po);
# 1  pi=13'b0110010101011;
#1 $display("%b", po);
# 1  pi=13'b0110010101100;
#1 $display("%b", po);
# 1  pi=13'b0110010101101;
#1 $display("%b", po);
# 1  pi=13'b0110010101110;
#1 $display("%b", po);
# 1  pi=13'b0110010101111;
#1 $display("%b", po);
# 1  pi=13'b0110010110000;
#1 $display("%b", po);
# 1  pi=13'b0110010110001;
#1 $display("%b", po);
# 1  pi=13'b0110010110010;
#1 $display("%b", po);
# 1  pi=13'b0110010110011;
#1 $display("%b", po);
# 1  pi=13'b0110010110100;
#1 $display("%b", po);
# 1  pi=13'b0110010110101;
#1 $display("%b", po);
# 1  pi=13'b0110010110110;
#1 $display("%b", po);
# 1  pi=13'b0110010110111;
#1 $display("%b", po);
# 1  pi=13'b0110010111000;
#1 $display("%b", po);
# 1  pi=13'b0110010111001;
#1 $display("%b", po);
# 1  pi=13'b0110010111010;
#1 $display("%b", po);
# 1  pi=13'b0110010111011;
#1 $display("%b", po);
# 1  pi=13'b0110010111100;
#1 $display("%b", po);
# 1  pi=13'b0110010111101;
#1 $display("%b", po);
# 1  pi=13'b0110010111110;
#1 $display("%b", po);
# 1  pi=13'b0110010111111;
#1 $display("%b", po);
# 1  pi=13'b0110011000000;
#1 $display("%b", po);
# 1  pi=13'b0110011000001;
#1 $display("%b", po);
# 1  pi=13'b0110011000010;
#1 $display("%b", po);
# 1  pi=13'b0110011000011;
#1 $display("%b", po);
# 1  pi=13'b0110011000100;
#1 $display("%b", po);
# 1  pi=13'b0110011000101;
#1 $display("%b", po);
# 1  pi=13'b0110011000110;
#1 $display("%b", po);
# 1  pi=13'b0110011000111;
#1 $display("%b", po);
# 1  pi=13'b0110011001000;
#1 $display("%b", po);
# 1  pi=13'b0110011001001;
#1 $display("%b", po);
# 1  pi=13'b0110011001010;
#1 $display("%b", po);
# 1  pi=13'b0110011001011;
#1 $display("%b", po);
# 1  pi=13'b0110011001100;
#1 $display("%b", po);
# 1  pi=13'b0110011001101;
#1 $display("%b", po);
# 1  pi=13'b0110011001110;
#1 $display("%b", po);
# 1  pi=13'b0110011001111;
#1 $display("%b", po);
# 1  pi=13'b0110011010000;
#1 $display("%b", po);
# 1  pi=13'b0110011010001;
#1 $display("%b", po);
# 1  pi=13'b0110011010010;
#1 $display("%b", po);
# 1  pi=13'b0110011010011;
#1 $display("%b", po);
# 1  pi=13'b0110011010100;
#1 $display("%b", po);
# 1  pi=13'b0110011010101;
#1 $display("%b", po);
# 1  pi=13'b0110011010110;
#1 $display("%b", po);
# 1  pi=13'b0110011010111;
#1 $display("%b", po);
# 1  pi=13'b0110011011000;
#1 $display("%b", po);
# 1  pi=13'b0110011011001;
#1 $display("%b", po);
# 1  pi=13'b0110011011010;
#1 $display("%b", po);
# 1  pi=13'b0110011011011;
#1 $display("%b", po);
# 1  pi=13'b0110011011100;
#1 $display("%b", po);
# 1  pi=13'b0110011011101;
#1 $display("%b", po);
# 1  pi=13'b0110011011110;
#1 $display("%b", po);
# 1  pi=13'b0110011011111;
#1 $display("%b", po);
# 1  pi=13'b0110011100000;
#1 $display("%b", po);
# 1  pi=13'b0110011100001;
#1 $display("%b", po);
# 1  pi=13'b0110011100010;
#1 $display("%b", po);
# 1  pi=13'b0110011100011;
#1 $display("%b", po);
# 1  pi=13'b0110011100100;
#1 $display("%b", po);
# 1  pi=13'b0110011100101;
#1 $display("%b", po);
# 1  pi=13'b0110011100110;
#1 $display("%b", po);
# 1  pi=13'b0110011100111;
#1 $display("%b", po);
# 1  pi=13'b0110011101000;
#1 $display("%b", po);
# 1  pi=13'b0110011101001;
#1 $display("%b", po);
# 1  pi=13'b0110011101010;
#1 $display("%b", po);
# 1  pi=13'b0110011101011;
#1 $display("%b", po);
# 1  pi=13'b0110011101100;
#1 $display("%b", po);
# 1  pi=13'b0110011101101;
#1 $display("%b", po);
# 1  pi=13'b0110011101110;
#1 $display("%b", po);
# 1  pi=13'b0110011101111;
#1 $display("%b", po);
# 1  pi=13'b0110011110000;
#1 $display("%b", po);
# 1  pi=13'b0110011110001;
#1 $display("%b", po);
# 1  pi=13'b0110011110010;
#1 $display("%b", po);
# 1  pi=13'b0110011110011;
#1 $display("%b", po);
# 1  pi=13'b0110011110100;
#1 $display("%b", po);
# 1  pi=13'b0110011110101;
#1 $display("%b", po);
# 1  pi=13'b0110011110110;
#1 $display("%b", po);
# 1  pi=13'b0110011110111;
#1 $display("%b", po);
# 1  pi=13'b0110011111000;
#1 $display("%b", po);
# 1  pi=13'b0110011111001;
#1 $display("%b", po);
# 1  pi=13'b0110011111010;
#1 $display("%b", po);
# 1  pi=13'b0110011111011;
#1 $display("%b", po);
# 1  pi=13'b0110011111100;
#1 $display("%b", po);
# 1  pi=13'b0110011111101;
#1 $display("%b", po);
# 1  pi=13'b0110011111110;
#1 $display("%b", po);
# 1  pi=13'b0110011111111;
#1 $display("%b", po);
# 1  pi=13'b0110100000000;
#1 $display("%b", po);
# 1  pi=13'b0110100000001;
#1 $display("%b", po);
# 1  pi=13'b0110100000010;
#1 $display("%b", po);
# 1  pi=13'b0110100000011;
#1 $display("%b", po);
# 1  pi=13'b0110100000100;
#1 $display("%b", po);
# 1  pi=13'b0110100000101;
#1 $display("%b", po);
# 1  pi=13'b0110100000110;
#1 $display("%b", po);
# 1  pi=13'b0110100000111;
#1 $display("%b", po);
# 1  pi=13'b0110100001000;
#1 $display("%b", po);
# 1  pi=13'b0110100001001;
#1 $display("%b", po);
# 1  pi=13'b0110100001010;
#1 $display("%b", po);
# 1  pi=13'b0110100001011;
#1 $display("%b", po);
# 1  pi=13'b0110100001100;
#1 $display("%b", po);
# 1  pi=13'b0110100001101;
#1 $display("%b", po);
# 1  pi=13'b0110100001110;
#1 $display("%b", po);
# 1  pi=13'b0110100001111;
#1 $display("%b", po);
# 1  pi=13'b0110100010000;
#1 $display("%b", po);
# 1  pi=13'b0110100010001;
#1 $display("%b", po);
# 1  pi=13'b0110100010010;
#1 $display("%b", po);
# 1  pi=13'b0110100010011;
#1 $display("%b", po);
# 1  pi=13'b0110100010100;
#1 $display("%b", po);
# 1  pi=13'b0110100010101;
#1 $display("%b", po);
# 1  pi=13'b0110100010110;
#1 $display("%b", po);
# 1  pi=13'b0110100010111;
#1 $display("%b", po);
# 1  pi=13'b0110100011000;
#1 $display("%b", po);
# 1  pi=13'b0110100011001;
#1 $display("%b", po);
# 1  pi=13'b0110100011010;
#1 $display("%b", po);
# 1  pi=13'b0110100011011;
#1 $display("%b", po);
# 1  pi=13'b0110100011100;
#1 $display("%b", po);
# 1  pi=13'b0110100011101;
#1 $display("%b", po);
# 1  pi=13'b0110100011110;
#1 $display("%b", po);
# 1  pi=13'b0110100011111;
#1 $display("%b", po);
# 1  pi=13'b0110100100000;
#1 $display("%b", po);
# 1  pi=13'b0110100100001;
#1 $display("%b", po);
# 1  pi=13'b0110100100010;
#1 $display("%b", po);
# 1  pi=13'b0110100100011;
#1 $display("%b", po);
# 1  pi=13'b0110100100100;
#1 $display("%b", po);
# 1  pi=13'b0110100100101;
#1 $display("%b", po);
# 1  pi=13'b0110100100110;
#1 $display("%b", po);
# 1  pi=13'b0110100100111;
#1 $display("%b", po);
# 1  pi=13'b0110100101000;
#1 $display("%b", po);
# 1  pi=13'b0110100101001;
#1 $display("%b", po);
# 1  pi=13'b0110100101010;
#1 $display("%b", po);
# 1  pi=13'b0110100101011;
#1 $display("%b", po);
# 1  pi=13'b0110100101100;
#1 $display("%b", po);
# 1  pi=13'b0110100101101;
#1 $display("%b", po);
# 1  pi=13'b0110100101110;
#1 $display("%b", po);
# 1  pi=13'b0110100101111;
#1 $display("%b", po);
# 1  pi=13'b0110100110000;
#1 $display("%b", po);
# 1  pi=13'b0110100110001;
#1 $display("%b", po);
# 1  pi=13'b0110100110010;
#1 $display("%b", po);
# 1  pi=13'b0110100110011;
#1 $display("%b", po);
# 1  pi=13'b0110100110100;
#1 $display("%b", po);
# 1  pi=13'b0110100110101;
#1 $display("%b", po);
# 1  pi=13'b0110100110110;
#1 $display("%b", po);
# 1  pi=13'b0110100110111;
#1 $display("%b", po);
# 1  pi=13'b0110100111000;
#1 $display("%b", po);
# 1  pi=13'b0110100111001;
#1 $display("%b", po);
# 1  pi=13'b0110100111010;
#1 $display("%b", po);
# 1  pi=13'b0110100111011;
#1 $display("%b", po);
# 1  pi=13'b0110100111100;
#1 $display("%b", po);
# 1  pi=13'b0110100111101;
#1 $display("%b", po);
# 1  pi=13'b0110100111110;
#1 $display("%b", po);
# 1  pi=13'b0110100111111;
#1 $display("%b", po);
# 1  pi=13'b0110101000000;
#1 $display("%b", po);
# 1  pi=13'b0110101000001;
#1 $display("%b", po);
# 1  pi=13'b0110101000010;
#1 $display("%b", po);
# 1  pi=13'b0110101000011;
#1 $display("%b", po);
# 1  pi=13'b0110101000100;
#1 $display("%b", po);
# 1  pi=13'b0110101000101;
#1 $display("%b", po);
# 1  pi=13'b0110101000110;
#1 $display("%b", po);
# 1  pi=13'b0110101000111;
#1 $display("%b", po);
# 1  pi=13'b0110101001000;
#1 $display("%b", po);
# 1  pi=13'b0110101001001;
#1 $display("%b", po);
# 1  pi=13'b0110101001010;
#1 $display("%b", po);
# 1  pi=13'b0110101001011;
#1 $display("%b", po);
# 1  pi=13'b0110101001100;
#1 $display("%b", po);
# 1  pi=13'b0110101001101;
#1 $display("%b", po);
# 1  pi=13'b0110101001110;
#1 $display("%b", po);
# 1  pi=13'b0110101001111;
#1 $display("%b", po);
# 1  pi=13'b0110101010000;
#1 $display("%b", po);
# 1  pi=13'b0110101010001;
#1 $display("%b", po);
# 1  pi=13'b0110101010010;
#1 $display("%b", po);
# 1  pi=13'b0110101010011;
#1 $display("%b", po);
# 1  pi=13'b0110101010100;
#1 $display("%b", po);
# 1  pi=13'b0110101010101;
#1 $display("%b", po);
# 1  pi=13'b0110101010110;
#1 $display("%b", po);
# 1  pi=13'b0110101010111;
#1 $display("%b", po);
# 1  pi=13'b0110101011000;
#1 $display("%b", po);
# 1  pi=13'b0110101011001;
#1 $display("%b", po);
# 1  pi=13'b0110101011010;
#1 $display("%b", po);
# 1  pi=13'b0110101011011;
#1 $display("%b", po);
# 1  pi=13'b0110101011100;
#1 $display("%b", po);
# 1  pi=13'b0110101011101;
#1 $display("%b", po);
# 1  pi=13'b0110101011110;
#1 $display("%b", po);
# 1  pi=13'b0110101011111;
#1 $display("%b", po);
# 1  pi=13'b0110101100000;
#1 $display("%b", po);
# 1  pi=13'b0110101100001;
#1 $display("%b", po);
# 1  pi=13'b0110101100010;
#1 $display("%b", po);
# 1  pi=13'b0110101100011;
#1 $display("%b", po);
# 1  pi=13'b0110101100100;
#1 $display("%b", po);
# 1  pi=13'b0110101100101;
#1 $display("%b", po);
# 1  pi=13'b0110101100110;
#1 $display("%b", po);
# 1  pi=13'b0110101100111;
#1 $display("%b", po);
# 1  pi=13'b0110101101000;
#1 $display("%b", po);
# 1  pi=13'b0110101101001;
#1 $display("%b", po);
# 1  pi=13'b0110101101010;
#1 $display("%b", po);
# 1  pi=13'b0110101101011;
#1 $display("%b", po);
# 1  pi=13'b0110101101100;
#1 $display("%b", po);
# 1  pi=13'b0110101101101;
#1 $display("%b", po);
# 1  pi=13'b0110101101110;
#1 $display("%b", po);
# 1  pi=13'b0110101101111;
#1 $display("%b", po);
# 1  pi=13'b0110101110000;
#1 $display("%b", po);
# 1  pi=13'b0110101110001;
#1 $display("%b", po);
# 1  pi=13'b0110101110010;
#1 $display("%b", po);
# 1  pi=13'b0110101110011;
#1 $display("%b", po);
# 1  pi=13'b0110101110100;
#1 $display("%b", po);
# 1  pi=13'b0110101110101;
#1 $display("%b", po);
# 1  pi=13'b0110101110110;
#1 $display("%b", po);
# 1  pi=13'b0110101110111;
#1 $display("%b", po);
# 1  pi=13'b0110101111000;
#1 $display("%b", po);
# 1  pi=13'b0110101111001;
#1 $display("%b", po);
# 1  pi=13'b0110101111010;
#1 $display("%b", po);
# 1  pi=13'b0110101111011;
#1 $display("%b", po);
# 1  pi=13'b0110101111100;
#1 $display("%b", po);
# 1  pi=13'b0110101111101;
#1 $display("%b", po);
# 1  pi=13'b0110101111110;
#1 $display("%b", po);
# 1  pi=13'b0110101111111;
#1 $display("%b", po);
# 1  pi=13'b0110110000000;
#1 $display("%b", po);
# 1  pi=13'b0110110000001;
#1 $display("%b", po);
# 1  pi=13'b0110110000010;
#1 $display("%b", po);
# 1  pi=13'b0110110000011;
#1 $display("%b", po);
# 1  pi=13'b0110110000100;
#1 $display("%b", po);
# 1  pi=13'b0110110000101;
#1 $display("%b", po);
# 1  pi=13'b0110110000110;
#1 $display("%b", po);
# 1  pi=13'b0110110000111;
#1 $display("%b", po);
# 1  pi=13'b0110110001000;
#1 $display("%b", po);
# 1  pi=13'b0110110001001;
#1 $display("%b", po);
# 1  pi=13'b0110110001010;
#1 $display("%b", po);
# 1  pi=13'b0110110001011;
#1 $display("%b", po);
# 1  pi=13'b0110110001100;
#1 $display("%b", po);
# 1  pi=13'b0110110001101;
#1 $display("%b", po);
# 1  pi=13'b0110110001110;
#1 $display("%b", po);
# 1  pi=13'b0110110001111;
#1 $display("%b", po);
# 1  pi=13'b0110110010000;
#1 $display("%b", po);
# 1  pi=13'b0110110010001;
#1 $display("%b", po);
# 1  pi=13'b0110110010010;
#1 $display("%b", po);
# 1  pi=13'b0110110010011;
#1 $display("%b", po);
# 1  pi=13'b0110110010100;
#1 $display("%b", po);
# 1  pi=13'b0110110010101;
#1 $display("%b", po);
# 1  pi=13'b0110110010110;
#1 $display("%b", po);
# 1  pi=13'b0110110010111;
#1 $display("%b", po);
# 1  pi=13'b0110110011000;
#1 $display("%b", po);
# 1  pi=13'b0110110011001;
#1 $display("%b", po);
# 1  pi=13'b0110110011010;
#1 $display("%b", po);
# 1  pi=13'b0110110011011;
#1 $display("%b", po);
# 1  pi=13'b0110110011100;
#1 $display("%b", po);
# 1  pi=13'b0110110011101;
#1 $display("%b", po);
# 1  pi=13'b0110110011110;
#1 $display("%b", po);
# 1  pi=13'b0110110011111;
#1 $display("%b", po);
# 1  pi=13'b0110110100000;
#1 $display("%b", po);
# 1  pi=13'b0110110100001;
#1 $display("%b", po);
# 1  pi=13'b0110110100010;
#1 $display("%b", po);
# 1  pi=13'b0110110100011;
#1 $display("%b", po);
# 1  pi=13'b0110110100100;
#1 $display("%b", po);
# 1  pi=13'b0110110100101;
#1 $display("%b", po);
# 1  pi=13'b0110110100110;
#1 $display("%b", po);
# 1  pi=13'b0110110100111;
#1 $display("%b", po);
# 1  pi=13'b0110110101000;
#1 $display("%b", po);
# 1  pi=13'b0110110101001;
#1 $display("%b", po);
# 1  pi=13'b0110110101010;
#1 $display("%b", po);
# 1  pi=13'b0110110101011;
#1 $display("%b", po);
# 1  pi=13'b0110110101100;
#1 $display("%b", po);
# 1  pi=13'b0110110101101;
#1 $display("%b", po);
# 1  pi=13'b0110110101110;
#1 $display("%b", po);
# 1  pi=13'b0110110101111;
#1 $display("%b", po);
# 1  pi=13'b0110110110000;
#1 $display("%b", po);
# 1  pi=13'b0110110110001;
#1 $display("%b", po);
# 1  pi=13'b0110110110010;
#1 $display("%b", po);
# 1  pi=13'b0110110110011;
#1 $display("%b", po);
# 1  pi=13'b0110110110100;
#1 $display("%b", po);
# 1  pi=13'b0110110110101;
#1 $display("%b", po);
# 1  pi=13'b0110110110110;
#1 $display("%b", po);
# 1  pi=13'b0110110110111;
#1 $display("%b", po);
# 1  pi=13'b0110110111000;
#1 $display("%b", po);
# 1  pi=13'b0110110111001;
#1 $display("%b", po);
# 1  pi=13'b0110110111010;
#1 $display("%b", po);
# 1  pi=13'b0110110111011;
#1 $display("%b", po);
# 1  pi=13'b0110110111100;
#1 $display("%b", po);
# 1  pi=13'b0110110111101;
#1 $display("%b", po);
# 1  pi=13'b0110110111110;
#1 $display("%b", po);
# 1  pi=13'b0110110111111;
#1 $display("%b", po);
# 1  pi=13'b0110111000000;
#1 $display("%b", po);
# 1  pi=13'b0110111000001;
#1 $display("%b", po);
# 1  pi=13'b0110111000010;
#1 $display("%b", po);
# 1  pi=13'b0110111000011;
#1 $display("%b", po);
# 1  pi=13'b0110111000100;
#1 $display("%b", po);
# 1  pi=13'b0110111000101;
#1 $display("%b", po);
# 1  pi=13'b0110111000110;
#1 $display("%b", po);
# 1  pi=13'b0110111000111;
#1 $display("%b", po);
# 1  pi=13'b0110111001000;
#1 $display("%b", po);
# 1  pi=13'b0110111001001;
#1 $display("%b", po);
# 1  pi=13'b0110111001010;
#1 $display("%b", po);
# 1  pi=13'b0110111001011;
#1 $display("%b", po);
# 1  pi=13'b0110111001100;
#1 $display("%b", po);
# 1  pi=13'b0110111001101;
#1 $display("%b", po);
# 1  pi=13'b0110111001110;
#1 $display("%b", po);
# 1  pi=13'b0110111001111;
#1 $display("%b", po);
# 1  pi=13'b0110111010000;
#1 $display("%b", po);
# 1  pi=13'b0110111010001;
#1 $display("%b", po);
# 1  pi=13'b0110111010010;
#1 $display("%b", po);
# 1  pi=13'b0110111010011;
#1 $display("%b", po);
# 1  pi=13'b0110111010100;
#1 $display("%b", po);
# 1  pi=13'b0110111010101;
#1 $display("%b", po);
# 1  pi=13'b0110111010110;
#1 $display("%b", po);
# 1  pi=13'b0110111010111;
#1 $display("%b", po);
# 1  pi=13'b0110111011000;
#1 $display("%b", po);
# 1  pi=13'b0110111011001;
#1 $display("%b", po);
# 1  pi=13'b0110111011010;
#1 $display("%b", po);
# 1  pi=13'b0110111011011;
#1 $display("%b", po);
# 1  pi=13'b0110111011100;
#1 $display("%b", po);
# 1  pi=13'b0110111011101;
#1 $display("%b", po);
# 1  pi=13'b0110111011110;
#1 $display("%b", po);
# 1  pi=13'b0110111011111;
#1 $display("%b", po);
# 1  pi=13'b0110111100000;
#1 $display("%b", po);
# 1  pi=13'b0110111100001;
#1 $display("%b", po);
# 1  pi=13'b0110111100010;
#1 $display("%b", po);
# 1  pi=13'b0110111100011;
#1 $display("%b", po);
# 1  pi=13'b0110111100100;
#1 $display("%b", po);
# 1  pi=13'b0110111100101;
#1 $display("%b", po);
# 1  pi=13'b0110111100110;
#1 $display("%b", po);
# 1  pi=13'b0110111100111;
#1 $display("%b", po);
# 1  pi=13'b0110111101000;
#1 $display("%b", po);
# 1  pi=13'b0110111101001;
#1 $display("%b", po);
# 1  pi=13'b0110111101010;
#1 $display("%b", po);
# 1  pi=13'b0110111101011;
#1 $display("%b", po);
# 1  pi=13'b0110111101100;
#1 $display("%b", po);
# 1  pi=13'b0110111101101;
#1 $display("%b", po);
# 1  pi=13'b0110111101110;
#1 $display("%b", po);
# 1  pi=13'b0110111101111;
#1 $display("%b", po);
# 1  pi=13'b0110111110000;
#1 $display("%b", po);
# 1  pi=13'b0110111110001;
#1 $display("%b", po);
# 1  pi=13'b0110111110010;
#1 $display("%b", po);
# 1  pi=13'b0110111110011;
#1 $display("%b", po);
# 1  pi=13'b0110111110100;
#1 $display("%b", po);
# 1  pi=13'b0110111110101;
#1 $display("%b", po);
# 1  pi=13'b0110111110110;
#1 $display("%b", po);
# 1  pi=13'b0110111110111;
#1 $display("%b", po);
# 1  pi=13'b0110111111000;
#1 $display("%b", po);
# 1  pi=13'b0110111111001;
#1 $display("%b", po);
# 1  pi=13'b0110111111010;
#1 $display("%b", po);
# 1  pi=13'b0110111111011;
#1 $display("%b", po);
# 1  pi=13'b0110111111100;
#1 $display("%b", po);
# 1  pi=13'b0110111111101;
#1 $display("%b", po);
# 1  pi=13'b0110111111110;
#1 $display("%b", po);
# 1  pi=13'b0110111111111;
#1 $display("%b", po);
# 1  pi=13'b0111000000000;
#1 $display("%b", po);
# 1  pi=13'b0111000000001;
#1 $display("%b", po);
# 1  pi=13'b0111000000010;
#1 $display("%b", po);
# 1  pi=13'b0111000000011;
#1 $display("%b", po);
# 1  pi=13'b0111000000100;
#1 $display("%b", po);
# 1  pi=13'b0111000000101;
#1 $display("%b", po);
# 1  pi=13'b0111000000110;
#1 $display("%b", po);
# 1  pi=13'b0111000000111;
#1 $display("%b", po);
# 1  pi=13'b0111000001000;
#1 $display("%b", po);
# 1  pi=13'b0111000001001;
#1 $display("%b", po);
# 1  pi=13'b0111000001010;
#1 $display("%b", po);
# 1  pi=13'b0111000001011;
#1 $display("%b", po);
# 1  pi=13'b0111000001100;
#1 $display("%b", po);
# 1  pi=13'b0111000001101;
#1 $display("%b", po);
# 1  pi=13'b0111000001110;
#1 $display("%b", po);
# 1  pi=13'b0111000001111;
#1 $display("%b", po);
# 1  pi=13'b0111000010000;
#1 $display("%b", po);
# 1  pi=13'b0111000010001;
#1 $display("%b", po);
# 1  pi=13'b0111000010010;
#1 $display("%b", po);
# 1  pi=13'b0111000010011;
#1 $display("%b", po);
# 1  pi=13'b0111000010100;
#1 $display("%b", po);
# 1  pi=13'b0111000010101;
#1 $display("%b", po);
# 1  pi=13'b0111000010110;
#1 $display("%b", po);
# 1  pi=13'b0111000010111;
#1 $display("%b", po);
# 1  pi=13'b0111000011000;
#1 $display("%b", po);
# 1  pi=13'b0111000011001;
#1 $display("%b", po);
# 1  pi=13'b0111000011010;
#1 $display("%b", po);
# 1  pi=13'b0111000011011;
#1 $display("%b", po);
# 1  pi=13'b0111000011100;
#1 $display("%b", po);
# 1  pi=13'b0111000011101;
#1 $display("%b", po);
# 1  pi=13'b0111000011110;
#1 $display("%b", po);
# 1  pi=13'b0111000011111;
#1 $display("%b", po);
# 1  pi=13'b0111000100000;
#1 $display("%b", po);
# 1  pi=13'b0111000100001;
#1 $display("%b", po);
# 1  pi=13'b0111000100010;
#1 $display("%b", po);
# 1  pi=13'b0111000100011;
#1 $display("%b", po);
# 1  pi=13'b0111000100100;
#1 $display("%b", po);
# 1  pi=13'b0111000100101;
#1 $display("%b", po);
# 1  pi=13'b0111000100110;
#1 $display("%b", po);
# 1  pi=13'b0111000100111;
#1 $display("%b", po);
# 1  pi=13'b0111000101000;
#1 $display("%b", po);
# 1  pi=13'b0111000101001;
#1 $display("%b", po);
# 1  pi=13'b0111000101010;
#1 $display("%b", po);
# 1  pi=13'b0111000101011;
#1 $display("%b", po);
# 1  pi=13'b0111000101100;
#1 $display("%b", po);
# 1  pi=13'b0111000101101;
#1 $display("%b", po);
# 1  pi=13'b0111000101110;
#1 $display("%b", po);
# 1  pi=13'b0111000101111;
#1 $display("%b", po);
# 1  pi=13'b0111000110000;
#1 $display("%b", po);
# 1  pi=13'b0111000110001;
#1 $display("%b", po);
# 1  pi=13'b0111000110010;
#1 $display("%b", po);
# 1  pi=13'b0111000110011;
#1 $display("%b", po);
# 1  pi=13'b0111000110100;
#1 $display("%b", po);
# 1  pi=13'b0111000110101;
#1 $display("%b", po);
# 1  pi=13'b0111000110110;
#1 $display("%b", po);
# 1  pi=13'b0111000110111;
#1 $display("%b", po);
# 1  pi=13'b0111000111000;
#1 $display("%b", po);
# 1  pi=13'b0111000111001;
#1 $display("%b", po);
# 1  pi=13'b0111000111010;
#1 $display("%b", po);
# 1  pi=13'b0111000111011;
#1 $display("%b", po);
# 1  pi=13'b0111000111100;
#1 $display("%b", po);
# 1  pi=13'b0111000111101;
#1 $display("%b", po);
# 1  pi=13'b0111000111110;
#1 $display("%b", po);
# 1  pi=13'b0111000111111;
#1 $display("%b", po);
# 1  pi=13'b0111001000000;
#1 $display("%b", po);
# 1  pi=13'b0111001000001;
#1 $display("%b", po);
# 1  pi=13'b0111001000010;
#1 $display("%b", po);
# 1  pi=13'b0111001000011;
#1 $display("%b", po);
# 1  pi=13'b0111001000100;
#1 $display("%b", po);
# 1  pi=13'b0111001000101;
#1 $display("%b", po);
# 1  pi=13'b0111001000110;
#1 $display("%b", po);
# 1  pi=13'b0111001000111;
#1 $display("%b", po);
# 1  pi=13'b0111001001000;
#1 $display("%b", po);
# 1  pi=13'b0111001001001;
#1 $display("%b", po);
# 1  pi=13'b0111001001010;
#1 $display("%b", po);
# 1  pi=13'b0111001001011;
#1 $display("%b", po);
# 1  pi=13'b0111001001100;
#1 $display("%b", po);
# 1  pi=13'b0111001001101;
#1 $display("%b", po);
# 1  pi=13'b0111001001110;
#1 $display("%b", po);
# 1  pi=13'b0111001001111;
#1 $display("%b", po);
# 1  pi=13'b0111001010000;
#1 $display("%b", po);
# 1  pi=13'b0111001010001;
#1 $display("%b", po);
# 1  pi=13'b0111001010010;
#1 $display("%b", po);
# 1  pi=13'b0111001010011;
#1 $display("%b", po);
# 1  pi=13'b0111001010100;
#1 $display("%b", po);
# 1  pi=13'b0111001010101;
#1 $display("%b", po);
# 1  pi=13'b0111001010110;
#1 $display("%b", po);
# 1  pi=13'b0111001010111;
#1 $display("%b", po);
# 1  pi=13'b0111001011000;
#1 $display("%b", po);
# 1  pi=13'b0111001011001;
#1 $display("%b", po);
# 1  pi=13'b0111001011010;
#1 $display("%b", po);
# 1  pi=13'b0111001011011;
#1 $display("%b", po);
# 1  pi=13'b0111001011100;
#1 $display("%b", po);
# 1  pi=13'b0111001011101;
#1 $display("%b", po);
# 1  pi=13'b0111001011110;
#1 $display("%b", po);
# 1  pi=13'b0111001011111;
#1 $display("%b", po);
# 1  pi=13'b0111001100000;
#1 $display("%b", po);
# 1  pi=13'b0111001100001;
#1 $display("%b", po);
# 1  pi=13'b0111001100010;
#1 $display("%b", po);
# 1  pi=13'b0111001100011;
#1 $display("%b", po);
# 1  pi=13'b0111001100100;
#1 $display("%b", po);
# 1  pi=13'b0111001100101;
#1 $display("%b", po);
# 1  pi=13'b0111001100110;
#1 $display("%b", po);
# 1  pi=13'b0111001100111;
#1 $display("%b", po);
# 1  pi=13'b0111001101000;
#1 $display("%b", po);
# 1  pi=13'b0111001101001;
#1 $display("%b", po);
# 1  pi=13'b0111001101010;
#1 $display("%b", po);
# 1  pi=13'b0111001101011;
#1 $display("%b", po);
# 1  pi=13'b0111001101100;
#1 $display("%b", po);
# 1  pi=13'b0111001101101;
#1 $display("%b", po);
# 1  pi=13'b0111001101110;
#1 $display("%b", po);
# 1  pi=13'b0111001101111;
#1 $display("%b", po);
# 1  pi=13'b0111001110000;
#1 $display("%b", po);
# 1  pi=13'b0111001110001;
#1 $display("%b", po);
# 1  pi=13'b0111001110010;
#1 $display("%b", po);
# 1  pi=13'b0111001110011;
#1 $display("%b", po);
# 1  pi=13'b0111001110100;
#1 $display("%b", po);
# 1  pi=13'b0111001110101;
#1 $display("%b", po);
# 1  pi=13'b0111001110110;
#1 $display("%b", po);
# 1  pi=13'b0111001110111;
#1 $display("%b", po);
# 1  pi=13'b0111001111000;
#1 $display("%b", po);
# 1  pi=13'b0111001111001;
#1 $display("%b", po);
# 1  pi=13'b0111001111010;
#1 $display("%b", po);
# 1  pi=13'b0111001111011;
#1 $display("%b", po);
# 1  pi=13'b0111001111100;
#1 $display("%b", po);
# 1  pi=13'b0111001111101;
#1 $display("%b", po);
# 1  pi=13'b0111001111110;
#1 $display("%b", po);
# 1  pi=13'b0111001111111;
#1 $display("%b", po);
# 1  pi=13'b0111010000000;
#1 $display("%b", po);
# 1  pi=13'b0111010000001;
#1 $display("%b", po);
# 1  pi=13'b0111010000010;
#1 $display("%b", po);
# 1  pi=13'b0111010000011;
#1 $display("%b", po);
# 1  pi=13'b0111010000100;
#1 $display("%b", po);
# 1  pi=13'b0111010000101;
#1 $display("%b", po);
# 1  pi=13'b0111010000110;
#1 $display("%b", po);
# 1  pi=13'b0111010000111;
#1 $display("%b", po);
# 1  pi=13'b0111010001000;
#1 $display("%b", po);
# 1  pi=13'b0111010001001;
#1 $display("%b", po);
# 1  pi=13'b0111010001010;
#1 $display("%b", po);
# 1  pi=13'b0111010001011;
#1 $display("%b", po);
# 1  pi=13'b0111010001100;
#1 $display("%b", po);
# 1  pi=13'b0111010001101;
#1 $display("%b", po);
# 1  pi=13'b0111010001110;
#1 $display("%b", po);
# 1  pi=13'b0111010001111;
#1 $display("%b", po);
# 1  pi=13'b0111010010000;
#1 $display("%b", po);
# 1  pi=13'b0111010010001;
#1 $display("%b", po);
# 1  pi=13'b0111010010010;
#1 $display("%b", po);
# 1  pi=13'b0111010010011;
#1 $display("%b", po);
# 1  pi=13'b0111010010100;
#1 $display("%b", po);
# 1  pi=13'b0111010010101;
#1 $display("%b", po);
# 1  pi=13'b0111010010110;
#1 $display("%b", po);
# 1  pi=13'b0111010010111;
#1 $display("%b", po);
# 1  pi=13'b0111010011000;
#1 $display("%b", po);
# 1  pi=13'b0111010011001;
#1 $display("%b", po);
# 1  pi=13'b0111010011010;
#1 $display("%b", po);
# 1  pi=13'b0111010011011;
#1 $display("%b", po);
# 1  pi=13'b0111010011100;
#1 $display("%b", po);
# 1  pi=13'b0111010011101;
#1 $display("%b", po);
# 1  pi=13'b0111010011110;
#1 $display("%b", po);
# 1  pi=13'b0111010011111;
#1 $display("%b", po);
# 1  pi=13'b0111010100000;
#1 $display("%b", po);
# 1  pi=13'b0111010100001;
#1 $display("%b", po);
# 1  pi=13'b0111010100010;
#1 $display("%b", po);
# 1  pi=13'b0111010100011;
#1 $display("%b", po);
# 1  pi=13'b0111010100100;
#1 $display("%b", po);
# 1  pi=13'b0111010100101;
#1 $display("%b", po);
# 1  pi=13'b0111010100110;
#1 $display("%b", po);
# 1  pi=13'b0111010100111;
#1 $display("%b", po);
# 1  pi=13'b0111010101000;
#1 $display("%b", po);
# 1  pi=13'b0111010101001;
#1 $display("%b", po);
# 1  pi=13'b0111010101010;
#1 $display("%b", po);
# 1  pi=13'b0111010101011;
#1 $display("%b", po);
# 1  pi=13'b0111010101100;
#1 $display("%b", po);
# 1  pi=13'b0111010101101;
#1 $display("%b", po);
# 1  pi=13'b0111010101110;
#1 $display("%b", po);
# 1  pi=13'b0111010101111;
#1 $display("%b", po);
# 1  pi=13'b0111010110000;
#1 $display("%b", po);
# 1  pi=13'b0111010110001;
#1 $display("%b", po);
# 1  pi=13'b0111010110010;
#1 $display("%b", po);
# 1  pi=13'b0111010110011;
#1 $display("%b", po);
# 1  pi=13'b0111010110100;
#1 $display("%b", po);
# 1  pi=13'b0111010110101;
#1 $display("%b", po);
# 1  pi=13'b0111010110110;
#1 $display("%b", po);
# 1  pi=13'b0111010110111;
#1 $display("%b", po);
# 1  pi=13'b0111010111000;
#1 $display("%b", po);
# 1  pi=13'b0111010111001;
#1 $display("%b", po);
# 1  pi=13'b0111010111010;
#1 $display("%b", po);
# 1  pi=13'b0111010111011;
#1 $display("%b", po);
# 1  pi=13'b0111010111100;
#1 $display("%b", po);
# 1  pi=13'b0111010111101;
#1 $display("%b", po);
# 1  pi=13'b0111010111110;
#1 $display("%b", po);
# 1  pi=13'b0111010111111;
#1 $display("%b", po);
# 1  pi=13'b0111011000000;
#1 $display("%b", po);
# 1  pi=13'b0111011000001;
#1 $display("%b", po);
# 1  pi=13'b0111011000010;
#1 $display("%b", po);
# 1  pi=13'b0111011000011;
#1 $display("%b", po);
# 1  pi=13'b0111011000100;
#1 $display("%b", po);
# 1  pi=13'b0111011000101;
#1 $display("%b", po);
# 1  pi=13'b0111011000110;
#1 $display("%b", po);
# 1  pi=13'b0111011000111;
#1 $display("%b", po);
# 1  pi=13'b0111011001000;
#1 $display("%b", po);
# 1  pi=13'b0111011001001;
#1 $display("%b", po);
# 1  pi=13'b0111011001010;
#1 $display("%b", po);
# 1  pi=13'b0111011001011;
#1 $display("%b", po);
# 1  pi=13'b0111011001100;
#1 $display("%b", po);
# 1  pi=13'b0111011001101;
#1 $display("%b", po);
# 1  pi=13'b0111011001110;
#1 $display("%b", po);
# 1  pi=13'b0111011001111;
#1 $display("%b", po);
# 1  pi=13'b0111011010000;
#1 $display("%b", po);
# 1  pi=13'b0111011010001;
#1 $display("%b", po);
# 1  pi=13'b0111011010010;
#1 $display("%b", po);
# 1  pi=13'b0111011010011;
#1 $display("%b", po);
# 1  pi=13'b0111011010100;
#1 $display("%b", po);
# 1  pi=13'b0111011010101;
#1 $display("%b", po);
# 1  pi=13'b0111011010110;
#1 $display("%b", po);
# 1  pi=13'b0111011010111;
#1 $display("%b", po);
# 1  pi=13'b0111011011000;
#1 $display("%b", po);
# 1  pi=13'b0111011011001;
#1 $display("%b", po);
# 1  pi=13'b0111011011010;
#1 $display("%b", po);
# 1  pi=13'b0111011011011;
#1 $display("%b", po);
# 1  pi=13'b0111011011100;
#1 $display("%b", po);
# 1  pi=13'b0111011011101;
#1 $display("%b", po);
# 1  pi=13'b0111011011110;
#1 $display("%b", po);
# 1  pi=13'b0111011011111;
#1 $display("%b", po);
# 1  pi=13'b0111011100000;
#1 $display("%b", po);
# 1  pi=13'b0111011100001;
#1 $display("%b", po);
# 1  pi=13'b0111011100010;
#1 $display("%b", po);
# 1  pi=13'b0111011100011;
#1 $display("%b", po);
# 1  pi=13'b0111011100100;
#1 $display("%b", po);
# 1  pi=13'b0111011100101;
#1 $display("%b", po);
# 1  pi=13'b0111011100110;
#1 $display("%b", po);
# 1  pi=13'b0111011100111;
#1 $display("%b", po);
# 1  pi=13'b0111011101000;
#1 $display("%b", po);
# 1  pi=13'b0111011101001;
#1 $display("%b", po);
# 1  pi=13'b0111011101010;
#1 $display("%b", po);
# 1  pi=13'b0111011101011;
#1 $display("%b", po);
# 1  pi=13'b0111011101100;
#1 $display("%b", po);
# 1  pi=13'b0111011101101;
#1 $display("%b", po);
# 1  pi=13'b0111011101110;
#1 $display("%b", po);
# 1  pi=13'b0111011101111;
#1 $display("%b", po);
# 1  pi=13'b0111011110000;
#1 $display("%b", po);
# 1  pi=13'b0111011110001;
#1 $display("%b", po);
# 1  pi=13'b0111011110010;
#1 $display("%b", po);
# 1  pi=13'b0111011110011;
#1 $display("%b", po);
# 1  pi=13'b0111011110100;
#1 $display("%b", po);
# 1  pi=13'b0111011110101;
#1 $display("%b", po);
# 1  pi=13'b0111011110110;
#1 $display("%b", po);
# 1  pi=13'b0111011110111;
#1 $display("%b", po);
# 1  pi=13'b0111011111000;
#1 $display("%b", po);
# 1  pi=13'b0111011111001;
#1 $display("%b", po);
# 1  pi=13'b0111011111010;
#1 $display("%b", po);
# 1  pi=13'b0111011111011;
#1 $display("%b", po);
# 1  pi=13'b0111011111100;
#1 $display("%b", po);
# 1  pi=13'b0111011111101;
#1 $display("%b", po);
# 1  pi=13'b0111011111110;
#1 $display("%b", po);
# 1  pi=13'b0111011111111;
#1 $display("%b", po);
# 1  pi=13'b0111100000000;
#1 $display("%b", po);
# 1  pi=13'b0111100000001;
#1 $display("%b", po);
# 1  pi=13'b0111100000010;
#1 $display("%b", po);
# 1  pi=13'b0111100000011;
#1 $display("%b", po);
# 1  pi=13'b0111100000100;
#1 $display("%b", po);
# 1  pi=13'b0111100000101;
#1 $display("%b", po);
# 1  pi=13'b0111100000110;
#1 $display("%b", po);
# 1  pi=13'b0111100000111;
#1 $display("%b", po);
# 1  pi=13'b0111100001000;
#1 $display("%b", po);
# 1  pi=13'b0111100001001;
#1 $display("%b", po);
# 1  pi=13'b0111100001010;
#1 $display("%b", po);
# 1  pi=13'b0111100001011;
#1 $display("%b", po);
# 1  pi=13'b0111100001100;
#1 $display("%b", po);
# 1  pi=13'b0111100001101;
#1 $display("%b", po);
# 1  pi=13'b0111100001110;
#1 $display("%b", po);
# 1  pi=13'b0111100001111;
#1 $display("%b", po);
# 1  pi=13'b0111100010000;
#1 $display("%b", po);
# 1  pi=13'b0111100010001;
#1 $display("%b", po);
# 1  pi=13'b0111100010010;
#1 $display("%b", po);
# 1  pi=13'b0111100010011;
#1 $display("%b", po);
# 1  pi=13'b0111100010100;
#1 $display("%b", po);
# 1  pi=13'b0111100010101;
#1 $display("%b", po);
# 1  pi=13'b0111100010110;
#1 $display("%b", po);
# 1  pi=13'b0111100010111;
#1 $display("%b", po);
# 1  pi=13'b0111100011000;
#1 $display("%b", po);
# 1  pi=13'b0111100011001;
#1 $display("%b", po);
# 1  pi=13'b0111100011010;
#1 $display("%b", po);
# 1  pi=13'b0111100011011;
#1 $display("%b", po);
# 1  pi=13'b0111100011100;
#1 $display("%b", po);
# 1  pi=13'b0111100011101;
#1 $display("%b", po);
# 1  pi=13'b0111100011110;
#1 $display("%b", po);
# 1  pi=13'b0111100011111;
#1 $display("%b", po);
# 1  pi=13'b0111100100000;
#1 $display("%b", po);
# 1  pi=13'b0111100100001;
#1 $display("%b", po);
# 1  pi=13'b0111100100010;
#1 $display("%b", po);
# 1  pi=13'b0111100100011;
#1 $display("%b", po);
# 1  pi=13'b0111100100100;
#1 $display("%b", po);
# 1  pi=13'b0111100100101;
#1 $display("%b", po);
# 1  pi=13'b0111100100110;
#1 $display("%b", po);
# 1  pi=13'b0111100100111;
#1 $display("%b", po);
# 1  pi=13'b0111100101000;
#1 $display("%b", po);
# 1  pi=13'b0111100101001;
#1 $display("%b", po);
# 1  pi=13'b0111100101010;
#1 $display("%b", po);
# 1  pi=13'b0111100101011;
#1 $display("%b", po);
# 1  pi=13'b0111100101100;
#1 $display("%b", po);
# 1  pi=13'b0111100101101;
#1 $display("%b", po);
# 1  pi=13'b0111100101110;
#1 $display("%b", po);
# 1  pi=13'b0111100101111;
#1 $display("%b", po);
# 1  pi=13'b0111100110000;
#1 $display("%b", po);
# 1  pi=13'b0111100110001;
#1 $display("%b", po);
# 1  pi=13'b0111100110010;
#1 $display("%b", po);
# 1  pi=13'b0111100110011;
#1 $display("%b", po);
# 1  pi=13'b0111100110100;
#1 $display("%b", po);
# 1  pi=13'b0111100110101;
#1 $display("%b", po);
# 1  pi=13'b0111100110110;
#1 $display("%b", po);
# 1  pi=13'b0111100110111;
#1 $display("%b", po);
# 1  pi=13'b0111100111000;
#1 $display("%b", po);
# 1  pi=13'b0111100111001;
#1 $display("%b", po);
# 1  pi=13'b0111100111010;
#1 $display("%b", po);
# 1  pi=13'b0111100111011;
#1 $display("%b", po);
# 1  pi=13'b0111100111100;
#1 $display("%b", po);
# 1  pi=13'b0111100111101;
#1 $display("%b", po);
# 1  pi=13'b0111100111110;
#1 $display("%b", po);
# 1  pi=13'b0111100111111;
#1 $display("%b", po);
# 1  pi=13'b0111101000000;
#1 $display("%b", po);
# 1  pi=13'b0111101000001;
#1 $display("%b", po);
# 1  pi=13'b0111101000010;
#1 $display("%b", po);
# 1  pi=13'b0111101000011;
#1 $display("%b", po);
# 1  pi=13'b0111101000100;
#1 $display("%b", po);
# 1  pi=13'b0111101000101;
#1 $display("%b", po);
# 1  pi=13'b0111101000110;
#1 $display("%b", po);
# 1  pi=13'b0111101000111;
#1 $display("%b", po);
# 1  pi=13'b0111101001000;
#1 $display("%b", po);
# 1  pi=13'b0111101001001;
#1 $display("%b", po);
# 1  pi=13'b0111101001010;
#1 $display("%b", po);
# 1  pi=13'b0111101001011;
#1 $display("%b", po);
# 1  pi=13'b0111101001100;
#1 $display("%b", po);
# 1  pi=13'b0111101001101;
#1 $display("%b", po);
# 1  pi=13'b0111101001110;
#1 $display("%b", po);
# 1  pi=13'b0111101001111;
#1 $display("%b", po);
# 1  pi=13'b0111101010000;
#1 $display("%b", po);
# 1  pi=13'b0111101010001;
#1 $display("%b", po);
# 1  pi=13'b0111101010010;
#1 $display("%b", po);
# 1  pi=13'b0111101010011;
#1 $display("%b", po);
# 1  pi=13'b0111101010100;
#1 $display("%b", po);
# 1  pi=13'b0111101010101;
#1 $display("%b", po);
# 1  pi=13'b0111101010110;
#1 $display("%b", po);
# 1  pi=13'b0111101010111;
#1 $display("%b", po);
# 1  pi=13'b0111101011000;
#1 $display("%b", po);
# 1  pi=13'b0111101011001;
#1 $display("%b", po);
# 1  pi=13'b0111101011010;
#1 $display("%b", po);
# 1  pi=13'b0111101011011;
#1 $display("%b", po);
# 1  pi=13'b0111101011100;
#1 $display("%b", po);
# 1  pi=13'b0111101011101;
#1 $display("%b", po);
# 1  pi=13'b0111101011110;
#1 $display("%b", po);
# 1  pi=13'b0111101011111;
#1 $display("%b", po);
# 1  pi=13'b0111101100000;
#1 $display("%b", po);
# 1  pi=13'b0111101100001;
#1 $display("%b", po);
# 1  pi=13'b0111101100010;
#1 $display("%b", po);
# 1  pi=13'b0111101100011;
#1 $display("%b", po);
# 1  pi=13'b0111101100100;
#1 $display("%b", po);
# 1  pi=13'b0111101100101;
#1 $display("%b", po);
# 1  pi=13'b0111101100110;
#1 $display("%b", po);
# 1  pi=13'b0111101100111;
#1 $display("%b", po);
# 1  pi=13'b0111101101000;
#1 $display("%b", po);
# 1  pi=13'b0111101101001;
#1 $display("%b", po);
# 1  pi=13'b0111101101010;
#1 $display("%b", po);
# 1  pi=13'b0111101101011;
#1 $display("%b", po);
# 1  pi=13'b0111101101100;
#1 $display("%b", po);
# 1  pi=13'b0111101101101;
#1 $display("%b", po);
# 1  pi=13'b0111101101110;
#1 $display("%b", po);
# 1  pi=13'b0111101101111;
#1 $display("%b", po);
# 1  pi=13'b0111101110000;
#1 $display("%b", po);
# 1  pi=13'b0111101110001;
#1 $display("%b", po);
# 1  pi=13'b0111101110010;
#1 $display("%b", po);
# 1  pi=13'b0111101110011;
#1 $display("%b", po);
# 1  pi=13'b0111101110100;
#1 $display("%b", po);
# 1  pi=13'b0111101110101;
#1 $display("%b", po);
# 1  pi=13'b0111101110110;
#1 $display("%b", po);
# 1  pi=13'b0111101110111;
#1 $display("%b", po);
# 1  pi=13'b0111101111000;
#1 $display("%b", po);
# 1  pi=13'b0111101111001;
#1 $display("%b", po);
# 1  pi=13'b0111101111010;
#1 $display("%b", po);
# 1  pi=13'b0111101111011;
#1 $display("%b", po);
# 1  pi=13'b0111101111100;
#1 $display("%b", po);
# 1  pi=13'b0111101111101;
#1 $display("%b", po);
# 1  pi=13'b0111101111110;
#1 $display("%b", po);
# 1  pi=13'b0111101111111;
#1 $display("%b", po);
# 1  pi=13'b0111110000000;
#1 $display("%b", po);
# 1  pi=13'b0111110000001;
#1 $display("%b", po);
# 1  pi=13'b0111110000010;
#1 $display("%b", po);
# 1  pi=13'b0111110000011;
#1 $display("%b", po);
# 1  pi=13'b0111110000100;
#1 $display("%b", po);
# 1  pi=13'b0111110000101;
#1 $display("%b", po);
# 1  pi=13'b0111110000110;
#1 $display("%b", po);
# 1  pi=13'b0111110000111;
#1 $display("%b", po);
# 1  pi=13'b0111110001000;
#1 $display("%b", po);
# 1  pi=13'b0111110001001;
#1 $display("%b", po);
# 1  pi=13'b0111110001010;
#1 $display("%b", po);
# 1  pi=13'b0111110001011;
#1 $display("%b", po);
# 1  pi=13'b0111110001100;
#1 $display("%b", po);
# 1  pi=13'b0111110001101;
#1 $display("%b", po);
# 1  pi=13'b0111110001110;
#1 $display("%b", po);
# 1  pi=13'b0111110001111;
#1 $display("%b", po);
# 1  pi=13'b0111110010000;
#1 $display("%b", po);
# 1  pi=13'b0111110010001;
#1 $display("%b", po);
# 1  pi=13'b0111110010010;
#1 $display("%b", po);
# 1  pi=13'b0111110010011;
#1 $display("%b", po);
# 1  pi=13'b0111110010100;
#1 $display("%b", po);
# 1  pi=13'b0111110010101;
#1 $display("%b", po);
# 1  pi=13'b0111110010110;
#1 $display("%b", po);
# 1  pi=13'b0111110010111;
#1 $display("%b", po);
# 1  pi=13'b0111110011000;
#1 $display("%b", po);
# 1  pi=13'b0111110011001;
#1 $display("%b", po);
# 1  pi=13'b0111110011010;
#1 $display("%b", po);
# 1  pi=13'b0111110011011;
#1 $display("%b", po);
# 1  pi=13'b0111110011100;
#1 $display("%b", po);
# 1  pi=13'b0111110011101;
#1 $display("%b", po);
# 1  pi=13'b0111110011110;
#1 $display("%b", po);
# 1  pi=13'b0111110011111;
#1 $display("%b", po);
# 1  pi=13'b0111110100000;
#1 $display("%b", po);
# 1  pi=13'b0111110100001;
#1 $display("%b", po);
# 1  pi=13'b0111110100010;
#1 $display("%b", po);
# 1  pi=13'b0111110100011;
#1 $display("%b", po);
# 1  pi=13'b0111110100100;
#1 $display("%b", po);
# 1  pi=13'b0111110100101;
#1 $display("%b", po);
# 1  pi=13'b0111110100110;
#1 $display("%b", po);
# 1  pi=13'b0111110100111;
#1 $display("%b", po);
# 1  pi=13'b0111110101000;
#1 $display("%b", po);
# 1  pi=13'b0111110101001;
#1 $display("%b", po);
# 1  pi=13'b0111110101010;
#1 $display("%b", po);
# 1  pi=13'b0111110101011;
#1 $display("%b", po);
# 1  pi=13'b0111110101100;
#1 $display("%b", po);
# 1  pi=13'b0111110101101;
#1 $display("%b", po);
# 1  pi=13'b0111110101110;
#1 $display("%b", po);
# 1  pi=13'b0111110101111;
#1 $display("%b", po);
# 1  pi=13'b0111110110000;
#1 $display("%b", po);
# 1  pi=13'b0111110110001;
#1 $display("%b", po);
# 1  pi=13'b0111110110010;
#1 $display("%b", po);
# 1  pi=13'b0111110110011;
#1 $display("%b", po);
# 1  pi=13'b0111110110100;
#1 $display("%b", po);
# 1  pi=13'b0111110110101;
#1 $display("%b", po);
# 1  pi=13'b0111110110110;
#1 $display("%b", po);
# 1  pi=13'b0111110110111;
#1 $display("%b", po);
# 1  pi=13'b0111110111000;
#1 $display("%b", po);
# 1  pi=13'b0111110111001;
#1 $display("%b", po);
# 1  pi=13'b0111110111010;
#1 $display("%b", po);
# 1  pi=13'b0111110111011;
#1 $display("%b", po);
# 1  pi=13'b0111110111100;
#1 $display("%b", po);
# 1  pi=13'b0111110111101;
#1 $display("%b", po);
# 1  pi=13'b0111110111110;
#1 $display("%b", po);
# 1  pi=13'b0111110111111;
#1 $display("%b", po);
# 1  pi=13'b0111111000000;
#1 $display("%b", po);
# 1  pi=13'b0111111000001;
#1 $display("%b", po);
# 1  pi=13'b0111111000010;
#1 $display("%b", po);
# 1  pi=13'b0111111000011;
#1 $display("%b", po);
# 1  pi=13'b0111111000100;
#1 $display("%b", po);
# 1  pi=13'b0111111000101;
#1 $display("%b", po);
# 1  pi=13'b0111111000110;
#1 $display("%b", po);
# 1  pi=13'b0111111000111;
#1 $display("%b", po);
# 1  pi=13'b0111111001000;
#1 $display("%b", po);
# 1  pi=13'b0111111001001;
#1 $display("%b", po);
# 1  pi=13'b0111111001010;
#1 $display("%b", po);
# 1  pi=13'b0111111001011;
#1 $display("%b", po);
# 1  pi=13'b0111111001100;
#1 $display("%b", po);
# 1  pi=13'b0111111001101;
#1 $display("%b", po);
# 1  pi=13'b0111111001110;
#1 $display("%b", po);
# 1  pi=13'b0111111001111;
#1 $display("%b", po);
# 1  pi=13'b0111111010000;
#1 $display("%b", po);
# 1  pi=13'b0111111010001;
#1 $display("%b", po);
# 1  pi=13'b0111111010010;
#1 $display("%b", po);
# 1  pi=13'b0111111010011;
#1 $display("%b", po);
# 1  pi=13'b0111111010100;
#1 $display("%b", po);
# 1  pi=13'b0111111010101;
#1 $display("%b", po);
# 1  pi=13'b0111111010110;
#1 $display("%b", po);
# 1  pi=13'b0111111010111;
#1 $display("%b", po);
# 1  pi=13'b0111111011000;
#1 $display("%b", po);
# 1  pi=13'b0111111011001;
#1 $display("%b", po);
# 1  pi=13'b0111111011010;
#1 $display("%b", po);
# 1  pi=13'b0111111011011;
#1 $display("%b", po);
# 1  pi=13'b0111111011100;
#1 $display("%b", po);
# 1  pi=13'b0111111011101;
#1 $display("%b", po);
# 1  pi=13'b0111111011110;
#1 $display("%b", po);
# 1  pi=13'b0111111011111;
#1 $display("%b", po);
# 1  pi=13'b0111111100000;
#1 $display("%b", po);
# 1  pi=13'b0111111100001;
#1 $display("%b", po);
# 1  pi=13'b0111111100010;
#1 $display("%b", po);
# 1  pi=13'b0111111100011;
#1 $display("%b", po);
# 1  pi=13'b0111111100100;
#1 $display("%b", po);
# 1  pi=13'b0111111100101;
#1 $display("%b", po);
# 1  pi=13'b0111111100110;
#1 $display("%b", po);
# 1  pi=13'b0111111100111;
#1 $display("%b", po);
# 1  pi=13'b0111111101000;
#1 $display("%b", po);
# 1  pi=13'b0111111101001;
#1 $display("%b", po);
# 1  pi=13'b0111111101010;
#1 $display("%b", po);
# 1  pi=13'b0111111101011;
#1 $display("%b", po);
# 1  pi=13'b0111111101100;
#1 $display("%b", po);
# 1  pi=13'b0111111101101;
#1 $display("%b", po);
# 1  pi=13'b0111111101110;
#1 $display("%b", po);
# 1  pi=13'b0111111101111;
#1 $display("%b", po);
# 1  pi=13'b0111111110000;
#1 $display("%b", po);
# 1  pi=13'b0111111110001;
#1 $display("%b", po);
# 1  pi=13'b0111111110010;
#1 $display("%b", po);
# 1  pi=13'b0111111110011;
#1 $display("%b", po);
# 1  pi=13'b0111111110100;
#1 $display("%b", po);
# 1  pi=13'b0111111110101;
#1 $display("%b", po);
# 1  pi=13'b0111111110110;
#1 $display("%b", po);
# 1  pi=13'b0111111110111;
#1 $display("%b", po);
# 1  pi=13'b0111111111000;
#1 $display("%b", po);
# 1  pi=13'b0111111111001;
#1 $display("%b", po);
# 1  pi=13'b0111111111010;
#1 $display("%b", po);
# 1  pi=13'b0111111111011;
#1 $display("%b", po);
# 1  pi=13'b0111111111100;
#1 $display("%b", po);
# 1  pi=13'b0111111111101;
#1 $display("%b", po);
# 1  pi=13'b0111111111110;
#1 $display("%b", po);
# 1  pi=13'b0111111111111;
#1 $display("%b", po);
# 1  pi=13'b1000000000000;
#1 $display("%b", po);
# 1  pi=13'b1000000000001;
#1 $display("%b", po);
# 1  pi=13'b1000000000010;
#1 $display("%b", po);
# 1  pi=13'b1000000000011;
#1 $display("%b", po);
# 1  pi=13'b1000000000100;
#1 $display("%b", po);
# 1  pi=13'b1000000000101;
#1 $display("%b", po);
# 1  pi=13'b1000000000110;
#1 $display("%b", po);
# 1  pi=13'b1000000000111;
#1 $display("%b", po);
# 1  pi=13'b1000000001000;
#1 $display("%b", po);
# 1  pi=13'b1000000001001;
#1 $display("%b", po);
# 1  pi=13'b1000000001010;
#1 $display("%b", po);
# 1  pi=13'b1000000001011;
#1 $display("%b", po);
# 1  pi=13'b1000000001100;
#1 $display("%b", po);
# 1  pi=13'b1000000001101;
#1 $display("%b", po);
# 1  pi=13'b1000000001110;
#1 $display("%b", po);
# 1  pi=13'b1000000001111;
#1 $display("%b", po);
# 1  pi=13'b1000000010000;
#1 $display("%b", po);
# 1  pi=13'b1000000010001;
#1 $display("%b", po);
# 1  pi=13'b1000000010010;
#1 $display("%b", po);
# 1  pi=13'b1000000010011;
#1 $display("%b", po);
# 1  pi=13'b1000000010100;
#1 $display("%b", po);
# 1  pi=13'b1000000010101;
#1 $display("%b", po);
# 1  pi=13'b1000000010110;
#1 $display("%b", po);
# 1  pi=13'b1000000010111;
#1 $display("%b", po);
# 1  pi=13'b1000000011000;
#1 $display("%b", po);
# 1  pi=13'b1000000011001;
#1 $display("%b", po);
# 1  pi=13'b1000000011010;
#1 $display("%b", po);
# 1  pi=13'b1000000011011;
#1 $display("%b", po);
# 1  pi=13'b1000000011100;
#1 $display("%b", po);
# 1  pi=13'b1000000011101;
#1 $display("%b", po);
# 1  pi=13'b1000000011110;
#1 $display("%b", po);
# 1  pi=13'b1000000011111;
#1 $display("%b", po);
# 1  pi=13'b1000000100000;
#1 $display("%b", po);
# 1  pi=13'b1000000100001;
#1 $display("%b", po);
# 1  pi=13'b1000000100010;
#1 $display("%b", po);
# 1  pi=13'b1000000100011;
#1 $display("%b", po);
# 1  pi=13'b1000000100100;
#1 $display("%b", po);
# 1  pi=13'b1000000100101;
#1 $display("%b", po);
# 1  pi=13'b1000000100110;
#1 $display("%b", po);
# 1  pi=13'b1000000100111;
#1 $display("%b", po);
# 1  pi=13'b1000000101000;
#1 $display("%b", po);
# 1  pi=13'b1000000101001;
#1 $display("%b", po);
# 1  pi=13'b1000000101010;
#1 $display("%b", po);
# 1  pi=13'b1000000101011;
#1 $display("%b", po);
# 1  pi=13'b1000000101100;
#1 $display("%b", po);
# 1  pi=13'b1000000101101;
#1 $display("%b", po);
# 1  pi=13'b1000000101110;
#1 $display("%b", po);
# 1  pi=13'b1000000101111;
#1 $display("%b", po);
# 1  pi=13'b1000000110000;
#1 $display("%b", po);
# 1  pi=13'b1000000110001;
#1 $display("%b", po);
# 1  pi=13'b1000000110010;
#1 $display("%b", po);
# 1  pi=13'b1000000110011;
#1 $display("%b", po);
# 1  pi=13'b1000000110100;
#1 $display("%b", po);
# 1  pi=13'b1000000110101;
#1 $display("%b", po);
# 1  pi=13'b1000000110110;
#1 $display("%b", po);
# 1  pi=13'b1000000110111;
#1 $display("%b", po);
# 1  pi=13'b1000000111000;
#1 $display("%b", po);
# 1  pi=13'b1000000111001;
#1 $display("%b", po);
# 1  pi=13'b1000000111010;
#1 $display("%b", po);
# 1  pi=13'b1000000111011;
#1 $display("%b", po);
# 1  pi=13'b1000000111100;
#1 $display("%b", po);
# 1  pi=13'b1000000111101;
#1 $display("%b", po);
# 1  pi=13'b1000000111110;
#1 $display("%b", po);
# 1  pi=13'b1000000111111;
#1 $display("%b", po);
# 1  pi=13'b1000001000000;
#1 $display("%b", po);
# 1  pi=13'b1000001000001;
#1 $display("%b", po);
# 1  pi=13'b1000001000010;
#1 $display("%b", po);
# 1  pi=13'b1000001000011;
#1 $display("%b", po);
# 1  pi=13'b1000001000100;
#1 $display("%b", po);
# 1  pi=13'b1000001000101;
#1 $display("%b", po);
# 1  pi=13'b1000001000110;
#1 $display("%b", po);
# 1  pi=13'b1000001000111;
#1 $display("%b", po);
# 1  pi=13'b1000001001000;
#1 $display("%b", po);
# 1  pi=13'b1000001001001;
#1 $display("%b", po);
# 1  pi=13'b1000001001010;
#1 $display("%b", po);
# 1  pi=13'b1000001001011;
#1 $display("%b", po);
# 1  pi=13'b1000001001100;
#1 $display("%b", po);
# 1  pi=13'b1000001001101;
#1 $display("%b", po);
# 1  pi=13'b1000001001110;
#1 $display("%b", po);
# 1  pi=13'b1000001001111;
#1 $display("%b", po);
# 1  pi=13'b1000001010000;
#1 $display("%b", po);
# 1  pi=13'b1000001010001;
#1 $display("%b", po);
# 1  pi=13'b1000001010010;
#1 $display("%b", po);
# 1  pi=13'b1000001010011;
#1 $display("%b", po);
# 1  pi=13'b1000001010100;
#1 $display("%b", po);
# 1  pi=13'b1000001010101;
#1 $display("%b", po);
# 1  pi=13'b1000001010110;
#1 $display("%b", po);
# 1  pi=13'b1000001010111;
#1 $display("%b", po);
# 1  pi=13'b1000001011000;
#1 $display("%b", po);
# 1  pi=13'b1000001011001;
#1 $display("%b", po);
# 1  pi=13'b1000001011010;
#1 $display("%b", po);
# 1  pi=13'b1000001011011;
#1 $display("%b", po);
# 1  pi=13'b1000001011100;
#1 $display("%b", po);
# 1  pi=13'b1000001011101;
#1 $display("%b", po);
# 1  pi=13'b1000001011110;
#1 $display("%b", po);
# 1  pi=13'b1000001011111;
#1 $display("%b", po);
# 1  pi=13'b1000001100000;
#1 $display("%b", po);
# 1  pi=13'b1000001100001;
#1 $display("%b", po);
# 1  pi=13'b1000001100010;
#1 $display("%b", po);
# 1  pi=13'b1000001100011;
#1 $display("%b", po);
# 1  pi=13'b1000001100100;
#1 $display("%b", po);
# 1  pi=13'b1000001100101;
#1 $display("%b", po);
# 1  pi=13'b1000001100110;
#1 $display("%b", po);
# 1  pi=13'b1000001100111;
#1 $display("%b", po);
# 1  pi=13'b1000001101000;
#1 $display("%b", po);
# 1  pi=13'b1000001101001;
#1 $display("%b", po);
# 1  pi=13'b1000001101010;
#1 $display("%b", po);
# 1  pi=13'b1000001101011;
#1 $display("%b", po);
# 1  pi=13'b1000001101100;
#1 $display("%b", po);
# 1  pi=13'b1000001101101;
#1 $display("%b", po);
# 1  pi=13'b1000001101110;
#1 $display("%b", po);
# 1  pi=13'b1000001101111;
#1 $display("%b", po);
# 1  pi=13'b1000001110000;
#1 $display("%b", po);
# 1  pi=13'b1000001110001;
#1 $display("%b", po);
# 1  pi=13'b1000001110010;
#1 $display("%b", po);
# 1  pi=13'b1000001110011;
#1 $display("%b", po);
# 1  pi=13'b1000001110100;
#1 $display("%b", po);
# 1  pi=13'b1000001110101;
#1 $display("%b", po);
# 1  pi=13'b1000001110110;
#1 $display("%b", po);
# 1  pi=13'b1000001110111;
#1 $display("%b", po);
# 1  pi=13'b1000001111000;
#1 $display("%b", po);
# 1  pi=13'b1000001111001;
#1 $display("%b", po);
# 1  pi=13'b1000001111010;
#1 $display("%b", po);
# 1  pi=13'b1000001111011;
#1 $display("%b", po);
# 1  pi=13'b1000001111100;
#1 $display("%b", po);
# 1  pi=13'b1000001111101;
#1 $display("%b", po);
# 1  pi=13'b1000001111110;
#1 $display("%b", po);
# 1  pi=13'b1000001111111;
#1 $display("%b", po);
# 1  pi=13'b1000010000000;
#1 $display("%b", po);
# 1  pi=13'b1000010000001;
#1 $display("%b", po);
# 1  pi=13'b1000010000010;
#1 $display("%b", po);
# 1  pi=13'b1000010000011;
#1 $display("%b", po);
# 1  pi=13'b1000010000100;
#1 $display("%b", po);
# 1  pi=13'b1000010000101;
#1 $display("%b", po);
# 1  pi=13'b1000010000110;
#1 $display("%b", po);
# 1  pi=13'b1000010000111;
#1 $display("%b", po);
# 1  pi=13'b1000010001000;
#1 $display("%b", po);
# 1  pi=13'b1000010001001;
#1 $display("%b", po);
# 1  pi=13'b1000010001010;
#1 $display("%b", po);
# 1  pi=13'b1000010001011;
#1 $display("%b", po);
# 1  pi=13'b1000010001100;
#1 $display("%b", po);
# 1  pi=13'b1000010001101;
#1 $display("%b", po);
# 1  pi=13'b1000010001110;
#1 $display("%b", po);
# 1  pi=13'b1000010001111;
#1 $display("%b", po);
# 1  pi=13'b1000010010000;
#1 $display("%b", po);
# 1  pi=13'b1000010010001;
#1 $display("%b", po);
# 1  pi=13'b1000010010010;
#1 $display("%b", po);
# 1  pi=13'b1000010010011;
#1 $display("%b", po);
# 1  pi=13'b1000010010100;
#1 $display("%b", po);
# 1  pi=13'b1000010010101;
#1 $display("%b", po);
# 1  pi=13'b1000010010110;
#1 $display("%b", po);
# 1  pi=13'b1000010010111;
#1 $display("%b", po);
# 1  pi=13'b1000010011000;
#1 $display("%b", po);
# 1  pi=13'b1000010011001;
#1 $display("%b", po);
# 1  pi=13'b1000010011010;
#1 $display("%b", po);
# 1  pi=13'b1000010011011;
#1 $display("%b", po);
# 1  pi=13'b1000010011100;
#1 $display("%b", po);
# 1  pi=13'b1000010011101;
#1 $display("%b", po);
# 1  pi=13'b1000010011110;
#1 $display("%b", po);
# 1  pi=13'b1000010011111;
#1 $display("%b", po);
# 1  pi=13'b1000010100000;
#1 $display("%b", po);
# 1  pi=13'b1000010100001;
#1 $display("%b", po);
# 1  pi=13'b1000010100010;
#1 $display("%b", po);
# 1  pi=13'b1000010100011;
#1 $display("%b", po);
# 1  pi=13'b1000010100100;
#1 $display("%b", po);
# 1  pi=13'b1000010100101;
#1 $display("%b", po);
# 1  pi=13'b1000010100110;
#1 $display("%b", po);
# 1  pi=13'b1000010100111;
#1 $display("%b", po);
# 1  pi=13'b1000010101000;
#1 $display("%b", po);
# 1  pi=13'b1000010101001;
#1 $display("%b", po);
# 1  pi=13'b1000010101010;
#1 $display("%b", po);
# 1  pi=13'b1000010101011;
#1 $display("%b", po);
# 1  pi=13'b1000010101100;
#1 $display("%b", po);
# 1  pi=13'b1000010101101;
#1 $display("%b", po);
# 1  pi=13'b1000010101110;
#1 $display("%b", po);
# 1  pi=13'b1000010101111;
#1 $display("%b", po);
# 1  pi=13'b1000010110000;
#1 $display("%b", po);
# 1  pi=13'b1000010110001;
#1 $display("%b", po);
# 1  pi=13'b1000010110010;
#1 $display("%b", po);
# 1  pi=13'b1000010110011;
#1 $display("%b", po);
# 1  pi=13'b1000010110100;
#1 $display("%b", po);
# 1  pi=13'b1000010110101;
#1 $display("%b", po);
# 1  pi=13'b1000010110110;
#1 $display("%b", po);
# 1  pi=13'b1000010110111;
#1 $display("%b", po);
# 1  pi=13'b1000010111000;
#1 $display("%b", po);
# 1  pi=13'b1000010111001;
#1 $display("%b", po);
# 1  pi=13'b1000010111010;
#1 $display("%b", po);
# 1  pi=13'b1000010111011;
#1 $display("%b", po);
# 1  pi=13'b1000010111100;
#1 $display("%b", po);
# 1  pi=13'b1000010111101;
#1 $display("%b", po);
# 1  pi=13'b1000010111110;
#1 $display("%b", po);
# 1  pi=13'b1000010111111;
#1 $display("%b", po);
# 1  pi=13'b1000011000000;
#1 $display("%b", po);
# 1  pi=13'b1000011000001;
#1 $display("%b", po);
# 1  pi=13'b1000011000010;
#1 $display("%b", po);
# 1  pi=13'b1000011000011;
#1 $display("%b", po);
# 1  pi=13'b1000011000100;
#1 $display("%b", po);
# 1  pi=13'b1000011000101;
#1 $display("%b", po);
# 1  pi=13'b1000011000110;
#1 $display("%b", po);
# 1  pi=13'b1000011000111;
#1 $display("%b", po);
# 1  pi=13'b1000011001000;
#1 $display("%b", po);
# 1  pi=13'b1000011001001;
#1 $display("%b", po);
# 1  pi=13'b1000011001010;
#1 $display("%b", po);
# 1  pi=13'b1000011001011;
#1 $display("%b", po);
# 1  pi=13'b1000011001100;
#1 $display("%b", po);
# 1  pi=13'b1000011001101;
#1 $display("%b", po);
# 1  pi=13'b1000011001110;
#1 $display("%b", po);
# 1  pi=13'b1000011001111;
#1 $display("%b", po);
# 1  pi=13'b1000011010000;
#1 $display("%b", po);
# 1  pi=13'b1000011010001;
#1 $display("%b", po);
# 1  pi=13'b1000011010010;
#1 $display("%b", po);
# 1  pi=13'b1000011010011;
#1 $display("%b", po);
# 1  pi=13'b1000011010100;
#1 $display("%b", po);
# 1  pi=13'b1000011010101;
#1 $display("%b", po);
# 1  pi=13'b1000011010110;
#1 $display("%b", po);
# 1  pi=13'b1000011010111;
#1 $display("%b", po);
# 1  pi=13'b1000011011000;
#1 $display("%b", po);
# 1  pi=13'b1000011011001;
#1 $display("%b", po);
# 1  pi=13'b1000011011010;
#1 $display("%b", po);
# 1  pi=13'b1000011011011;
#1 $display("%b", po);
# 1  pi=13'b1000011011100;
#1 $display("%b", po);
# 1  pi=13'b1000011011101;
#1 $display("%b", po);
# 1  pi=13'b1000011011110;
#1 $display("%b", po);
# 1  pi=13'b1000011011111;
#1 $display("%b", po);
# 1  pi=13'b1000011100000;
#1 $display("%b", po);
# 1  pi=13'b1000011100001;
#1 $display("%b", po);
# 1  pi=13'b1000011100010;
#1 $display("%b", po);
# 1  pi=13'b1000011100011;
#1 $display("%b", po);
# 1  pi=13'b1000011100100;
#1 $display("%b", po);
# 1  pi=13'b1000011100101;
#1 $display("%b", po);
# 1  pi=13'b1000011100110;
#1 $display("%b", po);
# 1  pi=13'b1000011100111;
#1 $display("%b", po);
# 1  pi=13'b1000011101000;
#1 $display("%b", po);
# 1  pi=13'b1000011101001;
#1 $display("%b", po);
# 1  pi=13'b1000011101010;
#1 $display("%b", po);
# 1  pi=13'b1000011101011;
#1 $display("%b", po);
# 1  pi=13'b1000011101100;
#1 $display("%b", po);
# 1  pi=13'b1000011101101;
#1 $display("%b", po);
# 1  pi=13'b1000011101110;
#1 $display("%b", po);
# 1  pi=13'b1000011101111;
#1 $display("%b", po);
# 1  pi=13'b1000011110000;
#1 $display("%b", po);
# 1  pi=13'b1000011110001;
#1 $display("%b", po);
# 1  pi=13'b1000011110010;
#1 $display("%b", po);
# 1  pi=13'b1000011110011;
#1 $display("%b", po);
# 1  pi=13'b1000011110100;
#1 $display("%b", po);
# 1  pi=13'b1000011110101;
#1 $display("%b", po);
# 1  pi=13'b1000011110110;
#1 $display("%b", po);
# 1  pi=13'b1000011110111;
#1 $display("%b", po);
# 1  pi=13'b1000011111000;
#1 $display("%b", po);
# 1  pi=13'b1000011111001;
#1 $display("%b", po);
# 1  pi=13'b1000011111010;
#1 $display("%b", po);
# 1  pi=13'b1000011111011;
#1 $display("%b", po);
# 1  pi=13'b1000011111100;
#1 $display("%b", po);
# 1  pi=13'b1000011111101;
#1 $display("%b", po);
# 1  pi=13'b1000011111110;
#1 $display("%b", po);
# 1  pi=13'b1000011111111;
#1 $display("%b", po);
# 1  pi=13'b1000100000000;
#1 $display("%b", po);
# 1  pi=13'b1000100000001;
#1 $display("%b", po);
# 1  pi=13'b1000100000010;
#1 $display("%b", po);
# 1  pi=13'b1000100000011;
#1 $display("%b", po);
# 1  pi=13'b1000100000100;
#1 $display("%b", po);
# 1  pi=13'b1000100000101;
#1 $display("%b", po);
# 1  pi=13'b1000100000110;
#1 $display("%b", po);
# 1  pi=13'b1000100000111;
#1 $display("%b", po);
# 1  pi=13'b1000100001000;
#1 $display("%b", po);
# 1  pi=13'b1000100001001;
#1 $display("%b", po);
# 1  pi=13'b1000100001010;
#1 $display("%b", po);
# 1  pi=13'b1000100001011;
#1 $display("%b", po);
# 1  pi=13'b1000100001100;
#1 $display("%b", po);
# 1  pi=13'b1000100001101;
#1 $display("%b", po);
# 1  pi=13'b1000100001110;
#1 $display("%b", po);
# 1  pi=13'b1000100001111;
#1 $display("%b", po);
# 1  pi=13'b1000100010000;
#1 $display("%b", po);
# 1  pi=13'b1000100010001;
#1 $display("%b", po);
# 1  pi=13'b1000100010010;
#1 $display("%b", po);
# 1  pi=13'b1000100010011;
#1 $display("%b", po);
# 1  pi=13'b1000100010100;
#1 $display("%b", po);
# 1  pi=13'b1000100010101;
#1 $display("%b", po);
# 1  pi=13'b1000100010110;
#1 $display("%b", po);
# 1  pi=13'b1000100010111;
#1 $display("%b", po);
# 1  pi=13'b1000100011000;
#1 $display("%b", po);
# 1  pi=13'b1000100011001;
#1 $display("%b", po);
# 1  pi=13'b1000100011010;
#1 $display("%b", po);
# 1  pi=13'b1000100011011;
#1 $display("%b", po);
# 1  pi=13'b1000100011100;
#1 $display("%b", po);
# 1  pi=13'b1000100011101;
#1 $display("%b", po);
# 1  pi=13'b1000100011110;
#1 $display("%b", po);
# 1  pi=13'b1000100011111;
#1 $display("%b", po);
# 1  pi=13'b1000100100000;
#1 $display("%b", po);
# 1  pi=13'b1000100100001;
#1 $display("%b", po);
# 1  pi=13'b1000100100010;
#1 $display("%b", po);
# 1  pi=13'b1000100100011;
#1 $display("%b", po);
# 1  pi=13'b1000100100100;
#1 $display("%b", po);
# 1  pi=13'b1000100100101;
#1 $display("%b", po);
# 1  pi=13'b1000100100110;
#1 $display("%b", po);
# 1  pi=13'b1000100100111;
#1 $display("%b", po);
# 1  pi=13'b1000100101000;
#1 $display("%b", po);
# 1  pi=13'b1000100101001;
#1 $display("%b", po);
# 1  pi=13'b1000100101010;
#1 $display("%b", po);
# 1  pi=13'b1000100101011;
#1 $display("%b", po);
# 1  pi=13'b1000100101100;
#1 $display("%b", po);
# 1  pi=13'b1000100101101;
#1 $display("%b", po);
# 1  pi=13'b1000100101110;
#1 $display("%b", po);
# 1  pi=13'b1000100101111;
#1 $display("%b", po);
# 1  pi=13'b1000100110000;
#1 $display("%b", po);
# 1  pi=13'b1000100110001;
#1 $display("%b", po);
# 1  pi=13'b1000100110010;
#1 $display("%b", po);
# 1  pi=13'b1000100110011;
#1 $display("%b", po);
# 1  pi=13'b1000100110100;
#1 $display("%b", po);
# 1  pi=13'b1000100110101;
#1 $display("%b", po);
# 1  pi=13'b1000100110110;
#1 $display("%b", po);
# 1  pi=13'b1000100110111;
#1 $display("%b", po);
# 1  pi=13'b1000100111000;
#1 $display("%b", po);
# 1  pi=13'b1000100111001;
#1 $display("%b", po);
# 1  pi=13'b1000100111010;
#1 $display("%b", po);
# 1  pi=13'b1000100111011;
#1 $display("%b", po);
# 1  pi=13'b1000100111100;
#1 $display("%b", po);
# 1  pi=13'b1000100111101;
#1 $display("%b", po);
# 1  pi=13'b1000100111110;
#1 $display("%b", po);
# 1  pi=13'b1000100111111;
#1 $display("%b", po);
# 1  pi=13'b1000101000000;
#1 $display("%b", po);
# 1  pi=13'b1000101000001;
#1 $display("%b", po);
# 1  pi=13'b1000101000010;
#1 $display("%b", po);
# 1  pi=13'b1000101000011;
#1 $display("%b", po);
# 1  pi=13'b1000101000100;
#1 $display("%b", po);
# 1  pi=13'b1000101000101;
#1 $display("%b", po);
# 1  pi=13'b1000101000110;
#1 $display("%b", po);
# 1  pi=13'b1000101000111;
#1 $display("%b", po);
# 1  pi=13'b1000101001000;
#1 $display("%b", po);
# 1  pi=13'b1000101001001;
#1 $display("%b", po);
# 1  pi=13'b1000101001010;
#1 $display("%b", po);
# 1  pi=13'b1000101001011;
#1 $display("%b", po);
# 1  pi=13'b1000101001100;
#1 $display("%b", po);
# 1  pi=13'b1000101001101;
#1 $display("%b", po);
# 1  pi=13'b1000101001110;
#1 $display("%b", po);
# 1  pi=13'b1000101001111;
#1 $display("%b", po);
# 1  pi=13'b1000101010000;
#1 $display("%b", po);
# 1  pi=13'b1000101010001;
#1 $display("%b", po);
# 1  pi=13'b1000101010010;
#1 $display("%b", po);
# 1  pi=13'b1000101010011;
#1 $display("%b", po);
# 1  pi=13'b1000101010100;
#1 $display("%b", po);
# 1  pi=13'b1000101010101;
#1 $display("%b", po);
# 1  pi=13'b1000101010110;
#1 $display("%b", po);
# 1  pi=13'b1000101010111;
#1 $display("%b", po);
# 1  pi=13'b1000101011000;
#1 $display("%b", po);
# 1  pi=13'b1000101011001;
#1 $display("%b", po);
# 1  pi=13'b1000101011010;
#1 $display("%b", po);
# 1  pi=13'b1000101011011;
#1 $display("%b", po);
# 1  pi=13'b1000101011100;
#1 $display("%b", po);
# 1  pi=13'b1000101011101;
#1 $display("%b", po);
# 1  pi=13'b1000101011110;
#1 $display("%b", po);
# 1  pi=13'b1000101011111;
#1 $display("%b", po);
# 1  pi=13'b1000101100000;
#1 $display("%b", po);
# 1  pi=13'b1000101100001;
#1 $display("%b", po);
# 1  pi=13'b1000101100010;
#1 $display("%b", po);
# 1  pi=13'b1000101100011;
#1 $display("%b", po);
# 1  pi=13'b1000101100100;
#1 $display("%b", po);
# 1  pi=13'b1000101100101;
#1 $display("%b", po);
# 1  pi=13'b1000101100110;
#1 $display("%b", po);
# 1  pi=13'b1000101100111;
#1 $display("%b", po);
# 1  pi=13'b1000101101000;
#1 $display("%b", po);
# 1  pi=13'b1000101101001;
#1 $display("%b", po);
# 1  pi=13'b1000101101010;
#1 $display("%b", po);
# 1  pi=13'b1000101101011;
#1 $display("%b", po);
# 1  pi=13'b1000101101100;
#1 $display("%b", po);
# 1  pi=13'b1000101101101;
#1 $display("%b", po);
# 1  pi=13'b1000101101110;
#1 $display("%b", po);
# 1  pi=13'b1000101101111;
#1 $display("%b", po);
# 1  pi=13'b1000101110000;
#1 $display("%b", po);
# 1  pi=13'b1000101110001;
#1 $display("%b", po);
# 1  pi=13'b1000101110010;
#1 $display("%b", po);
# 1  pi=13'b1000101110011;
#1 $display("%b", po);
# 1  pi=13'b1000101110100;
#1 $display("%b", po);
# 1  pi=13'b1000101110101;
#1 $display("%b", po);
# 1  pi=13'b1000101110110;
#1 $display("%b", po);
# 1  pi=13'b1000101110111;
#1 $display("%b", po);
# 1  pi=13'b1000101111000;
#1 $display("%b", po);
# 1  pi=13'b1000101111001;
#1 $display("%b", po);
# 1  pi=13'b1000101111010;
#1 $display("%b", po);
# 1  pi=13'b1000101111011;
#1 $display("%b", po);
# 1  pi=13'b1000101111100;
#1 $display("%b", po);
# 1  pi=13'b1000101111101;
#1 $display("%b", po);
# 1  pi=13'b1000101111110;
#1 $display("%b", po);
# 1  pi=13'b1000101111111;
#1 $display("%b", po);
# 1  pi=13'b1000110000000;
#1 $display("%b", po);
# 1  pi=13'b1000110000001;
#1 $display("%b", po);
# 1  pi=13'b1000110000010;
#1 $display("%b", po);
# 1  pi=13'b1000110000011;
#1 $display("%b", po);
# 1  pi=13'b1000110000100;
#1 $display("%b", po);
# 1  pi=13'b1000110000101;
#1 $display("%b", po);
# 1  pi=13'b1000110000110;
#1 $display("%b", po);
# 1  pi=13'b1000110000111;
#1 $display("%b", po);
# 1  pi=13'b1000110001000;
#1 $display("%b", po);
# 1  pi=13'b1000110001001;
#1 $display("%b", po);
# 1  pi=13'b1000110001010;
#1 $display("%b", po);
# 1  pi=13'b1000110001011;
#1 $display("%b", po);
# 1  pi=13'b1000110001100;
#1 $display("%b", po);
# 1  pi=13'b1000110001101;
#1 $display("%b", po);
# 1  pi=13'b1000110001110;
#1 $display("%b", po);
# 1  pi=13'b1000110001111;
#1 $display("%b", po);
# 1  pi=13'b1000110010000;
#1 $display("%b", po);
# 1  pi=13'b1000110010001;
#1 $display("%b", po);
# 1  pi=13'b1000110010010;
#1 $display("%b", po);
# 1  pi=13'b1000110010011;
#1 $display("%b", po);
# 1  pi=13'b1000110010100;
#1 $display("%b", po);
# 1  pi=13'b1000110010101;
#1 $display("%b", po);
# 1  pi=13'b1000110010110;
#1 $display("%b", po);
# 1  pi=13'b1000110010111;
#1 $display("%b", po);
# 1  pi=13'b1000110011000;
#1 $display("%b", po);
# 1  pi=13'b1000110011001;
#1 $display("%b", po);
# 1  pi=13'b1000110011010;
#1 $display("%b", po);
# 1  pi=13'b1000110011011;
#1 $display("%b", po);
# 1  pi=13'b1000110011100;
#1 $display("%b", po);
# 1  pi=13'b1000110011101;
#1 $display("%b", po);
# 1  pi=13'b1000110011110;
#1 $display("%b", po);
# 1  pi=13'b1000110011111;
#1 $display("%b", po);
# 1  pi=13'b1000110100000;
#1 $display("%b", po);
# 1  pi=13'b1000110100001;
#1 $display("%b", po);
# 1  pi=13'b1000110100010;
#1 $display("%b", po);
# 1  pi=13'b1000110100011;
#1 $display("%b", po);
# 1  pi=13'b1000110100100;
#1 $display("%b", po);
# 1  pi=13'b1000110100101;
#1 $display("%b", po);
# 1  pi=13'b1000110100110;
#1 $display("%b", po);
# 1  pi=13'b1000110100111;
#1 $display("%b", po);
# 1  pi=13'b1000110101000;
#1 $display("%b", po);
# 1  pi=13'b1000110101001;
#1 $display("%b", po);
# 1  pi=13'b1000110101010;
#1 $display("%b", po);
# 1  pi=13'b1000110101011;
#1 $display("%b", po);
# 1  pi=13'b1000110101100;
#1 $display("%b", po);
# 1  pi=13'b1000110101101;
#1 $display("%b", po);
# 1  pi=13'b1000110101110;
#1 $display("%b", po);
# 1  pi=13'b1000110101111;
#1 $display("%b", po);
# 1  pi=13'b1000110110000;
#1 $display("%b", po);
# 1  pi=13'b1000110110001;
#1 $display("%b", po);
# 1  pi=13'b1000110110010;
#1 $display("%b", po);
# 1  pi=13'b1000110110011;
#1 $display("%b", po);
# 1  pi=13'b1000110110100;
#1 $display("%b", po);
# 1  pi=13'b1000110110101;
#1 $display("%b", po);
# 1  pi=13'b1000110110110;
#1 $display("%b", po);
# 1  pi=13'b1000110110111;
#1 $display("%b", po);
# 1  pi=13'b1000110111000;
#1 $display("%b", po);
# 1  pi=13'b1000110111001;
#1 $display("%b", po);
# 1  pi=13'b1000110111010;
#1 $display("%b", po);
# 1  pi=13'b1000110111011;
#1 $display("%b", po);
# 1  pi=13'b1000110111100;
#1 $display("%b", po);
# 1  pi=13'b1000110111101;
#1 $display("%b", po);
# 1  pi=13'b1000110111110;
#1 $display("%b", po);
# 1  pi=13'b1000110111111;
#1 $display("%b", po);
# 1  pi=13'b1000111000000;
#1 $display("%b", po);
# 1  pi=13'b1000111000001;
#1 $display("%b", po);
# 1  pi=13'b1000111000010;
#1 $display("%b", po);
# 1  pi=13'b1000111000011;
#1 $display("%b", po);
# 1  pi=13'b1000111000100;
#1 $display("%b", po);
# 1  pi=13'b1000111000101;
#1 $display("%b", po);
# 1  pi=13'b1000111000110;
#1 $display("%b", po);
# 1  pi=13'b1000111000111;
#1 $display("%b", po);
# 1  pi=13'b1000111001000;
#1 $display("%b", po);
# 1  pi=13'b1000111001001;
#1 $display("%b", po);
# 1  pi=13'b1000111001010;
#1 $display("%b", po);
# 1  pi=13'b1000111001011;
#1 $display("%b", po);
# 1  pi=13'b1000111001100;
#1 $display("%b", po);
# 1  pi=13'b1000111001101;
#1 $display("%b", po);
# 1  pi=13'b1000111001110;
#1 $display("%b", po);
# 1  pi=13'b1000111001111;
#1 $display("%b", po);
# 1  pi=13'b1000111010000;
#1 $display("%b", po);
# 1  pi=13'b1000111010001;
#1 $display("%b", po);
# 1  pi=13'b1000111010010;
#1 $display("%b", po);
# 1  pi=13'b1000111010011;
#1 $display("%b", po);
# 1  pi=13'b1000111010100;
#1 $display("%b", po);
# 1  pi=13'b1000111010101;
#1 $display("%b", po);
# 1  pi=13'b1000111010110;
#1 $display("%b", po);
# 1  pi=13'b1000111010111;
#1 $display("%b", po);
# 1  pi=13'b1000111011000;
#1 $display("%b", po);
# 1  pi=13'b1000111011001;
#1 $display("%b", po);
# 1  pi=13'b1000111011010;
#1 $display("%b", po);
# 1  pi=13'b1000111011011;
#1 $display("%b", po);
# 1  pi=13'b1000111011100;
#1 $display("%b", po);
# 1  pi=13'b1000111011101;
#1 $display("%b", po);
# 1  pi=13'b1000111011110;
#1 $display("%b", po);
# 1  pi=13'b1000111011111;
#1 $display("%b", po);
# 1  pi=13'b1000111100000;
#1 $display("%b", po);
# 1  pi=13'b1000111100001;
#1 $display("%b", po);
# 1  pi=13'b1000111100010;
#1 $display("%b", po);
# 1  pi=13'b1000111100011;
#1 $display("%b", po);
# 1  pi=13'b1000111100100;
#1 $display("%b", po);
# 1  pi=13'b1000111100101;
#1 $display("%b", po);
# 1  pi=13'b1000111100110;
#1 $display("%b", po);
# 1  pi=13'b1000111100111;
#1 $display("%b", po);
# 1  pi=13'b1000111101000;
#1 $display("%b", po);
# 1  pi=13'b1000111101001;
#1 $display("%b", po);
# 1  pi=13'b1000111101010;
#1 $display("%b", po);
# 1  pi=13'b1000111101011;
#1 $display("%b", po);
# 1  pi=13'b1000111101100;
#1 $display("%b", po);
# 1  pi=13'b1000111101101;
#1 $display("%b", po);
# 1  pi=13'b1000111101110;
#1 $display("%b", po);
# 1  pi=13'b1000111101111;
#1 $display("%b", po);
# 1  pi=13'b1000111110000;
#1 $display("%b", po);
# 1  pi=13'b1000111110001;
#1 $display("%b", po);
# 1  pi=13'b1000111110010;
#1 $display("%b", po);
# 1  pi=13'b1000111110011;
#1 $display("%b", po);
# 1  pi=13'b1000111110100;
#1 $display("%b", po);
# 1  pi=13'b1000111110101;
#1 $display("%b", po);
# 1  pi=13'b1000111110110;
#1 $display("%b", po);
# 1  pi=13'b1000111110111;
#1 $display("%b", po);
# 1  pi=13'b1000111111000;
#1 $display("%b", po);
# 1  pi=13'b1000111111001;
#1 $display("%b", po);
# 1  pi=13'b1000111111010;
#1 $display("%b", po);
# 1  pi=13'b1000111111011;
#1 $display("%b", po);
# 1  pi=13'b1000111111100;
#1 $display("%b", po);
# 1  pi=13'b1000111111101;
#1 $display("%b", po);
# 1  pi=13'b1000111111110;
#1 $display("%b", po);
# 1  pi=13'b1000111111111;
#1 $display("%b", po);
# 1  pi=13'b1001000000000;
#1 $display("%b", po);
# 1  pi=13'b1001000000001;
#1 $display("%b", po);
# 1  pi=13'b1001000000010;
#1 $display("%b", po);
# 1  pi=13'b1001000000011;
#1 $display("%b", po);
# 1  pi=13'b1001000000100;
#1 $display("%b", po);
# 1  pi=13'b1001000000101;
#1 $display("%b", po);
# 1  pi=13'b1001000000110;
#1 $display("%b", po);
# 1  pi=13'b1001000000111;
#1 $display("%b", po);
# 1  pi=13'b1001000001000;
#1 $display("%b", po);
# 1  pi=13'b1001000001001;
#1 $display("%b", po);
# 1  pi=13'b1001000001010;
#1 $display("%b", po);
# 1  pi=13'b1001000001011;
#1 $display("%b", po);
# 1  pi=13'b1001000001100;
#1 $display("%b", po);
# 1  pi=13'b1001000001101;
#1 $display("%b", po);
# 1  pi=13'b1001000001110;
#1 $display("%b", po);
# 1  pi=13'b1001000001111;
#1 $display("%b", po);
# 1  pi=13'b1001000010000;
#1 $display("%b", po);
# 1  pi=13'b1001000010001;
#1 $display("%b", po);
# 1  pi=13'b1001000010010;
#1 $display("%b", po);
# 1  pi=13'b1001000010011;
#1 $display("%b", po);
# 1  pi=13'b1001000010100;
#1 $display("%b", po);
# 1  pi=13'b1001000010101;
#1 $display("%b", po);
# 1  pi=13'b1001000010110;
#1 $display("%b", po);
# 1  pi=13'b1001000010111;
#1 $display("%b", po);
# 1  pi=13'b1001000011000;
#1 $display("%b", po);
# 1  pi=13'b1001000011001;
#1 $display("%b", po);
# 1  pi=13'b1001000011010;
#1 $display("%b", po);
# 1  pi=13'b1001000011011;
#1 $display("%b", po);
# 1  pi=13'b1001000011100;
#1 $display("%b", po);
# 1  pi=13'b1001000011101;
#1 $display("%b", po);
# 1  pi=13'b1001000011110;
#1 $display("%b", po);
# 1  pi=13'b1001000011111;
#1 $display("%b", po);
# 1  pi=13'b1001000100000;
#1 $display("%b", po);
# 1  pi=13'b1001000100001;
#1 $display("%b", po);
# 1  pi=13'b1001000100010;
#1 $display("%b", po);
# 1  pi=13'b1001000100011;
#1 $display("%b", po);
# 1  pi=13'b1001000100100;
#1 $display("%b", po);
# 1  pi=13'b1001000100101;
#1 $display("%b", po);
# 1  pi=13'b1001000100110;
#1 $display("%b", po);
# 1  pi=13'b1001000100111;
#1 $display("%b", po);
# 1  pi=13'b1001000101000;
#1 $display("%b", po);
# 1  pi=13'b1001000101001;
#1 $display("%b", po);
# 1  pi=13'b1001000101010;
#1 $display("%b", po);
# 1  pi=13'b1001000101011;
#1 $display("%b", po);
# 1  pi=13'b1001000101100;
#1 $display("%b", po);
# 1  pi=13'b1001000101101;
#1 $display("%b", po);
# 1  pi=13'b1001000101110;
#1 $display("%b", po);
# 1  pi=13'b1001000101111;
#1 $display("%b", po);
# 1  pi=13'b1001000110000;
#1 $display("%b", po);
# 1  pi=13'b1001000110001;
#1 $display("%b", po);
# 1  pi=13'b1001000110010;
#1 $display("%b", po);
# 1  pi=13'b1001000110011;
#1 $display("%b", po);
# 1  pi=13'b1001000110100;
#1 $display("%b", po);
# 1  pi=13'b1001000110101;
#1 $display("%b", po);
# 1  pi=13'b1001000110110;
#1 $display("%b", po);
# 1  pi=13'b1001000110111;
#1 $display("%b", po);
# 1  pi=13'b1001000111000;
#1 $display("%b", po);
# 1  pi=13'b1001000111001;
#1 $display("%b", po);
# 1  pi=13'b1001000111010;
#1 $display("%b", po);
# 1  pi=13'b1001000111011;
#1 $display("%b", po);
# 1  pi=13'b1001000111100;
#1 $display("%b", po);
# 1  pi=13'b1001000111101;
#1 $display("%b", po);
# 1  pi=13'b1001000111110;
#1 $display("%b", po);
# 1  pi=13'b1001000111111;
#1 $display("%b", po);
# 1  pi=13'b1001001000000;
#1 $display("%b", po);
# 1  pi=13'b1001001000001;
#1 $display("%b", po);
# 1  pi=13'b1001001000010;
#1 $display("%b", po);
# 1  pi=13'b1001001000011;
#1 $display("%b", po);
# 1  pi=13'b1001001000100;
#1 $display("%b", po);
# 1  pi=13'b1001001000101;
#1 $display("%b", po);
# 1  pi=13'b1001001000110;
#1 $display("%b", po);
# 1  pi=13'b1001001000111;
#1 $display("%b", po);
# 1  pi=13'b1001001001000;
#1 $display("%b", po);
# 1  pi=13'b1001001001001;
#1 $display("%b", po);
# 1  pi=13'b1001001001010;
#1 $display("%b", po);
# 1  pi=13'b1001001001011;
#1 $display("%b", po);
# 1  pi=13'b1001001001100;
#1 $display("%b", po);
# 1  pi=13'b1001001001101;
#1 $display("%b", po);
# 1  pi=13'b1001001001110;
#1 $display("%b", po);
# 1  pi=13'b1001001001111;
#1 $display("%b", po);
# 1  pi=13'b1001001010000;
#1 $display("%b", po);
# 1  pi=13'b1001001010001;
#1 $display("%b", po);
# 1  pi=13'b1001001010010;
#1 $display("%b", po);
# 1  pi=13'b1001001010011;
#1 $display("%b", po);
# 1  pi=13'b1001001010100;
#1 $display("%b", po);
# 1  pi=13'b1001001010101;
#1 $display("%b", po);
# 1  pi=13'b1001001010110;
#1 $display("%b", po);
# 1  pi=13'b1001001010111;
#1 $display("%b", po);
# 1  pi=13'b1001001011000;
#1 $display("%b", po);
# 1  pi=13'b1001001011001;
#1 $display("%b", po);
# 1  pi=13'b1001001011010;
#1 $display("%b", po);
# 1  pi=13'b1001001011011;
#1 $display("%b", po);
# 1  pi=13'b1001001011100;
#1 $display("%b", po);
# 1  pi=13'b1001001011101;
#1 $display("%b", po);
# 1  pi=13'b1001001011110;
#1 $display("%b", po);
# 1  pi=13'b1001001011111;
#1 $display("%b", po);
# 1  pi=13'b1001001100000;
#1 $display("%b", po);
# 1  pi=13'b1001001100001;
#1 $display("%b", po);
# 1  pi=13'b1001001100010;
#1 $display("%b", po);
# 1  pi=13'b1001001100011;
#1 $display("%b", po);
# 1  pi=13'b1001001100100;
#1 $display("%b", po);
# 1  pi=13'b1001001100101;
#1 $display("%b", po);
# 1  pi=13'b1001001100110;
#1 $display("%b", po);
# 1  pi=13'b1001001100111;
#1 $display("%b", po);
# 1  pi=13'b1001001101000;
#1 $display("%b", po);
# 1  pi=13'b1001001101001;
#1 $display("%b", po);
# 1  pi=13'b1001001101010;
#1 $display("%b", po);
# 1  pi=13'b1001001101011;
#1 $display("%b", po);
# 1  pi=13'b1001001101100;
#1 $display("%b", po);
# 1  pi=13'b1001001101101;
#1 $display("%b", po);
# 1  pi=13'b1001001101110;
#1 $display("%b", po);
# 1  pi=13'b1001001101111;
#1 $display("%b", po);
# 1  pi=13'b1001001110000;
#1 $display("%b", po);
# 1  pi=13'b1001001110001;
#1 $display("%b", po);
# 1  pi=13'b1001001110010;
#1 $display("%b", po);
# 1  pi=13'b1001001110011;
#1 $display("%b", po);
# 1  pi=13'b1001001110100;
#1 $display("%b", po);
# 1  pi=13'b1001001110101;
#1 $display("%b", po);
# 1  pi=13'b1001001110110;
#1 $display("%b", po);
# 1  pi=13'b1001001110111;
#1 $display("%b", po);
# 1  pi=13'b1001001111000;
#1 $display("%b", po);
# 1  pi=13'b1001001111001;
#1 $display("%b", po);
# 1  pi=13'b1001001111010;
#1 $display("%b", po);
# 1  pi=13'b1001001111011;
#1 $display("%b", po);
# 1  pi=13'b1001001111100;
#1 $display("%b", po);
# 1  pi=13'b1001001111101;
#1 $display("%b", po);
# 1  pi=13'b1001001111110;
#1 $display("%b", po);
# 1  pi=13'b1001001111111;
#1 $display("%b", po);
# 1  pi=13'b1001010000000;
#1 $display("%b", po);
# 1  pi=13'b1001010000001;
#1 $display("%b", po);
# 1  pi=13'b1001010000010;
#1 $display("%b", po);
# 1  pi=13'b1001010000011;
#1 $display("%b", po);
# 1  pi=13'b1001010000100;
#1 $display("%b", po);
# 1  pi=13'b1001010000101;
#1 $display("%b", po);
# 1  pi=13'b1001010000110;
#1 $display("%b", po);
# 1  pi=13'b1001010000111;
#1 $display("%b", po);
# 1  pi=13'b1001010001000;
#1 $display("%b", po);
# 1  pi=13'b1001010001001;
#1 $display("%b", po);
# 1  pi=13'b1001010001010;
#1 $display("%b", po);
# 1  pi=13'b1001010001011;
#1 $display("%b", po);
# 1  pi=13'b1001010001100;
#1 $display("%b", po);
# 1  pi=13'b1001010001101;
#1 $display("%b", po);
# 1  pi=13'b1001010001110;
#1 $display("%b", po);
# 1  pi=13'b1001010001111;
#1 $display("%b", po);
# 1  pi=13'b1001010010000;
#1 $display("%b", po);
# 1  pi=13'b1001010010001;
#1 $display("%b", po);
# 1  pi=13'b1001010010010;
#1 $display("%b", po);
# 1  pi=13'b1001010010011;
#1 $display("%b", po);
# 1  pi=13'b1001010010100;
#1 $display("%b", po);
# 1  pi=13'b1001010010101;
#1 $display("%b", po);
# 1  pi=13'b1001010010110;
#1 $display("%b", po);
# 1  pi=13'b1001010010111;
#1 $display("%b", po);
# 1  pi=13'b1001010011000;
#1 $display("%b", po);
# 1  pi=13'b1001010011001;
#1 $display("%b", po);
# 1  pi=13'b1001010011010;
#1 $display("%b", po);
# 1  pi=13'b1001010011011;
#1 $display("%b", po);
# 1  pi=13'b1001010011100;
#1 $display("%b", po);
# 1  pi=13'b1001010011101;
#1 $display("%b", po);
# 1  pi=13'b1001010011110;
#1 $display("%b", po);
# 1  pi=13'b1001010011111;
#1 $display("%b", po);
# 1  pi=13'b1001010100000;
#1 $display("%b", po);
# 1  pi=13'b1001010100001;
#1 $display("%b", po);
# 1  pi=13'b1001010100010;
#1 $display("%b", po);
# 1  pi=13'b1001010100011;
#1 $display("%b", po);
# 1  pi=13'b1001010100100;
#1 $display("%b", po);
# 1  pi=13'b1001010100101;
#1 $display("%b", po);
# 1  pi=13'b1001010100110;
#1 $display("%b", po);
# 1  pi=13'b1001010100111;
#1 $display("%b", po);
# 1  pi=13'b1001010101000;
#1 $display("%b", po);
# 1  pi=13'b1001010101001;
#1 $display("%b", po);
# 1  pi=13'b1001010101010;
#1 $display("%b", po);
# 1  pi=13'b1001010101011;
#1 $display("%b", po);
# 1  pi=13'b1001010101100;
#1 $display("%b", po);
# 1  pi=13'b1001010101101;
#1 $display("%b", po);
# 1  pi=13'b1001010101110;
#1 $display("%b", po);
# 1  pi=13'b1001010101111;
#1 $display("%b", po);
# 1  pi=13'b1001010110000;
#1 $display("%b", po);
# 1  pi=13'b1001010110001;
#1 $display("%b", po);
# 1  pi=13'b1001010110010;
#1 $display("%b", po);
# 1  pi=13'b1001010110011;
#1 $display("%b", po);
# 1  pi=13'b1001010110100;
#1 $display("%b", po);
# 1  pi=13'b1001010110101;
#1 $display("%b", po);
# 1  pi=13'b1001010110110;
#1 $display("%b", po);
# 1  pi=13'b1001010110111;
#1 $display("%b", po);
# 1  pi=13'b1001010111000;
#1 $display("%b", po);
# 1  pi=13'b1001010111001;
#1 $display("%b", po);
# 1  pi=13'b1001010111010;
#1 $display("%b", po);
# 1  pi=13'b1001010111011;
#1 $display("%b", po);
# 1  pi=13'b1001010111100;
#1 $display("%b", po);
# 1  pi=13'b1001010111101;
#1 $display("%b", po);
# 1  pi=13'b1001010111110;
#1 $display("%b", po);
# 1  pi=13'b1001010111111;
#1 $display("%b", po);
# 1  pi=13'b1001011000000;
#1 $display("%b", po);
# 1  pi=13'b1001011000001;
#1 $display("%b", po);
# 1  pi=13'b1001011000010;
#1 $display("%b", po);
# 1  pi=13'b1001011000011;
#1 $display("%b", po);
# 1  pi=13'b1001011000100;
#1 $display("%b", po);
# 1  pi=13'b1001011000101;
#1 $display("%b", po);
# 1  pi=13'b1001011000110;
#1 $display("%b", po);
# 1  pi=13'b1001011000111;
#1 $display("%b", po);
# 1  pi=13'b1001011001000;
#1 $display("%b", po);
# 1  pi=13'b1001011001001;
#1 $display("%b", po);
# 1  pi=13'b1001011001010;
#1 $display("%b", po);
# 1  pi=13'b1001011001011;
#1 $display("%b", po);
# 1  pi=13'b1001011001100;
#1 $display("%b", po);
# 1  pi=13'b1001011001101;
#1 $display("%b", po);
# 1  pi=13'b1001011001110;
#1 $display("%b", po);
# 1  pi=13'b1001011001111;
#1 $display("%b", po);
# 1  pi=13'b1001011010000;
#1 $display("%b", po);
# 1  pi=13'b1001011010001;
#1 $display("%b", po);
# 1  pi=13'b1001011010010;
#1 $display("%b", po);
# 1  pi=13'b1001011010011;
#1 $display("%b", po);
# 1  pi=13'b1001011010100;
#1 $display("%b", po);
# 1  pi=13'b1001011010101;
#1 $display("%b", po);
# 1  pi=13'b1001011010110;
#1 $display("%b", po);
# 1  pi=13'b1001011010111;
#1 $display("%b", po);
# 1  pi=13'b1001011011000;
#1 $display("%b", po);
# 1  pi=13'b1001011011001;
#1 $display("%b", po);
# 1  pi=13'b1001011011010;
#1 $display("%b", po);
# 1  pi=13'b1001011011011;
#1 $display("%b", po);
# 1  pi=13'b1001011011100;
#1 $display("%b", po);
# 1  pi=13'b1001011011101;
#1 $display("%b", po);
# 1  pi=13'b1001011011110;
#1 $display("%b", po);
# 1  pi=13'b1001011011111;
#1 $display("%b", po);
# 1  pi=13'b1001011100000;
#1 $display("%b", po);
# 1  pi=13'b1001011100001;
#1 $display("%b", po);
# 1  pi=13'b1001011100010;
#1 $display("%b", po);
# 1  pi=13'b1001011100011;
#1 $display("%b", po);
# 1  pi=13'b1001011100100;
#1 $display("%b", po);
# 1  pi=13'b1001011100101;
#1 $display("%b", po);
# 1  pi=13'b1001011100110;
#1 $display("%b", po);
# 1  pi=13'b1001011100111;
#1 $display("%b", po);
# 1  pi=13'b1001011101000;
#1 $display("%b", po);
# 1  pi=13'b1001011101001;
#1 $display("%b", po);
# 1  pi=13'b1001011101010;
#1 $display("%b", po);
# 1  pi=13'b1001011101011;
#1 $display("%b", po);
# 1  pi=13'b1001011101100;
#1 $display("%b", po);
# 1  pi=13'b1001011101101;
#1 $display("%b", po);
# 1  pi=13'b1001011101110;
#1 $display("%b", po);
# 1  pi=13'b1001011101111;
#1 $display("%b", po);
# 1  pi=13'b1001011110000;
#1 $display("%b", po);
# 1  pi=13'b1001011110001;
#1 $display("%b", po);
# 1  pi=13'b1001011110010;
#1 $display("%b", po);
# 1  pi=13'b1001011110011;
#1 $display("%b", po);
# 1  pi=13'b1001011110100;
#1 $display("%b", po);
# 1  pi=13'b1001011110101;
#1 $display("%b", po);
# 1  pi=13'b1001011110110;
#1 $display("%b", po);
# 1  pi=13'b1001011110111;
#1 $display("%b", po);
# 1  pi=13'b1001011111000;
#1 $display("%b", po);
# 1  pi=13'b1001011111001;
#1 $display("%b", po);
# 1  pi=13'b1001011111010;
#1 $display("%b", po);
# 1  pi=13'b1001011111011;
#1 $display("%b", po);
# 1  pi=13'b1001011111100;
#1 $display("%b", po);
# 1  pi=13'b1001011111101;
#1 $display("%b", po);
# 1  pi=13'b1001011111110;
#1 $display("%b", po);
# 1  pi=13'b1001011111111;
#1 $display("%b", po);
# 1  pi=13'b1001100000000;
#1 $display("%b", po);
# 1  pi=13'b1001100000001;
#1 $display("%b", po);
# 1  pi=13'b1001100000010;
#1 $display("%b", po);
# 1  pi=13'b1001100000011;
#1 $display("%b", po);
# 1  pi=13'b1001100000100;
#1 $display("%b", po);
# 1  pi=13'b1001100000101;
#1 $display("%b", po);
# 1  pi=13'b1001100000110;
#1 $display("%b", po);
# 1  pi=13'b1001100000111;
#1 $display("%b", po);
# 1  pi=13'b1001100001000;
#1 $display("%b", po);
# 1  pi=13'b1001100001001;
#1 $display("%b", po);
# 1  pi=13'b1001100001010;
#1 $display("%b", po);
# 1  pi=13'b1001100001011;
#1 $display("%b", po);
# 1  pi=13'b1001100001100;
#1 $display("%b", po);
# 1  pi=13'b1001100001101;
#1 $display("%b", po);
# 1  pi=13'b1001100001110;
#1 $display("%b", po);
# 1  pi=13'b1001100001111;
#1 $display("%b", po);
# 1  pi=13'b1001100010000;
#1 $display("%b", po);
# 1  pi=13'b1001100010001;
#1 $display("%b", po);
# 1  pi=13'b1001100010010;
#1 $display("%b", po);
# 1  pi=13'b1001100010011;
#1 $display("%b", po);
# 1  pi=13'b1001100010100;
#1 $display("%b", po);
# 1  pi=13'b1001100010101;
#1 $display("%b", po);
# 1  pi=13'b1001100010110;
#1 $display("%b", po);
# 1  pi=13'b1001100010111;
#1 $display("%b", po);
# 1  pi=13'b1001100011000;
#1 $display("%b", po);
# 1  pi=13'b1001100011001;
#1 $display("%b", po);
# 1  pi=13'b1001100011010;
#1 $display("%b", po);
# 1  pi=13'b1001100011011;
#1 $display("%b", po);
# 1  pi=13'b1001100011100;
#1 $display("%b", po);
# 1  pi=13'b1001100011101;
#1 $display("%b", po);
# 1  pi=13'b1001100011110;
#1 $display("%b", po);
# 1  pi=13'b1001100011111;
#1 $display("%b", po);
# 1  pi=13'b1001100100000;
#1 $display("%b", po);
# 1  pi=13'b1001100100001;
#1 $display("%b", po);
# 1  pi=13'b1001100100010;
#1 $display("%b", po);
# 1  pi=13'b1001100100011;
#1 $display("%b", po);
# 1  pi=13'b1001100100100;
#1 $display("%b", po);
# 1  pi=13'b1001100100101;
#1 $display("%b", po);
# 1  pi=13'b1001100100110;
#1 $display("%b", po);
# 1  pi=13'b1001100100111;
#1 $display("%b", po);
# 1  pi=13'b1001100101000;
#1 $display("%b", po);
# 1  pi=13'b1001100101001;
#1 $display("%b", po);
# 1  pi=13'b1001100101010;
#1 $display("%b", po);
# 1  pi=13'b1001100101011;
#1 $display("%b", po);
# 1  pi=13'b1001100101100;
#1 $display("%b", po);
# 1  pi=13'b1001100101101;
#1 $display("%b", po);
# 1  pi=13'b1001100101110;
#1 $display("%b", po);
# 1  pi=13'b1001100101111;
#1 $display("%b", po);
# 1  pi=13'b1001100110000;
#1 $display("%b", po);
# 1  pi=13'b1001100110001;
#1 $display("%b", po);
# 1  pi=13'b1001100110010;
#1 $display("%b", po);
# 1  pi=13'b1001100110011;
#1 $display("%b", po);
# 1  pi=13'b1001100110100;
#1 $display("%b", po);
# 1  pi=13'b1001100110101;
#1 $display("%b", po);
# 1  pi=13'b1001100110110;
#1 $display("%b", po);
# 1  pi=13'b1001100110111;
#1 $display("%b", po);
# 1  pi=13'b1001100111000;
#1 $display("%b", po);
# 1  pi=13'b1001100111001;
#1 $display("%b", po);
# 1  pi=13'b1001100111010;
#1 $display("%b", po);
# 1  pi=13'b1001100111011;
#1 $display("%b", po);
# 1  pi=13'b1001100111100;
#1 $display("%b", po);
# 1  pi=13'b1001100111101;
#1 $display("%b", po);
# 1  pi=13'b1001100111110;
#1 $display("%b", po);
# 1  pi=13'b1001100111111;
#1 $display("%b", po);
# 1  pi=13'b1001101000000;
#1 $display("%b", po);
# 1  pi=13'b1001101000001;
#1 $display("%b", po);
# 1  pi=13'b1001101000010;
#1 $display("%b", po);
# 1  pi=13'b1001101000011;
#1 $display("%b", po);
# 1  pi=13'b1001101000100;
#1 $display("%b", po);
# 1  pi=13'b1001101000101;
#1 $display("%b", po);
# 1  pi=13'b1001101000110;
#1 $display("%b", po);
# 1  pi=13'b1001101000111;
#1 $display("%b", po);
# 1  pi=13'b1001101001000;
#1 $display("%b", po);
# 1  pi=13'b1001101001001;
#1 $display("%b", po);
# 1  pi=13'b1001101001010;
#1 $display("%b", po);
# 1  pi=13'b1001101001011;
#1 $display("%b", po);
# 1  pi=13'b1001101001100;
#1 $display("%b", po);
# 1  pi=13'b1001101001101;
#1 $display("%b", po);
# 1  pi=13'b1001101001110;
#1 $display("%b", po);
# 1  pi=13'b1001101001111;
#1 $display("%b", po);
# 1  pi=13'b1001101010000;
#1 $display("%b", po);
# 1  pi=13'b1001101010001;
#1 $display("%b", po);
# 1  pi=13'b1001101010010;
#1 $display("%b", po);
# 1  pi=13'b1001101010011;
#1 $display("%b", po);
# 1  pi=13'b1001101010100;
#1 $display("%b", po);
# 1  pi=13'b1001101010101;
#1 $display("%b", po);
# 1  pi=13'b1001101010110;
#1 $display("%b", po);
# 1  pi=13'b1001101010111;
#1 $display("%b", po);
# 1  pi=13'b1001101011000;
#1 $display("%b", po);
# 1  pi=13'b1001101011001;
#1 $display("%b", po);
# 1  pi=13'b1001101011010;
#1 $display("%b", po);
# 1  pi=13'b1001101011011;
#1 $display("%b", po);
# 1  pi=13'b1001101011100;
#1 $display("%b", po);
# 1  pi=13'b1001101011101;
#1 $display("%b", po);
# 1  pi=13'b1001101011110;
#1 $display("%b", po);
# 1  pi=13'b1001101011111;
#1 $display("%b", po);
# 1  pi=13'b1001101100000;
#1 $display("%b", po);
# 1  pi=13'b1001101100001;
#1 $display("%b", po);
# 1  pi=13'b1001101100010;
#1 $display("%b", po);
# 1  pi=13'b1001101100011;
#1 $display("%b", po);
# 1  pi=13'b1001101100100;
#1 $display("%b", po);
# 1  pi=13'b1001101100101;
#1 $display("%b", po);
# 1  pi=13'b1001101100110;
#1 $display("%b", po);
# 1  pi=13'b1001101100111;
#1 $display("%b", po);
# 1  pi=13'b1001101101000;
#1 $display("%b", po);
# 1  pi=13'b1001101101001;
#1 $display("%b", po);
# 1  pi=13'b1001101101010;
#1 $display("%b", po);
# 1  pi=13'b1001101101011;
#1 $display("%b", po);
# 1  pi=13'b1001101101100;
#1 $display("%b", po);
# 1  pi=13'b1001101101101;
#1 $display("%b", po);
# 1  pi=13'b1001101101110;
#1 $display("%b", po);
# 1  pi=13'b1001101101111;
#1 $display("%b", po);
# 1  pi=13'b1001101110000;
#1 $display("%b", po);
# 1  pi=13'b1001101110001;
#1 $display("%b", po);
# 1  pi=13'b1001101110010;
#1 $display("%b", po);
# 1  pi=13'b1001101110011;
#1 $display("%b", po);
# 1  pi=13'b1001101110100;
#1 $display("%b", po);
# 1  pi=13'b1001101110101;
#1 $display("%b", po);
# 1  pi=13'b1001101110110;
#1 $display("%b", po);
# 1  pi=13'b1001101110111;
#1 $display("%b", po);
# 1  pi=13'b1001101111000;
#1 $display("%b", po);
# 1  pi=13'b1001101111001;
#1 $display("%b", po);
# 1  pi=13'b1001101111010;
#1 $display("%b", po);
# 1  pi=13'b1001101111011;
#1 $display("%b", po);
# 1  pi=13'b1001101111100;
#1 $display("%b", po);
# 1  pi=13'b1001101111101;
#1 $display("%b", po);
# 1  pi=13'b1001101111110;
#1 $display("%b", po);
# 1  pi=13'b1001101111111;
#1 $display("%b", po);
# 1  pi=13'b1001110000000;
#1 $display("%b", po);
# 1  pi=13'b1001110000001;
#1 $display("%b", po);
# 1  pi=13'b1001110000010;
#1 $display("%b", po);
# 1  pi=13'b1001110000011;
#1 $display("%b", po);
# 1  pi=13'b1001110000100;
#1 $display("%b", po);
# 1  pi=13'b1001110000101;
#1 $display("%b", po);
# 1  pi=13'b1001110000110;
#1 $display("%b", po);
# 1  pi=13'b1001110000111;
#1 $display("%b", po);
# 1  pi=13'b1001110001000;
#1 $display("%b", po);
# 1  pi=13'b1001110001001;
#1 $display("%b", po);
# 1  pi=13'b1001110001010;
#1 $display("%b", po);
# 1  pi=13'b1001110001011;
#1 $display("%b", po);
# 1  pi=13'b1001110001100;
#1 $display("%b", po);
# 1  pi=13'b1001110001101;
#1 $display("%b", po);
# 1  pi=13'b1001110001110;
#1 $display("%b", po);
# 1  pi=13'b1001110001111;
#1 $display("%b", po);
# 1  pi=13'b1001110010000;
#1 $display("%b", po);
# 1  pi=13'b1001110010001;
#1 $display("%b", po);
# 1  pi=13'b1001110010010;
#1 $display("%b", po);
# 1  pi=13'b1001110010011;
#1 $display("%b", po);
# 1  pi=13'b1001110010100;
#1 $display("%b", po);
# 1  pi=13'b1001110010101;
#1 $display("%b", po);
# 1  pi=13'b1001110010110;
#1 $display("%b", po);
# 1  pi=13'b1001110010111;
#1 $display("%b", po);
# 1  pi=13'b1001110011000;
#1 $display("%b", po);
# 1  pi=13'b1001110011001;
#1 $display("%b", po);
# 1  pi=13'b1001110011010;
#1 $display("%b", po);
# 1  pi=13'b1001110011011;
#1 $display("%b", po);
# 1  pi=13'b1001110011100;
#1 $display("%b", po);
# 1  pi=13'b1001110011101;
#1 $display("%b", po);
# 1  pi=13'b1001110011110;
#1 $display("%b", po);
# 1  pi=13'b1001110011111;
#1 $display("%b", po);
# 1  pi=13'b1001110100000;
#1 $display("%b", po);
# 1  pi=13'b1001110100001;
#1 $display("%b", po);
# 1  pi=13'b1001110100010;
#1 $display("%b", po);
# 1  pi=13'b1001110100011;
#1 $display("%b", po);
# 1  pi=13'b1001110100100;
#1 $display("%b", po);
# 1  pi=13'b1001110100101;
#1 $display("%b", po);
# 1  pi=13'b1001110100110;
#1 $display("%b", po);
# 1  pi=13'b1001110100111;
#1 $display("%b", po);
# 1  pi=13'b1001110101000;
#1 $display("%b", po);
# 1  pi=13'b1001110101001;
#1 $display("%b", po);
# 1  pi=13'b1001110101010;
#1 $display("%b", po);
# 1  pi=13'b1001110101011;
#1 $display("%b", po);
# 1  pi=13'b1001110101100;
#1 $display("%b", po);
# 1  pi=13'b1001110101101;
#1 $display("%b", po);
# 1  pi=13'b1001110101110;
#1 $display("%b", po);
# 1  pi=13'b1001110101111;
#1 $display("%b", po);
# 1  pi=13'b1001110110000;
#1 $display("%b", po);
# 1  pi=13'b1001110110001;
#1 $display("%b", po);
# 1  pi=13'b1001110110010;
#1 $display("%b", po);
# 1  pi=13'b1001110110011;
#1 $display("%b", po);
# 1  pi=13'b1001110110100;
#1 $display("%b", po);
# 1  pi=13'b1001110110101;
#1 $display("%b", po);
# 1  pi=13'b1001110110110;
#1 $display("%b", po);
# 1  pi=13'b1001110110111;
#1 $display("%b", po);
# 1  pi=13'b1001110111000;
#1 $display("%b", po);
# 1  pi=13'b1001110111001;
#1 $display("%b", po);
# 1  pi=13'b1001110111010;
#1 $display("%b", po);
# 1  pi=13'b1001110111011;
#1 $display("%b", po);
# 1  pi=13'b1001110111100;
#1 $display("%b", po);
# 1  pi=13'b1001110111101;
#1 $display("%b", po);
# 1  pi=13'b1001110111110;
#1 $display("%b", po);
# 1  pi=13'b1001110111111;
#1 $display("%b", po);
# 1  pi=13'b1001111000000;
#1 $display("%b", po);
# 1  pi=13'b1001111000001;
#1 $display("%b", po);
# 1  pi=13'b1001111000010;
#1 $display("%b", po);
# 1  pi=13'b1001111000011;
#1 $display("%b", po);
# 1  pi=13'b1001111000100;
#1 $display("%b", po);
# 1  pi=13'b1001111000101;
#1 $display("%b", po);
# 1  pi=13'b1001111000110;
#1 $display("%b", po);
# 1  pi=13'b1001111000111;
#1 $display("%b", po);
# 1  pi=13'b1001111001000;
#1 $display("%b", po);
# 1  pi=13'b1001111001001;
#1 $display("%b", po);
# 1  pi=13'b1001111001010;
#1 $display("%b", po);
# 1  pi=13'b1001111001011;
#1 $display("%b", po);
# 1  pi=13'b1001111001100;
#1 $display("%b", po);
# 1  pi=13'b1001111001101;
#1 $display("%b", po);
# 1  pi=13'b1001111001110;
#1 $display("%b", po);
# 1  pi=13'b1001111001111;
#1 $display("%b", po);
# 1  pi=13'b1001111010000;
#1 $display("%b", po);
# 1  pi=13'b1001111010001;
#1 $display("%b", po);
# 1  pi=13'b1001111010010;
#1 $display("%b", po);
# 1  pi=13'b1001111010011;
#1 $display("%b", po);
# 1  pi=13'b1001111010100;
#1 $display("%b", po);
# 1  pi=13'b1001111010101;
#1 $display("%b", po);
# 1  pi=13'b1001111010110;
#1 $display("%b", po);
# 1  pi=13'b1001111010111;
#1 $display("%b", po);
# 1  pi=13'b1001111011000;
#1 $display("%b", po);
# 1  pi=13'b1001111011001;
#1 $display("%b", po);
# 1  pi=13'b1001111011010;
#1 $display("%b", po);
# 1  pi=13'b1001111011011;
#1 $display("%b", po);
# 1  pi=13'b1001111011100;
#1 $display("%b", po);
# 1  pi=13'b1001111011101;
#1 $display("%b", po);
# 1  pi=13'b1001111011110;
#1 $display("%b", po);
# 1  pi=13'b1001111011111;
#1 $display("%b", po);
# 1  pi=13'b1001111100000;
#1 $display("%b", po);
# 1  pi=13'b1001111100001;
#1 $display("%b", po);
# 1  pi=13'b1001111100010;
#1 $display("%b", po);
# 1  pi=13'b1001111100011;
#1 $display("%b", po);
# 1  pi=13'b1001111100100;
#1 $display("%b", po);
# 1  pi=13'b1001111100101;
#1 $display("%b", po);
# 1  pi=13'b1001111100110;
#1 $display("%b", po);
# 1  pi=13'b1001111100111;
#1 $display("%b", po);
# 1  pi=13'b1001111101000;
#1 $display("%b", po);
# 1  pi=13'b1001111101001;
#1 $display("%b", po);
# 1  pi=13'b1001111101010;
#1 $display("%b", po);
# 1  pi=13'b1001111101011;
#1 $display("%b", po);
# 1  pi=13'b1001111101100;
#1 $display("%b", po);
# 1  pi=13'b1001111101101;
#1 $display("%b", po);
# 1  pi=13'b1001111101110;
#1 $display("%b", po);
# 1  pi=13'b1001111101111;
#1 $display("%b", po);
# 1  pi=13'b1001111110000;
#1 $display("%b", po);
# 1  pi=13'b1001111110001;
#1 $display("%b", po);
# 1  pi=13'b1001111110010;
#1 $display("%b", po);
# 1  pi=13'b1001111110011;
#1 $display("%b", po);
# 1  pi=13'b1001111110100;
#1 $display("%b", po);
# 1  pi=13'b1001111110101;
#1 $display("%b", po);
# 1  pi=13'b1001111110110;
#1 $display("%b", po);
# 1  pi=13'b1001111110111;
#1 $display("%b", po);
# 1  pi=13'b1001111111000;
#1 $display("%b", po);
# 1  pi=13'b1001111111001;
#1 $display("%b", po);
# 1  pi=13'b1001111111010;
#1 $display("%b", po);
# 1  pi=13'b1001111111011;
#1 $display("%b", po);
# 1  pi=13'b1001111111100;
#1 $display("%b", po);
# 1  pi=13'b1001111111101;
#1 $display("%b", po);
# 1  pi=13'b1001111111110;
#1 $display("%b", po);
# 1  pi=13'b1001111111111;
#1 $display("%b", po);
# 1  pi=13'b1010000000000;
#1 $display("%b", po);
# 1  pi=13'b1010000000001;
#1 $display("%b", po);
# 1  pi=13'b1010000000010;
#1 $display("%b", po);
# 1  pi=13'b1010000000011;
#1 $display("%b", po);
# 1  pi=13'b1010000000100;
#1 $display("%b", po);
# 1  pi=13'b1010000000101;
#1 $display("%b", po);
# 1  pi=13'b1010000000110;
#1 $display("%b", po);
# 1  pi=13'b1010000000111;
#1 $display("%b", po);
# 1  pi=13'b1010000001000;
#1 $display("%b", po);
# 1  pi=13'b1010000001001;
#1 $display("%b", po);
# 1  pi=13'b1010000001010;
#1 $display("%b", po);
# 1  pi=13'b1010000001011;
#1 $display("%b", po);
# 1  pi=13'b1010000001100;
#1 $display("%b", po);
# 1  pi=13'b1010000001101;
#1 $display("%b", po);
# 1  pi=13'b1010000001110;
#1 $display("%b", po);
# 1  pi=13'b1010000001111;
#1 $display("%b", po);
# 1  pi=13'b1010000010000;
#1 $display("%b", po);
# 1  pi=13'b1010000010001;
#1 $display("%b", po);
# 1  pi=13'b1010000010010;
#1 $display("%b", po);
# 1  pi=13'b1010000010011;
#1 $display("%b", po);
# 1  pi=13'b1010000010100;
#1 $display("%b", po);
# 1  pi=13'b1010000010101;
#1 $display("%b", po);
# 1  pi=13'b1010000010110;
#1 $display("%b", po);
# 1  pi=13'b1010000010111;
#1 $display("%b", po);
# 1  pi=13'b1010000011000;
#1 $display("%b", po);
# 1  pi=13'b1010000011001;
#1 $display("%b", po);
# 1  pi=13'b1010000011010;
#1 $display("%b", po);
# 1  pi=13'b1010000011011;
#1 $display("%b", po);
# 1  pi=13'b1010000011100;
#1 $display("%b", po);
# 1  pi=13'b1010000011101;
#1 $display("%b", po);
# 1  pi=13'b1010000011110;
#1 $display("%b", po);
# 1  pi=13'b1010000011111;
#1 $display("%b", po);
# 1  pi=13'b1010000100000;
#1 $display("%b", po);
# 1  pi=13'b1010000100001;
#1 $display("%b", po);
# 1  pi=13'b1010000100010;
#1 $display("%b", po);
# 1  pi=13'b1010000100011;
#1 $display("%b", po);
# 1  pi=13'b1010000100100;
#1 $display("%b", po);
# 1  pi=13'b1010000100101;
#1 $display("%b", po);
# 1  pi=13'b1010000100110;
#1 $display("%b", po);
# 1  pi=13'b1010000100111;
#1 $display("%b", po);
# 1  pi=13'b1010000101000;
#1 $display("%b", po);
# 1  pi=13'b1010000101001;
#1 $display("%b", po);
# 1  pi=13'b1010000101010;
#1 $display("%b", po);
# 1  pi=13'b1010000101011;
#1 $display("%b", po);
# 1  pi=13'b1010000101100;
#1 $display("%b", po);
# 1  pi=13'b1010000101101;
#1 $display("%b", po);
# 1  pi=13'b1010000101110;
#1 $display("%b", po);
# 1  pi=13'b1010000101111;
#1 $display("%b", po);
# 1  pi=13'b1010000110000;
#1 $display("%b", po);
# 1  pi=13'b1010000110001;
#1 $display("%b", po);
# 1  pi=13'b1010000110010;
#1 $display("%b", po);
# 1  pi=13'b1010000110011;
#1 $display("%b", po);
# 1  pi=13'b1010000110100;
#1 $display("%b", po);
# 1  pi=13'b1010000110101;
#1 $display("%b", po);
# 1  pi=13'b1010000110110;
#1 $display("%b", po);
# 1  pi=13'b1010000110111;
#1 $display("%b", po);
# 1  pi=13'b1010000111000;
#1 $display("%b", po);
# 1  pi=13'b1010000111001;
#1 $display("%b", po);
# 1  pi=13'b1010000111010;
#1 $display("%b", po);
# 1  pi=13'b1010000111011;
#1 $display("%b", po);
# 1  pi=13'b1010000111100;
#1 $display("%b", po);
# 1  pi=13'b1010000111101;
#1 $display("%b", po);
# 1  pi=13'b1010000111110;
#1 $display("%b", po);
# 1  pi=13'b1010000111111;
#1 $display("%b", po);
# 1  pi=13'b1010001000000;
#1 $display("%b", po);
# 1  pi=13'b1010001000001;
#1 $display("%b", po);
# 1  pi=13'b1010001000010;
#1 $display("%b", po);
# 1  pi=13'b1010001000011;
#1 $display("%b", po);
# 1  pi=13'b1010001000100;
#1 $display("%b", po);
# 1  pi=13'b1010001000101;
#1 $display("%b", po);
# 1  pi=13'b1010001000110;
#1 $display("%b", po);
# 1  pi=13'b1010001000111;
#1 $display("%b", po);
# 1  pi=13'b1010001001000;
#1 $display("%b", po);
# 1  pi=13'b1010001001001;
#1 $display("%b", po);
# 1  pi=13'b1010001001010;
#1 $display("%b", po);
# 1  pi=13'b1010001001011;
#1 $display("%b", po);
# 1  pi=13'b1010001001100;
#1 $display("%b", po);
# 1  pi=13'b1010001001101;
#1 $display("%b", po);
# 1  pi=13'b1010001001110;
#1 $display("%b", po);
# 1  pi=13'b1010001001111;
#1 $display("%b", po);
# 1  pi=13'b1010001010000;
#1 $display("%b", po);
# 1  pi=13'b1010001010001;
#1 $display("%b", po);
# 1  pi=13'b1010001010010;
#1 $display("%b", po);
# 1  pi=13'b1010001010011;
#1 $display("%b", po);
# 1  pi=13'b1010001010100;
#1 $display("%b", po);
# 1  pi=13'b1010001010101;
#1 $display("%b", po);
# 1  pi=13'b1010001010110;
#1 $display("%b", po);
# 1  pi=13'b1010001010111;
#1 $display("%b", po);
# 1  pi=13'b1010001011000;
#1 $display("%b", po);
# 1  pi=13'b1010001011001;
#1 $display("%b", po);
# 1  pi=13'b1010001011010;
#1 $display("%b", po);
# 1  pi=13'b1010001011011;
#1 $display("%b", po);
# 1  pi=13'b1010001011100;
#1 $display("%b", po);
# 1  pi=13'b1010001011101;
#1 $display("%b", po);
# 1  pi=13'b1010001011110;
#1 $display("%b", po);
# 1  pi=13'b1010001011111;
#1 $display("%b", po);
# 1  pi=13'b1010001100000;
#1 $display("%b", po);
# 1  pi=13'b1010001100001;
#1 $display("%b", po);
# 1  pi=13'b1010001100010;
#1 $display("%b", po);
# 1  pi=13'b1010001100011;
#1 $display("%b", po);
# 1  pi=13'b1010001100100;
#1 $display("%b", po);
# 1  pi=13'b1010001100101;
#1 $display("%b", po);
# 1  pi=13'b1010001100110;
#1 $display("%b", po);
# 1  pi=13'b1010001100111;
#1 $display("%b", po);
# 1  pi=13'b1010001101000;
#1 $display("%b", po);
# 1  pi=13'b1010001101001;
#1 $display("%b", po);
# 1  pi=13'b1010001101010;
#1 $display("%b", po);
# 1  pi=13'b1010001101011;
#1 $display("%b", po);
# 1  pi=13'b1010001101100;
#1 $display("%b", po);
# 1  pi=13'b1010001101101;
#1 $display("%b", po);
# 1  pi=13'b1010001101110;
#1 $display("%b", po);
# 1  pi=13'b1010001101111;
#1 $display("%b", po);
# 1  pi=13'b1010001110000;
#1 $display("%b", po);
# 1  pi=13'b1010001110001;
#1 $display("%b", po);
# 1  pi=13'b1010001110010;
#1 $display("%b", po);
# 1  pi=13'b1010001110011;
#1 $display("%b", po);
# 1  pi=13'b1010001110100;
#1 $display("%b", po);
# 1  pi=13'b1010001110101;
#1 $display("%b", po);
# 1  pi=13'b1010001110110;
#1 $display("%b", po);
# 1  pi=13'b1010001110111;
#1 $display("%b", po);
# 1  pi=13'b1010001111000;
#1 $display("%b", po);
# 1  pi=13'b1010001111001;
#1 $display("%b", po);
# 1  pi=13'b1010001111010;
#1 $display("%b", po);
# 1  pi=13'b1010001111011;
#1 $display("%b", po);
# 1  pi=13'b1010001111100;
#1 $display("%b", po);
# 1  pi=13'b1010001111101;
#1 $display("%b", po);
# 1  pi=13'b1010001111110;
#1 $display("%b", po);
# 1  pi=13'b1010001111111;
#1 $display("%b", po);
# 1  pi=13'b1010010000000;
#1 $display("%b", po);
# 1  pi=13'b1010010000001;
#1 $display("%b", po);
# 1  pi=13'b1010010000010;
#1 $display("%b", po);
# 1  pi=13'b1010010000011;
#1 $display("%b", po);
# 1  pi=13'b1010010000100;
#1 $display("%b", po);
# 1  pi=13'b1010010000101;
#1 $display("%b", po);
# 1  pi=13'b1010010000110;
#1 $display("%b", po);
# 1  pi=13'b1010010000111;
#1 $display("%b", po);
# 1  pi=13'b1010010001000;
#1 $display("%b", po);
# 1  pi=13'b1010010001001;
#1 $display("%b", po);
# 1  pi=13'b1010010001010;
#1 $display("%b", po);
# 1  pi=13'b1010010001011;
#1 $display("%b", po);
# 1  pi=13'b1010010001100;
#1 $display("%b", po);
# 1  pi=13'b1010010001101;
#1 $display("%b", po);
# 1  pi=13'b1010010001110;
#1 $display("%b", po);
# 1  pi=13'b1010010001111;
#1 $display("%b", po);
# 1  pi=13'b1010010010000;
#1 $display("%b", po);
# 1  pi=13'b1010010010001;
#1 $display("%b", po);
# 1  pi=13'b1010010010010;
#1 $display("%b", po);
# 1  pi=13'b1010010010011;
#1 $display("%b", po);
# 1  pi=13'b1010010010100;
#1 $display("%b", po);
# 1  pi=13'b1010010010101;
#1 $display("%b", po);
# 1  pi=13'b1010010010110;
#1 $display("%b", po);
# 1  pi=13'b1010010010111;
#1 $display("%b", po);
# 1  pi=13'b1010010011000;
#1 $display("%b", po);
# 1  pi=13'b1010010011001;
#1 $display("%b", po);
# 1  pi=13'b1010010011010;
#1 $display("%b", po);
# 1  pi=13'b1010010011011;
#1 $display("%b", po);
# 1  pi=13'b1010010011100;
#1 $display("%b", po);
# 1  pi=13'b1010010011101;
#1 $display("%b", po);
# 1  pi=13'b1010010011110;
#1 $display("%b", po);
# 1  pi=13'b1010010011111;
#1 $display("%b", po);
# 1  pi=13'b1010010100000;
#1 $display("%b", po);
# 1  pi=13'b1010010100001;
#1 $display("%b", po);
# 1  pi=13'b1010010100010;
#1 $display("%b", po);
# 1  pi=13'b1010010100011;
#1 $display("%b", po);
# 1  pi=13'b1010010100100;
#1 $display("%b", po);
# 1  pi=13'b1010010100101;
#1 $display("%b", po);
# 1  pi=13'b1010010100110;
#1 $display("%b", po);
# 1  pi=13'b1010010100111;
#1 $display("%b", po);
# 1  pi=13'b1010010101000;
#1 $display("%b", po);
# 1  pi=13'b1010010101001;
#1 $display("%b", po);
# 1  pi=13'b1010010101010;
#1 $display("%b", po);
# 1  pi=13'b1010010101011;
#1 $display("%b", po);
# 1  pi=13'b1010010101100;
#1 $display("%b", po);
# 1  pi=13'b1010010101101;
#1 $display("%b", po);
# 1  pi=13'b1010010101110;
#1 $display("%b", po);
# 1  pi=13'b1010010101111;
#1 $display("%b", po);
# 1  pi=13'b1010010110000;
#1 $display("%b", po);
# 1  pi=13'b1010010110001;
#1 $display("%b", po);
# 1  pi=13'b1010010110010;
#1 $display("%b", po);
# 1  pi=13'b1010010110011;
#1 $display("%b", po);
# 1  pi=13'b1010010110100;
#1 $display("%b", po);
# 1  pi=13'b1010010110101;
#1 $display("%b", po);
# 1  pi=13'b1010010110110;
#1 $display("%b", po);
# 1  pi=13'b1010010110111;
#1 $display("%b", po);
# 1  pi=13'b1010010111000;
#1 $display("%b", po);
# 1  pi=13'b1010010111001;
#1 $display("%b", po);
# 1  pi=13'b1010010111010;
#1 $display("%b", po);
# 1  pi=13'b1010010111011;
#1 $display("%b", po);
# 1  pi=13'b1010010111100;
#1 $display("%b", po);
# 1  pi=13'b1010010111101;
#1 $display("%b", po);
# 1  pi=13'b1010010111110;
#1 $display("%b", po);
# 1  pi=13'b1010010111111;
#1 $display("%b", po);
# 1  pi=13'b1010011000000;
#1 $display("%b", po);
# 1  pi=13'b1010011000001;
#1 $display("%b", po);
# 1  pi=13'b1010011000010;
#1 $display("%b", po);
# 1  pi=13'b1010011000011;
#1 $display("%b", po);
# 1  pi=13'b1010011000100;
#1 $display("%b", po);
# 1  pi=13'b1010011000101;
#1 $display("%b", po);
# 1  pi=13'b1010011000110;
#1 $display("%b", po);
# 1  pi=13'b1010011000111;
#1 $display("%b", po);
# 1  pi=13'b1010011001000;
#1 $display("%b", po);
# 1  pi=13'b1010011001001;
#1 $display("%b", po);
# 1  pi=13'b1010011001010;
#1 $display("%b", po);
# 1  pi=13'b1010011001011;
#1 $display("%b", po);
# 1  pi=13'b1010011001100;
#1 $display("%b", po);
# 1  pi=13'b1010011001101;
#1 $display("%b", po);
# 1  pi=13'b1010011001110;
#1 $display("%b", po);
# 1  pi=13'b1010011001111;
#1 $display("%b", po);
# 1  pi=13'b1010011010000;
#1 $display("%b", po);
# 1  pi=13'b1010011010001;
#1 $display("%b", po);
# 1  pi=13'b1010011010010;
#1 $display("%b", po);
# 1  pi=13'b1010011010011;
#1 $display("%b", po);
# 1  pi=13'b1010011010100;
#1 $display("%b", po);
# 1  pi=13'b1010011010101;
#1 $display("%b", po);
# 1  pi=13'b1010011010110;
#1 $display("%b", po);
# 1  pi=13'b1010011010111;
#1 $display("%b", po);
# 1  pi=13'b1010011011000;
#1 $display("%b", po);
# 1  pi=13'b1010011011001;
#1 $display("%b", po);
# 1  pi=13'b1010011011010;
#1 $display("%b", po);
# 1  pi=13'b1010011011011;
#1 $display("%b", po);
# 1  pi=13'b1010011011100;
#1 $display("%b", po);
# 1  pi=13'b1010011011101;
#1 $display("%b", po);
# 1  pi=13'b1010011011110;
#1 $display("%b", po);
# 1  pi=13'b1010011011111;
#1 $display("%b", po);
# 1  pi=13'b1010011100000;
#1 $display("%b", po);
# 1  pi=13'b1010011100001;
#1 $display("%b", po);
# 1  pi=13'b1010011100010;
#1 $display("%b", po);
# 1  pi=13'b1010011100011;
#1 $display("%b", po);
# 1  pi=13'b1010011100100;
#1 $display("%b", po);
# 1  pi=13'b1010011100101;
#1 $display("%b", po);
# 1  pi=13'b1010011100110;
#1 $display("%b", po);
# 1  pi=13'b1010011100111;
#1 $display("%b", po);
# 1  pi=13'b1010011101000;
#1 $display("%b", po);
# 1  pi=13'b1010011101001;
#1 $display("%b", po);
# 1  pi=13'b1010011101010;
#1 $display("%b", po);
# 1  pi=13'b1010011101011;
#1 $display("%b", po);
# 1  pi=13'b1010011101100;
#1 $display("%b", po);
# 1  pi=13'b1010011101101;
#1 $display("%b", po);
# 1  pi=13'b1010011101110;
#1 $display("%b", po);
# 1  pi=13'b1010011101111;
#1 $display("%b", po);
# 1  pi=13'b1010011110000;
#1 $display("%b", po);
# 1  pi=13'b1010011110001;
#1 $display("%b", po);
# 1  pi=13'b1010011110010;
#1 $display("%b", po);
# 1  pi=13'b1010011110011;
#1 $display("%b", po);
# 1  pi=13'b1010011110100;
#1 $display("%b", po);
# 1  pi=13'b1010011110101;
#1 $display("%b", po);
# 1  pi=13'b1010011110110;
#1 $display("%b", po);
# 1  pi=13'b1010011110111;
#1 $display("%b", po);
# 1  pi=13'b1010011111000;
#1 $display("%b", po);
# 1  pi=13'b1010011111001;
#1 $display("%b", po);
# 1  pi=13'b1010011111010;
#1 $display("%b", po);
# 1  pi=13'b1010011111011;
#1 $display("%b", po);
# 1  pi=13'b1010011111100;
#1 $display("%b", po);
# 1  pi=13'b1010011111101;
#1 $display("%b", po);
# 1  pi=13'b1010011111110;
#1 $display("%b", po);
# 1  pi=13'b1010011111111;
#1 $display("%b", po);
# 1  pi=13'b1010100000000;
#1 $display("%b", po);
# 1  pi=13'b1010100000001;
#1 $display("%b", po);
# 1  pi=13'b1010100000010;
#1 $display("%b", po);
# 1  pi=13'b1010100000011;
#1 $display("%b", po);
# 1  pi=13'b1010100000100;
#1 $display("%b", po);
# 1  pi=13'b1010100000101;
#1 $display("%b", po);
# 1  pi=13'b1010100000110;
#1 $display("%b", po);
# 1  pi=13'b1010100000111;
#1 $display("%b", po);
# 1  pi=13'b1010100001000;
#1 $display("%b", po);
# 1  pi=13'b1010100001001;
#1 $display("%b", po);
# 1  pi=13'b1010100001010;
#1 $display("%b", po);
# 1  pi=13'b1010100001011;
#1 $display("%b", po);
# 1  pi=13'b1010100001100;
#1 $display("%b", po);
# 1  pi=13'b1010100001101;
#1 $display("%b", po);
# 1  pi=13'b1010100001110;
#1 $display("%b", po);
# 1  pi=13'b1010100001111;
#1 $display("%b", po);
# 1  pi=13'b1010100010000;
#1 $display("%b", po);
# 1  pi=13'b1010100010001;
#1 $display("%b", po);
# 1  pi=13'b1010100010010;
#1 $display("%b", po);
# 1  pi=13'b1010100010011;
#1 $display("%b", po);
# 1  pi=13'b1010100010100;
#1 $display("%b", po);
# 1  pi=13'b1010100010101;
#1 $display("%b", po);
# 1  pi=13'b1010100010110;
#1 $display("%b", po);
# 1  pi=13'b1010100010111;
#1 $display("%b", po);
# 1  pi=13'b1010100011000;
#1 $display("%b", po);
# 1  pi=13'b1010100011001;
#1 $display("%b", po);
# 1  pi=13'b1010100011010;
#1 $display("%b", po);
# 1  pi=13'b1010100011011;
#1 $display("%b", po);
# 1  pi=13'b1010100011100;
#1 $display("%b", po);
# 1  pi=13'b1010100011101;
#1 $display("%b", po);
# 1  pi=13'b1010100011110;
#1 $display("%b", po);
# 1  pi=13'b1010100011111;
#1 $display("%b", po);
# 1  pi=13'b1010100100000;
#1 $display("%b", po);
# 1  pi=13'b1010100100001;
#1 $display("%b", po);
# 1  pi=13'b1010100100010;
#1 $display("%b", po);
# 1  pi=13'b1010100100011;
#1 $display("%b", po);
# 1  pi=13'b1010100100100;
#1 $display("%b", po);
# 1  pi=13'b1010100100101;
#1 $display("%b", po);
# 1  pi=13'b1010100100110;
#1 $display("%b", po);
# 1  pi=13'b1010100100111;
#1 $display("%b", po);
# 1  pi=13'b1010100101000;
#1 $display("%b", po);
# 1  pi=13'b1010100101001;
#1 $display("%b", po);
# 1  pi=13'b1010100101010;
#1 $display("%b", po);
# 1  pi=13'b1010100101011;
#1 $display("%b", po);
# 1  pi=13'b1010100101100;
#1 $display("%b", po);
# 1  pi=13'b1010100101101;
#1 $display("%b", po);
# 1  pi=13'b1010100101110;
#1 $display("%b", po);
# 1  pi=13'b1010100101111;
#1 $display("%b", po);
# 1  pi=13'b1010100110000;
#1 $display("%b", po);
# 1  pi=13'b1010100110001;
#1 $display("%b", po);
# 1  pi=13'b1010100110010;
#1 $display("%b", po);
# 1  pi=13'b1010100110011;
#1 $display("%b", po);
# 1  pi=13'b1010100110100;
#1 $display("%b", po);
# 1  pi=13'b1010100110101;
#1 $display("%b", po);
# 1  pi=13'b1010100110110;
#1 $display("%b", po);
# 1  pi=13'b1010100110111;
#1 $display("%b", po);
# 1  pi=13'b1010100111000;
#1 $display("%b", po);
# 1  pi=13'b1010100111001;
#1 $display("%b", po);
# 1  pi=13'b1010100111010;
#1 $display("%b", po);
# 1  pi=13'b1010100111011;
#1 $display("%b", po);
# 1  pi=13'b1010100111100;
#1 $display("%b", po);
# 1  pi=13'b1010100111101;
#1 $display("%b", po);
# 1  pi=13'b1010100111110;
#1 $display("%b", po);
# 1  pi=13'b1010100111111;
#1 $display("%b", po);
# 1  pi=13'b1010101000000;
#1 $display("%b", po);
# 1  pi=13'b1010101000001;
#1 $display("%b", po);
# 1  pi=13'b1010101000010;
#1 $display("%b", po);
# 1  pi=13'b1010101000011;
#1 $display("%b", po);
# 1  pi=13'b1010101000100;
#1 $display("%b", po);
# 1  pi=13'b1010101000101;
#1 $display("%b", po);
# 1  pi=13'b1010101000110;
#1 $display("%b", po);
# 1  pi=13'b1010101000111;
#1 $display("%b", po);
# 1  pi=13'b1010101001000;
#1 $display("%b", po);
# 1  pi=13'b1010101001001;
#1 $display("%b", po);
# 1  pi=13'b1010101001010;
#1 $display("%b", po);
# 1  pi=13'b1010101001011;
#1 $display("%b", po);
# 1  pi=13'b1010101001100;
#1 $display("%b", po);
# 1  pi=13'b1010101001101;
#1 $display("%b", po);
# 1  pi=13'b1010101001110;
#1 $display("%b", po);
# 1  pi=13'b1010101001111;
#1 $display("%b", po);
# 1  pi=13'b1010101010000;
#1 $display("%b", po);
# 1  pi=13'b1010101010001;
#1 $display("%b", po);
# 1  pi=13'b1010101010010;
#1 $display("%b", po);
# 1  pi=13'b1010101010011;
#1 $display("%b", po);
# 1  pi=13'b1010101010100;
#1 $display("%b", po);
# 1  pi=13'b1010101010101;
#1 $display("%b", po);
# 1  pi=13'b1010101010110;
#1 $display("%b", po);
# 1  pi=13'b1010101010111;
#1 $display("%b", po);
# 1  pi=13'b1010101011000;
#1 $display("%b", po);
# 1  pi=13'b1010101011001;
#1 $display("%b", po);
# 1  pi=13'b1010101011010;
#1 $display("%b", po);
# 1  pi=13'b1010101011011;
#1 $display("%b", po);
# 1  pi=13'b1010101011100;
#1 $display("%b", po);
# 1  pi=13'b1010101011101;
#1 $display("%b", po);
# 1  pi=13'b1010101011110;
#1 $display("%b", po);
# 1  pi=13'b1010101011111;
#1 $display("%b", po);
# 1  pi=13'b1010101100000;
#1 $display("%b", po);
# 1  pi=13'b1010101100001;
#1 $display("%b", po);
# 1  pi=13'b1010101100010;
#1 $display("%b", po);
# 1  pi=13'b1010101100011;
#1 $display("%b", po);
# 1  pi=13'b1010101100100;
#1 $display("%b", po);
# 1  pi=13'b1010101100101;
#1 $display("%b", po);
# 1  pi=13'b1010101100110;
#1 $display("%b", po);
# 1  pi=13'b1010101100111;
#1 $display("%b", po);
# 1  pi=13'b1010101101000;
#1 $display("%b", po);
# 1  pi=13'b1010101101001;
#1 $display("%b", po);
# 1  pi=13'b1010101101010;
#1 $display("%b", po);
# 1  pi=13'b1010101101011;
#1 $display("%b", po);
# 1  pi=13'b1010101101100;
#1 $display("%b", po);
# 1  pi=13'b1010101101101;
#1 $display("%b", po);
# 1  pi=13'b1010101101110;
#1 $display("%b", po);
# 1  pi=13'b1010101101111;
#1 $display("%b", po);
# 1  pi=13'b1010101110000;
#1 $display("%b", po);
# 1  pi=13'b1010101110001;
#1 $display("%b", po);
# 1  pi=13'b1010101110010;
#1 $display("%b", po);
# 1  pi=13'b1010101110011;
#1 $display("%b", po);
# 1  pi=13'b1010101110100;
#1 $display("%b", po);
# 1  pi=13'b1010101110101;
#1 $display("%b", po);
# 1  pi=13'b1010101110110;
#1 $display("%b", po);
# 1  pi=13'b1010101110111;
#1 $display("%b", po);
# 1  pi=13'b1010101111000;
#1 $display("%b", po);
# 1  pi=13'b1010101111001;
#1 $display("%b", po);
# 1  pi=13'b1010101111010;
#1 $display("%b", po);
# 1  pi=13'b1010101111011;
#1 $display("%b", po);
# 1  pi=13'b1010101111100;
#1 $display("%b", po);
# 1  pi=13'b1010101111101;
#1 $display("%b", po);
# 1  pi=13'b1010101111110;
#1 $display("%b", po);
# 1  pi=13'b1010101111111;
#1 $display("%b", po);
# 1  pi=13'b1010110000000;
#1 $display("%b", po);
# 1  pi=13'b1010110000001;
#1 $display("%b", po);
# 1  pi=13'b1010110000010;
#1 $display("%b", po);
# 1  pi=13'b1010110000011;
#1 $display("%b", po);
# 1  pi=13'b1010110000100;
#1 $display("%b", po);
# 1  pi=13'b1010110000101;
#1 $display("%b", po);
# 1  pi=13'b1010110000110;
#1 $display("%b", po);
# 1  pi=13'b1010110000111;
#1 $display("%b", po);
# 1  pi=13'b1010110001000;
#1 $display("%b", po);
# 1  pi=13'b1010110001001;
#1 $display("%b", po);
# 1  pi=13'b1010110001010;
#1 $display("%b", po);
# 1  pi=13'b1010110001011;
#1 $display("%b", po);
# 1  pi=13'b1010110001100;
#1 $display("%b", po);
# 1  pi=13'b1010110001101;
#1 $display("%b", po);
# 1  pi=13'b1010110001110;
#1 $display("%b", po);
# 1  pi=13'b1010110001111;
#1 $display("%b", po);
# 1  pi=13'b1010110010000;
#1 $display("%b", po);
# 1  pi=13'b1010110010001;
#1 $display("%b", po);
# 1  pi=13'b1010110010010;
#1 $display("%b", po);
# 1  pi=13'b1010110010011;
#1 $display("%b", po);
# 1  pi=13'b1010110010100;
#1 $display("%b", po);
# 1  pi=13'b1010110010101;
#1 $display("%b", po);
# 1  pi=13'b1010110010110;
#1 $display("%b", po);
# 1  pi=13'b1010110010111;
#1 $display("%b", po);
# 1  pi=13'b1010110011000;
#1 $display("%b", po);
# 1  pi=13'b1010110011001;
#1 $display("%b", po);
# 1  pi=13'b1010110011010;
#1 $display("%b", po);
# 1  pi=13'b1010110011011;
#1 $display("%b", po);
# 1  pi=13'b1010110011100;
#1 $display("%b", po);
# 1  pi=13'b1010110011101;
#1 $display("%b", po);
# 1  pi=13'b1010110011110;
#1 $display("%b", po);
# 1  pi=13'b1010110011111;
#1 $display("%b", po);
# 1  pi=13'b1010110100000;
#1 $display("%b", po);
# 1  pi=13'b1010110100001;
#1 $display("%b", po);
# 1  pi=13'b1010110100010;
#1 $display("%b", po);
# 1  pi=13'b1010110100011;
#1 $display("%b", po);
# 1  pi=13'b1010110100100;
#1 $display("%b", po);
# 1  pi=13'b1010110100101;
#1 $display("%b", po);
# 1  pi=13'b1010110100110;
#1 $display("%b", po);
# 1  pi=13'b1010110100111;
#1 $display("%b", po);
# 1  pi=13'b1010110101000;
#1 $display("%b", po);
# 1  pi=13'b1010110101001;
#1 $display("%b", po);
# 1  pi=13'b1010110101010;
#1 $display("%b", po);
# 1  pi=13'b1010110101011;
#1 $display("%b", po);
# 1  pi=13'b1010110101100;
#1 $display("%b", po);
# 1  pi=13'b1010110101101;
#1 $display("%b", po);
# 1  pi=13'b1010110101110;
#1 $display("%b", po);
# 1  pi=13'b1010110101111;
#1 $display("%b", po);
# 1  pi=13'b1010110110000;
#1 $display("%b", po);
# 1  pi=13'b1010110110001;
#1 $display("%b", po);
# 1  pi=13'b1010110110010;
#1 $display("%b", po);
# 1  pi=13'b1010110110011;
#1 $display("%b", po);
# 1  pi=13'b1010110110100;
#1 $display("%b", po);
# 1  pi=13'b1010110110101;
#1 $display("%b", po);
# 1  pi=13'b1010110110110;
#1 $display("%b", po);
# 1  pi=13'b1010110110111;
#1 $display("%b", po);
# 1  pi=13'b1010110111000;
#1 $display("%b", po);
# 1  pi=13'b1010110111001;
#1 $display("%b", po);
# 1  pi=13'b1010110111010;
#1 $display("%b", po);
# 1  pi=13'b1010110111011;
#1 $display("%b", po);
# 1  pi=13'b1010110111100;
#1 $display("%b", po);
# 1  pi=13'b1010110111101;
#1 $display("%b", po);
# 1  pi=13'b1010110111110;
#1 $display("%b", po);
# 1  pi=13'b1010110111111;
#1 $display("%b", po);
# 1  pi=13'b1010111000000;
#1 $display("%b", po);
# 1  pi=13'b1010111000001;
#1 $display("%b", po);
# 1  pi=13'b1010111000010;
#1 $display("%b", po);
# 1  pi=13'b1010111000011;
#1 $display("%b", po);
# 1  pi=13'b1010111000100;
#1 $display("%b", po);
# 1  pi=13'b1010111000101;
#1 $display("%b", po);
# 1  pi=13'b1010111000110;
#1 $display("%b", po);
# 1  pi=13'b1010111000111;
#1 $display("%b", po);
# 1  pi=13'b1010111001000;
#1 $display("%b", po);
# 1  pi=13'b1010111001001;
#1 $display("%b", po);
# 1  pi=13'b1010111001010;
#1 $display("%b", po);
# 1  pi=13'b1010111001011;
#1 $display("%b", po);
# 1  pi=13'b1010111001100;
#1 $display("%b", po);
# 1  pi=13'b1010111001101;
#1 $display("%b", po);
# 1  pi=13'b1010111001110;
#1 $display("%b", po);
# 1  pi=13'b1010111001111;
#1 $display("%b", po);
# 1  pi=13'b1010111010000;
#1 $display("%b", po);
# 1  pi=13'b1010111010001;
#1 $display("%b", po);
# 1  pi=13'b1010111010010;
#1 $display("%b", po);
# 1  pi=13'b1010111010011;
#1 $display("%b", po);
# 1  pi=13'b1010111010100;
#1 $display("%b", po);
# 1  pi=13'b1010111010101;
#1 $display("%b", po);
# 1  pi=13'b1010111010110;
#1 $display("%b", po);
# 1  pi=13'b1010111010111;
#1 $display("%b", po);
# 1  pi=13'b1010111011000;
#1 $display("%b", po);
# 1  pi=13'b1010111011001;
#1 $display("%b", po);
# 1  pi=13'b1010111011010;
#1 $display("%b", po);
# 1  pi=13'b1010111011011;
#1 $display("%b", po);
# 1  pi=13'b1010111011100;
#1 $display("%b", po);
# 1  pi=13'b1010111011101;
#1 $display("%b", po);
# 1  pi=13'b1010111011110;
#1 $display("%b", po);
# 1  pi=13'b1010111011111;
#1 $display("%b", po);
# 1  pi=13'b1010111100000;
#1 $display("%b", po);
# 1  pi=13'b1010111100001;
#1 $display("%b", po);
# 1  pi=13'b1010111100010;
#1 $display("%b", po);
# 1  pi=13'b1010111100011;
#1 $display("%b", po);
# 1  pi=13'b1010111100100;
#1 $display("%b", po);
# 1  pi=13'b1010111100101;
#1 $display("%b", po);
# 1  pi=13'b1010111100110;
#1 $display("%b", po);
# 1  pi=13'b1010111100111;
#1 $display("%b", po);
# 1  pi=13'b1010111101000;
#1 $display("%b", po);
# 1  pi=13'b1010111101001;
#1 $display("%b", po);
# 1  pi=13'b1010111101010;
#1 $display("%b", po);
# 1  pi=13'b1010111101011;
#1 $display("%b", po);
# 1  pi=13'b1010111101100;
#1 $display("%b", po);
# 1  pi=13'b1010111101101;
#1 $display("%b", po);
# 1  pi=13'b1010111101110;
#1 $display("%b", po);
# 1  pi=13'b1010111101111;
#1 $display("%b", po);
# 1  pi=13'b1010111110000;
#1 $display("%b", po);
# 1  pi=13'b1010111110001;
#1 $display("%b", po);
# 1  pi=13'b1010111110010;
#1 $display("%b", po);
# 1  pi=13'b1010111110011;
#1 $display("%b", po);
# 1  pi=13'b1010111110100;
#1 $display("%b", po);
# 1  pi=13'b1010111110101;
#1 $display("%b", po);
# 1  pi=13'b1010111110110;
#1 $display("%b", po);
# 1  pi=13'b1010111110111;
#1 $display("%b", po);
# 1  pi=13'b1010111111000;
#1 $display("%b", po);
# 1  pi=13'b1010111111001;
#1 $display("%b", po);
# 1  pi=13'b1010111111010;
#1 $display("%b", po);
# 1  pi=13'b1010111111011;
#1 $display("%b", po);
# 1  pi=13'b1010111111100;
#1 $display("%b", po);
# 1  pi=13'b1010111111101;
#1 $display("%b", po);
# 1  pi=13'b1010111111110;
#1 $display("%b", po);
# 1  pi=13'b1010111111111;
#1 $display("%b", po);
# 1  pi=13'b1011000000000;
#1 $display("%b", po);
# 1  pi=13'b1011000000001;
#1 $display("%b", po);
# 1  pi=13'b1011000000010;
#1 $display("%b", po);
# 1  pi=13'b1011000000011;
#1 $display("%b", po);
# 1  pi=13'b1011000000100;
#1 $display("%b", po);
# 1  pi=13'b1011000000101;
#1 $display("%b", po);
# 1  pi=13'b1011000000110;
#1 $display("%b", po);
# 1  pi=13'b1011000000111;
#1 $display("%b", po);
# 1  pi=13'b1011000001000;
#1 $display("%b", po);
# 1  pi=13'b1011000001001;
#1 $display("%b", po);
# 1  pi=13'b1011000001010;
#1 $display("%b", po);
# 1  pi=13'b1011000001011;
#1 $display("%b", po);
# 1  pi=13'b1011000001100;
#1 $display("%b", po);
# 1  pi=13'b1011000001101;
#1 $display("%b", po);
# 1  pi=13'b1011000001110;
#1 $display("%b", po);
# 1  pi=13'b1011000001111;
#1 $display("%b", po);
# 1  pi=13'b1011000010000;
#1 $display("%b", po);
# 1  pi=13'b1011000010001;
#1 $display("%b", po);
# 1  pi=13'b1011000010010;
#1 $display("%b", po);
# 1  pi=13'b1011000010011;
#1 $display("%b", po);
# 1  pi=13'b1011000010100;
#1 $display("%b", po);
# 1  pi=13'b1011000010101;
#1 $display("%b", po);
# 1  pi=13'b1011000010110;
#1 $display("%b", po);
# 1  pi=13'b1011000010111;
#1 $display("%b", po);
# 1  pi=13'b1011000011000;
#1 $display("%b", po);
# 1  pi=13'b1011000011001;
#1 $display("%b", po);
# 1  pi=13'b1011000011010;
#1 $display("%b", po);
# 1  pi=13'b1011000011011;
#1 $display("%b", po);
# 1  pi=13'b1011000011100;
#1 $display("%b", po);
# 1  pi=13'b1011000011101;
#1 $display("%b", po);
# 1  pi=13'b1011000011110;
#1 $display("%b", po);
# 1  pi=13'b1011000011111;
#1 $display("%b", po);
# 1  pi=13'b1011000100000;
#1 $display("%b", po);
# 1  pi=13'b1011000100001;
#1 $display("%b", po);
# 1  pi=13'b1011000100010;
#1 $display("%b", po);
# 1  pi=13'b1011000100011;
#1 $display("%b", po);
# 1  pi=13'b1011000100100;
#1 $display("%b", po);
# 1  pi=13'b1011000100101;
#1 $display("%b", po);
# 1  pi=13'b1011000100110;
#1 $display("%b", po);
# 1  pi=13'b1011000100111;
#1 $display("%b", po);
# 1  pi=13'b1011000101000;
#1 $display("%b", po);
# 1  pi=13'b1011000101001;
#1 $display("%b", po);
# 1  pi=13'b1011000101010;
#1 $display("%b", po);
# 1  pi=13'b1011000101011;
#1 $display("%b", po);
# 1  pi=13'b1011000101100;
#1 $display("%b", po);
# 1  pi=13'b1011000101101;
#1 $display("%b", po);
# 1  pi=13'b1011000101110;
#1 $display("%b", po);
# 1  pi=13'b1011000101111;
#1 $display("%b", po);
# 1  pi=13'b1011000110000;
#1 $display("%b", po);
# 1  pi=13'b1011000110001;
#1 $display("%b", po);
# 1  pi=13'b1011000110010;
#1 $display("%b", po);
# 1  pi=13'b1011000110011;
#1 $display("%b", po);
# 1  pi=13'b1011000110100;
#1 $display("%b", po);
# 1  pi=13'b1011000110101;
#1 $display("%b", po);
# 1  pi=13'b1011000110110;
#1 $display("%b", po);
# 1  pi=13'b1011000110111;
#1 $display("%b", po);
# 1  pi=13'b1011000111000;
#1 $display("%b", po);
# 1  pi=13'b1011000111001;
#1 $display("%b", po);
# 1  pi=13'b1011000111010;
#1 $display("%b", po);
# 1  pi=13'b1011000111011;
#1 $display("%b", po);
# 1  pi=13'b1011000111100;
#1 $display("%b", po);
# 1  pi=13'b1011000111101;
#1 $display("%b", po);
# 1  pi=13'b1011000111110;
#1 $display("%b", po);
# 1  pi=13'b1011000111111;
#1 $display("%b", po);
# 1  pi=13'b1011001000000;
#1 $display("%b", po);
# 1  pi=13'b1011001000001;
#1 $display("%b", po);
# 1  pi=13'b1011001000010;
#1 $display("%b", po);
# 1  pi=13'b1011001000011;
#1 $display("%b", po);
# 1  pi=13'b1011001000100;
#1 $display("%b", po);
# 1  pi=13'b1011001000101;
#1 $display("%b", po);
# 1  pi=13'b1011001000110;
#1 $display("%b", po);
# 1  pi=13'b1011001000111;
#1 $display("%b", po);
# 1  pi=13'b1011001001000;
#1 $display("%b", po);
# 1  pi=13'b1011001001001;
#1 $display("%b", po);
# 1  pi=13'b1011001001010;
#1 $display("%b", po);
# 1  pi=13'b1011001001011;
#1 $display("%b", po);
# 1  pi=13'b1011001001100;
#1 $display("%b", po);
# 1  pi=13'b1011001001101;
#1 $display("%b", po);
# 1  pi=13'b1011001001110;
#1 $display("%b", po);
# 1  pi=13'b1011001001111;
#1 $display("%b", po);
# 1  pi=13'b1011001010000;
#1 $display("%b", po);
# 1  pi=13'b1011001010001;
#1 $display("%b", po);
# 1  pi=13'b1011001010010;
#1 $display("%b", po);
# 1  pi=13'b1011001010011;
#1 $display("%b", po);
# 1  pi=13'b1011001010100;
#1 $display("%b", po);
# 1  pi=13'b1011001010101;
#1 $display("%b", po);
# 1  pi=13'b1011001010110;
#1 $display("%b", po);
# 1  pi=13'b1011001010111;
#1 $display("%b", po);
# 1  pi=13'b1011001011000;
#1 $display("%b", po);
# 1  pi=13'b1011001011001;
#1 $display("%b", po);
# 1  pi=13'b1011001011010;
#1 $display("%b", po);
# 1  pi=13'b1011001011011;
#1 $display("%b", po);
# 1  pi=13'b1011001011100;
#1 $display("%b", po);
# 1  pi=13'b1011001011101;
#1 $display("%b", po);
# 1  pi=13'b1011001011110;
#1 $display("%b", po);
# 1  pi=13'b1011001011111;
#1 $display("%b", po);
# 1  pi=13'b1011001100000;
#1 $display("%b", po);
# 1  pi=13'b1011001100001;
#1 $display("%b", po);
# 1  pi=13'b1011001100010;
#1 $display("%b", po);
# 1  pi=13'b1011001100011;
#1 $display("%b", po);
# 1  pi=13'b1011001100100;
#1 $display("%b", po);
# 1  pi=13'b1011001100101;
#1 $display("%b", po);
# 1  pi=13'b1011001100110;
#1 $display("%b", po);
# 1  pi=13'b1011001100111;
#1 $display("%b", po);
# 1  pi=13'b1011001101000;
#1 $display("%b", po);
# 1  pi=13'b1011001101001;
#1 $display("%b", po);
# 1  pi=13'b1011001101010;
#1 $display("%b", po);
# 1  pi=13'b1011001101011;
#1 $display("%b", po);
# 1  pi=13'b1011001101100;
#1 $display("%b", po);
# 1  pi=13'b1011001101101;
#1 $display("%b", po);
# 1  pi=13'b1011001101110;
#1 $display("%b", po);
# 1  pi=13'b1011001101111;
#1 $display("%b", po);
# 1  pi=13'b1011001110000;
#1 $display("%b", po);
# 1  pi=13'b1011001110001;
#1 $display("%b", po);
# 1  pi=13'b1011001110010;
#1 $display("%b", po);
# 1  pi=13'b1011001110011;
#1 $display("%b", po);
# 1  pi=13'b1011001110100;
#1 $display("%b", po);
# 1  pi=13'b1011001110101;
#1 $display("%b", po);
# 1  pi=13'b1011001110110;
#1 $display("%b", po);
# 1  pi=13'b1011001110111;
#1 $display("%b", po);
# 1  pi=13'b1011001111000;
#1 $display("%b", po);
# 1  pi=13'b1011001111001;
#1 $display("%b", po);
# 1  pi=13'b1011001111010;
#1 $display("%b", po);
# 1  pi=13'b1011001111011;
#1 $display("%b", po);
# 1  pi=13'b1011001111100;
#1 $display("%b", po);
# 1  pi=13'b1011001111101;
#1 $display("%b", po);
# 1  pi=13'b1011001111110;
#1 $display("%b", po);
# 1  pi=13'b1011001111111;
#1 $display("%b", po);
# 1  pi=13'b1011010000000;
#1 $display("%b", po);
# 1  pi=13'b1011010000001;
#1 $display("%b", po);
# 1  pi=13'b1011010000010;
#1 $display("%b", po);
# 1  pi=13'b1011010000011;
#1 $display("%b", po);
# 1  pi=13'b1011010000100;
#1 $display("%b", po);
# 1  pi=13'b1011010000101;
#1 $display("%b", po);
# 1  pi=13'b1011010000110;
#1 $display("%b", po);
# 1  pi=13'b1011010000111;
#1 $display("%b", po);
# 1  pi=13'b1011010001000;
#1 $display("%b", po);
# 1  pi=13'b1011010001001;
#1 $display("%b", po);
# 1  pi=13'b1011010001010;
#1 $display("%b", po);
# 1  pi=13'b1011010001011;
#1 $display("%b", po);
# 1  pi=13'b1011010001100;
#1 $display("%b", po);
# 1  pi=13'b1011010001101;
#1 $display("%b", po);
# 1  pi=13'b1011010001110;
#1 $display("%b", po);
# 1  pi=13'b1011010001111;
#1 $display("%b", po);
# 1  pi=13'b1011010010000;
#1 $display("%b", po);
# 1  pi=13'b1011010010001;
#1 $display("%b", po);
# 1  pi=13'b1011010010010;
#1 $display("%b", po);
# 1  pi=13'b1011010010011;
#1 $display("%b", po);
# 1  pi=13'b1011010010100;
#1 $display("%b", po);
# 1  pi=13'b1011010010101;
#1 $display("%b", po);
# 1  pi=13'b1011010010110;
#1 $display("%b", po);
# 1  pi=13'b1011010010111;
#1 $display("%b", po);
# 1  pi=13'b1011010011000;
#1 $display("%b", po);
# 1  pi=13'b1011010011001;
#1 $display("%b", po);
# 1  pi=13'b1011010011010;
#1 $display("%b", po);
# 1  pi=13'b1011010011011;
#1 $display("%b", po);
# 1  pi=13'b1011010011100;
#1 $display("%b", po);
# 1  pi=13'b1011010011101;
#1 $display("%b", po);
# 1  pi=13'b1011010011110;
#1 $display("%b", po);
# 1  pi=13'b1011010011111;
#1 $display("%b", po);
# 1  pi=13'b1011010100000;
#1 $display("%b", po);
# 1  pi=13'b1011010100001;
#1 $display("%b", po);
# 1  pi=13'b1011010100010;
#1 $display("%b", po);
# 1  pi=13'b1011010100011;
#1 $display("%b", po);
# 1  pi=13'b1011010100100;
#1 $display("%b", po);
# 1  pi=13'b1011010100101;
#1 $display("%b", po);
# 1  pi=13'b1011010100110;
#1 $display("%b", po);
# 1  pi=13'b1011010100111;
#1 $display("%b", po);
# 1  pi=13'b1011010101000;
#1 $display("%b", po);
# 1  pi=13'b1011010101001;
#1 $display("%b", po);
# 1  pi=13'b1011010101010;
#1 $display("%b", po);
# 1  pi=13'b1011010101011;
#1 $display("%b", po);
# 1  pi=13'b1011010101100;
#1 $display("%b", po);
# 1  pi=13'b1011010101101;
#1 $display("%b", po);
# 1  pi=13'b1011010101110;
#1 $display("%b", po);
# 1  pi=13'b1011010101111;
#1 $display("%b", po);
# 1  pi=13'b1011010110000;
#1 $display("%b", po);
# 1  pi=13'b1011010110001;
#1 $display("%b", po);
# 1  pi=13'b1011010110010;
#1 $display("%b", po);
# 1  pi=13'b1011010110011;
#1 $display("%b", po);
# 1  pi=13'b1011010110100;
#1 $display("%b", po);
# 1  pi=13'b1011010110101;
#1 $display("%b", po);
# 1  pi=13'b1011010110110;
#1 $display("%b", po);
# 1  pi=13'b1011010110111;
#1 $display("%b", po);
# 1  pi=13'b1011010111000;
#1 $display("%b", po);
# 1  pi=13'b1011010111001;
#1 $display("%b", po);
# 1  pi=13'b1011010111010;
#1 $display("%b", po);
# 1  pi=13'b1011010111011;
#1 $display("%b", po);
# 1  pi=13'b1011010111100;
#1 $display("%b", po);
# 1  pi=13'b1011010111101;
#1 $display("%b", po);
# 1  pi=13'b1011010111110;
#1 $display("%b", po);
# 1  pi=13'b1011010111111;
#1 $display("%b", po);
# 1  pi=13'b1011011000000;
#1 $display("%b", po);
# 1  pi=13'b1011011000001;
#1 $display("%b", po);
# 1  pi=13'b1011011000010;
#1 $display("%b", po);
# 1  pi=13'b1011011000011;
#1 $display("%b", po);
# 1  pi=13'b1011011000100;
#1 $display("%b", po);
# 1  pi=13'b1011011000101;
#1 $display("%b", po);
# 1  pi=13'b1011011000110;
#1 $display("%b", po);
# 1  pi=13'b1011011000111;
#1 $display("%b", po);
# 1  pi=13'b1011011001000;
#1 $display("%b", po);
# 1  pi=13'b1011011001001;
#1 $display("%b", po);
# 1  pi=13'b1011011001010;
#1 $display("%b", po);
# 1  pi=13'b1011011001011;
#1 $display("%b", po);
# 1  pi=13'b1011011001100;
#1 $display("%b", po);
# 1  pi=13'b1011011001101;
#1 $display("%b", po);
# 1  pi=13'b1011011001110;
#1 $display("%b", po);
# 1  pi=13'b1011011001111;
#1 $display("%b", po);
# 1  pi=13'b1011011010000;
#1 $display("%b", po);
# 1  pi=13'b1011011010001;
#1 $display("%b", po);
# 1  pi=13'b1011011010010;
#1 $display("%b", po);
# 1  pi=13'b1011011010011;
#1 $display("%b", po);
# 1  pi=13'b1011011010100;
#1 $display("%b", po);
# 1  pi=13'b1011011010101;
#1 $display("%b", po);
# 1  pi=13'b1011011010110;
#1 $display("%b", po);
# 1  pi=13'b1011011010111;
#1 $display("%b", po);
# 1  pi=13'b1011011011000;
#1 $display("%b", po);
# 1  pi=13'b1011011011001;
#1 $display("%b", po);
# 1  pi=13'b1011011011010;
#1 $display("%b", po);
# 1  pi=13'b1011011011011;
#1 $display("%b", po);
# 1  pi=13'b1011011011100;
#1 $display("%b", po);
# 1  pi=13'b1011011011101;
#1 $display("%b", po);
# 1  pi=13'b1011011011110;
#1 $display("%b", po);
# 1  pi=13'b1011011011111;
#1 $display("%b", po);
# 1  pi=13'b1011011100000;
#1 $display("%b", po);
# 1  pi=13'b1011011100001;
#1 $display("%b", po);
# 1  pi=13'b1011011100010;
#1 $display("%b", po);
# 1  pi=13'b1011011100011;
#1 $display("%b", po);
# 1  pi=13'b1011011100100;
#1 $display("%b", po);
# 1  pi=13'b1011011100101;
#1 $display("%b", po);
# 1  pi=13'b1011011100110;
#1 $display("%b", po);
# 1  pi=13'b1011011100111;
#1 $display("%b", po);
# 1  pi=13'b1011011101000;
#1 $display("%b", po);
# 1  pi=13'b1011011101001;
#1 $display("%b", po);
# 1  pi=13'b1011011101010;
#1 $display("%b", po);
# 1  pi=13'b1011011101011;
#1 $display("%b", po);
# 1  pi=13'b1011011101100;
#1 $display("%b", po);
# 1  pi=13'b1011011101101;
#1 $display("%b", po);
# 1  pi=13'b1011011101110;
#1 $display("%b", po);
# 1  pi=13'b1011011101111;
#1 $display("%b", po);
# 1  pi=13'b1011011110000;
#1 $display("%b", po);
# 1  pi=13'b1011011110001;
#1 $display("%b", po);
# 1  pi=13'b1011011110010;
#1 $display("%b", po);
# 1  pi=13'b1011011110011;
#1 $display("%b", po);
# 1  pi=13'b1011011110100;
#1 $display("%b", po);
# 1  pi=13'b1011011110101;
#1 $display("%b", po);
# 1  pi=13'b1011011110110;
#1 $display("%b", po);
# 1  pi=13'b1011011110111;
#1 $display("%b", po);
# 1  pi=13'b1011011111000;
#1 $display("%b", po);
# 1  pi=13'b1011011111001;
#1 $display("%b", po);
# 1  pi=13'b1011011111010;
#1 $display("%b", po);
# 1  pi=13'b1011011111011;
#1 $display("%b", po);
# 1  pi=13'b1011011111100;
#1 $display("%b", po);
# 1  pi=13'b1011011111101;
#1 $display("%b", po);
# 1  pi=13'b1011011111110;
#1 $display("%b", po);
# 1  pi=13'b1011011111111;
#1 $display("%b", po);
# 1  pi=13'b1011100000000;
#1 $display("%b", po);
# 1  pi=13'b1011100000001;
#1 $display("%b", po);
# 1  pi=13'b1011100000010;
#1 $display("%b", po);
# 1  pi=13'b1011100000011;
#1 $display("%b", po);
# 1  pi=13'b1011100000100;
#1 $display("%b", po);
# 1  pi=13'b1011100000101;
#1 $display("%b", po);
# 1  pi=13'b1011100000110;
#1 $display("%b", po);
# 1  pi=13'b1011100000111;
#1 $display("%b", po);
# 1  pi=13'b1011100001000;
#1 $display("%b", po);
# 1  pi=13'b1011100001001;
#1 $display("%b", po);
# 1  pi=13'b1011100001010;
#1 $display("%b", po);
# 1  pi=13'b1011100001011;
#1 $display("%b", po);
# 1  pi=13'b1011100001100;
#1 $display("%b", po);
# 1  pi=13'b1011100001101;
#1 $display("%b", po);
# 1  pi=13'b1011100001110;
#1 $display("%b", po);
# 1  pi=13'b1011100001111;
#1 $display("%b", po);
# 1  pi=13'b1011100010000;
#1 $display("%b", po);
# 1  pi=13'b1011100010001;
#1 $display("%b", po);
# 1  pi=13'b1011100010010;
#1 $display("%b", po);
# 1  pi=13'b1011100010011;
#1 $display("%b", po);
# 1  pi=13'b1011100010100;
#1 $display("%b", po);
# 1  pi=13'b1011100010101;
#1 $display("%b", po);
# 1  pi=13'b1011100010110;
#1 $display("%b", po);
# 1  pi=13'b1011100010111;
#1 $display("%b", po);
# 1  pi=13'b1011100011000;
#1 $display("%b", po);
# 1  pi=13'b1011100011001;
#1 $display("%b", po);
# 1  pi=13'b1011100011010;
#1 $display("%b", po);
# 1  pi=13'b1011100011011;
#1 $display("%b", po);
# 1  pi=13'b1011100011100;
#1 $display("%b", po);
# 1  pi=13'b1011100011101;
#1 $display("%b", po);
# 1  pi=13'b1011100011110;
#1 $display("%b", po);
# 1  pi=13'b1011100011111;
#1 $display("%b", po);
# 1  pi=13'b1011100100000;
#1 $display("%b", po);
# 1  pi=13'b1011100100001;
#1 $display("%b", po);
# 1  pi=13'b1011100100010;
#1 $display("%b", po);
# 1  pi=13'b1011100100011;
#1 $display("%b", po);
# 1  pi=13'b1011100100100;
#1 $display("%b", po);
# 1  pi=13'b1011100100101;
#1 $display("%b", po);
# 1  pi=13'b1011100100110;
#1 $display("%b", po);
# 1  pi=13'b1011100100111;
#1 $display("%b", po);
# 1  pi=13'b1011100101000;
#1 $display("%b", po);
# 1  pi=13'b1011100101001;
#1 $display("%b", po);
# 1  pi=13'b1011100101010;
#1 $display("%b", po);
# 1  pi=13'b1011100101011;
#1 $display("%b", po);
# 1  pi=13'b1011100101100;
#1 $display("%b", po);
# 1  pi=13'b1011100101101;
#1 $display("%b", po);
# 1  pi=13'b1011100101110;
#1 $display("%b", po);
# 1  pi=13'b1011100101111;
#1 $display("%b", po);
# 1  pi=13'b1011100110000;
#1 $display("%b", po);
# 1  pi=13'b1011100110001;
#1 $display("%b", po);
# 1  pi=13'b1011100110010;
#1 $display("%b", po);
# 1  pi=13'b1011100110011;
#1 $display("%b", po);
# 1  pi=13'b1011100110100;
#1 $display("%b", po);
# 1  pi=13'b1011100110101;
#1 $display("%b", po);
# 1  pi=13'b1011100110110;
#1 $display("%b", po);
# 1  pi=13'b1011100110111;
#1 $display("%b", po);
# 1  pi=13'b1011100111000;
#1 $display("%b", po);
# 1  pi=13'b1011100111001;
#1 $display("%b", po);
# 1  pi=13'b1011100111010;
#1 $display("%b", po);
# 1  pi=13'b1011100111011;
#1 $display("%b", po);
# 1  pi=13'b1011100111100;
#1 $display("%b", po);
# 1  pi=13'b1011100111101;
#1 $display("%b", po);
# 1  pi=13'b1011100111110;
#1 $display("%b", po);
# 1  pi=13'b1011100111111;
#1 $display("%b", po);
# 1  pi=13'b1011101000000;
#1 $display("%b", po);
# 1  pi=13'b1011101000001;
#1 $display("%b", po);
# 1  pi=13'b1011101000010;
#1 $display("%b", po);
# 1  pi=13'b1011101000011;
#1 $display("%b", po);
# 1  pi=13'b1011101000100;
#1 $display("%b", po);
# 1  pi=13'b1011101000101;
#1 $display("%b", po);
# 1  pi=13'b1011101000110;
#1 $display("%b", po);
# 1  pi=13'b1011101000111;
#1 $display("%b", po);
# 1  pi=13'b1011101001000;
#1 $display("%b", po);
# 1  pi=13'b1011101001001;
#1 $display("%b", po);
# 1  pi=13'b1011101001010;
#1 $display("%b", po);
# 1  pi=13'b1011101001011;
#1 $display("%b", po);
# 1  pi=13'b1011101001100;
#1 $display("%b", po);
# 1  pi=13'b1011101001101;
#1 $display("%b", po);
# 1  pi=13'b1011101001110;
#1 $display("%b", po);
# 1  pi=13'b1011101001111;
#1 $display("%b", po);
# 1  pi=13'b1011101010000;
#1 $display("%b", po);
# 1  pi=13'b1011101010001;
#1 $display("%b", po);
# 1  pi=13'b1011101010010;
#1 $display("%b", po);
# 1  pi=13'b1011101010011;
#1 $display("%b", po);
# 1  pi=13'b1011101010100;
#1 $display("%b", po);
# 1  pi=13'b1011101010101;
#1 $display("%b", po);
# 1  pi=13'b1011101010110;
#1 $display("%b", po);
# 1  pi=13'b1011101010111;
#1 $display("%b", po);
# 1  pi=13'b1011101011000;
#1 $display("%b", po);
# 1  pi=13'b1011101011001;
#1 $display("%b", po);
# 1  pi=13'b1011101011010;
#1 $display("%b", po);
# 1  pi=13'b1011101011011;
#1 $display("%b", po);
# 1  pi=13'b1011101011100;
#1 $display("%b", po);
# 1  pi=13'b1011101011101;
#1 $display("%b", po);
# 1  pi=13'b1011101011110;
#1 $display("%b", po);
# 1  pi=13'b1011101011111;
#1 $display("%b", po);
# 1  pi=13'b1011101100000;
#1 $display("%b", po);
# 1  pi=13'b1011101100001;
#1 $display("%b", po);
# 1  pi=13'b1011101100010;
#1 $display("%b", po);
# 1  pi=13'b1011101100011;
#1 $display("%b", po);
# 1  pi=13'b1011101100100;
#1 $display("%b", po);
# 1  pi=13'b1011101100101;
#1 $display("%b", po);
# 1  pi=13'b1011101100110;
#1 $display("%b", po);
# 1  pi=13'b1011101100111;
#1 $display("%b", po);
# 1  pi=13'b1011101101000;
#1 $display("%b", po);
# 1  pi=13'b1011101101001;
#1 $display("%b", po);
# 1  pi=13'b1011101101010;
#1 $display("%b", po);
# 1  pi=13'b1011101101011;
#1 $display("%b", po);
# 1  pi=13'b1011101101100;
#1 $display("%b", po);
# 1  pi=13'b1011101101101;
#1 $display("%b", po);
# 1  pi=13'b1011101101110;
#1 $display("%b", po);
# 1  pi=13'b1011101101111;
#1 $display("%b", po);
# 1  pi=13'b1011101110000;
#1 $display("%b", po);
# 1  pi=13'b1011101110001;
#1 $display("%b", po);
# 1  pi=13'b1011101110010;
#1 $display("%b", po);
# 1  pi=13'b1011101110011;
#1 $display("%b", po);
# 1  pi=13'b1011101110100;
#1 $display("%b", po);
# 1  pi=13'b1011101110101;
#1 $display("%b", po);
# 1  pi=13'b1011101110110;
#1 $display("%b", po);
# 1  pi=13'b1011101110111;
#1 $display("%b", po);
# 1  pi=13'b1011101111000;
#1 $display("%b", po);
# 1  pi=13'b1011101111001;
#1 $display("%b", po);
# 1  pi=13'b1011101111010;
#1 $display("%b", po);
# 1  pi=13'b1011101111011;
#1 $display("%b", po);
# 1  pi=13'b1011101111100;
#1 $display("%b", po);
# 1  pi=13'b1011101111101;
#1 $display("%b", po);
# 1  pi=13'b1011101111110;
#1 $display("%b", po);
# 1  pi=13'b1011101111111;
#1 $display("%b", po);
# 1  pi=13'b1011110000000;
#1 $display("%b", po);
# 1  pi=13'b1011110000001;
#1 $display("%b", po);
# 1  pi=13'b1011110000010;
#1 $display("%b", po);
# 1  pi=13'b1011110000011;
#1 $display("%b", po);
# 1  pi=13'b1011110000100;
#1 $display("%b", po);
# 1  pi=13'b1011110000101;
#1 $display("%b", po);
# 1  pi=13'b1011110000110;
#1 $display("%b", po);
# 1  pi=13'b1011110000111;
#1 $display("%b", po);
# 1  pi=13'b1011110001000;
#1 $display("%b", po);
# 1  pi=13'b1011110001001;
#1 $display("%b", po);
# 1  pi=13'b1011110001010;
#1 $display("%b", po);
# 1  pi=13'b1011110001011;
#1 $display("%b", po);
# 1  pi=13'b1011110001100;
#1 $display("%b", po);
# 1  pi=13'b1011110001101;
#1 $display("%b", po);
# 1  pi=13'b1011110001110;
#1 $display("%b", po);
# 1  pi=13'b1011110001111;
#1 $display("%b", po);
# 1  pi=13'b1011110010000;
#1 $display("%b", po);
# 1  pi=13'b1011110010001;
#1 $display("%b", po);
# 1  pi=13'b1011110010010;
#1 $display("%b", po);
# 1  pi=13'b1011110010011;
#1 $display("%b", po);
# 1  pi=13'b1011110010100;
#1 $display("%b", po);
# 1  pi=13'b1011110010101;
#1 $display("%b", po);
# 1  pi=13'b1011110010110;
#1 $display("%b", po);
# 1  pi=13'b1011110010111;
#1 $display("%b", po);
# 1  pi=13'b1011110011000;
#1 $display("%b", po);
# 1  pi=13'b1011110011001;
#1 $display("%b", po);
# 1  pi=13'b1011110011010;
#1 $display("%b", po);
# 1  pi=13'b1011110011011;
#1 $display("%b", po);
# 1  pi=13'b1011110011100;
#1 $display("%b", po);
# 1  pi=13'b1011110011101;
#1 $display("%b", po);
# 1  pi=13'b1011110011110;
#1 $display("%b", po);
# 1  pi=13'b1011110011111;
#1 $display("%b", po);
# 1  pi=13'b1011110100000;
#1 $display("%b", po);
# 1  pi=13'b1011110100001;
#1 $display("%b", po);
# 1  pi=13'b1011110100010;
#1 $display("%b", po);
# 1  pi=13'b1011110100011;
#1 $display("%b", po);
# 1  pi=13'b1011110100100;
#1 $display("%b", po);
# 1  pi=13'b1011110100101;
#1 $display("%b", po);
# 1  pi=13'b1011110100110;
#1 $display("%b", po);
# 1  pi=13'b1011110100111;
#1 $display("%b", po);
# 1  pi=13'b1011110101000;
#1 $display("%b", po);
# 1  pi=13'b1011110101001;
#1 $display("%b", po);
# 1  pi=13'b1011110101010;
#1 $display("%b", po);
# 1  pi=13'b1011110101011;
#1 $display("%b", po);
# 1  pi=13'b1011110101100;
#1 $display("%b", po);
# 1  pi=13'b1011110101101;
#1 $display("%b", po);
# 1  pi=13'b1011110101110;
#1 $display("%b", po);
# 1  pi=13'b1011110101111;
#1 $display("%b", po);
# 1  pi=13'b1011110110000;
#1 $display("%b", po);
# 1  pi=13'b1011110110001;
#1 $display("%b", po);
# 1  pi=13'b1011110110010;
#1 $display("%b", po);
# 1  pi=13'b1011110110011;
#1 $display("%b", po);
# 1  pi=13'b1011110110100;
#1 $display("%b", po);
# 1  pi=13'b1011110110101;
#1 $display("%b", po);
# 1  pi=13'b1011110110110;
#1 $display("%b", po);
# 1  pi=13'b1011110110111;
#1 $display("%b", po);
# 1  pi=13'b1011110111000;
#1 $display("%b", po);
# 1  pi=13'b1011110111001;
#1 $display("%b", po);
# 1  pi=13'b1011110111010;
#1 $display("%b", po);
# 1  pi=13'b1011110111011;
#1 $display("%b", po);
# 1  pi=13'b1011110111100;
#1 $display("%b", po);
# 1  pi=13'b1011110111101;
#1 $display("%b", po);
# 1  pi=13'b1011110111110;
#1 $display("%b", po);
# 1  pi=13'b1011110111111;
#1 $display("%b", po);
# 1  pi=13'b1011111000000;
#1 $display("%b", po);
# 1  pi=13'b1011111000001;
#1 $display("%b", po);
# 1  pi=13'b1011111000010;
#1 $display("%b", po);
# 1  pi=13'b1011111000011;
#1 $display("%b", po);
# 1  pi=13'b1011111000100;
#1 $display("%b", po);
# 1  pi=13'b1011111000101;
#1 $display("%b", po);
# 1  pi=13'b1011111000110;
#1 $display("%b", po);
# 1  pi=13'b1011111000111;
#1 $display("%b", po);
# 1  pi=13'b1011111001000;
#1 $display("%b", po);
# 1  pi=13'b1011111001001;
#1 $display("%b", po);
# 1  pi=13'b1011111001010;
#1 $display("%b", po);
# 1  pi=13'b1011111001011;
#1 $display("%b", po);
# 1  pi=13'b1011111001100;
#1 $display("%b", po);
# 1  pi=13'b1011111001101;
#1 $display("%b", po);
# 1  pi=13'b1011111001110;
#1 $display("%b", po);
# 1  pi=13'b1011111001111;
#1 $display("%b", po);
# 1  pi=13'b1011111010000;
#1 $display("%b", po);
# 1  pi=13'b1011111010001;
#1 $display("%b", po);
# 1  pi=13'b1011111010010;
#1 $display("%b", po);
# 1  pi=13'b1011111010011;
#1 $display("%b", po);
# 1  pi=13'b1011111010100;
#1 $display("%b", po);
# 1  pi=13'b1011111010101;
#1 $display("%b", po);
# 1  pi=13'b1011111010110;
#1 $display("%b", po);
# 1  pi=13'b1011111010111;
#1 $display("%b", po);
# 1  pi=13'b1011111011000;
#1 $display("%b", po);
# 1  pi=13'b1011111011001;
#1 $display("%b", po);
# 1  pi=13'b1011111011010;
#1 $display("%b", po);
# 1  pi=13'b1011111011011;
#1 $display("%b", po);
# 1  pi=13'b1011111011100;
#1 $display("%b", po);
# 1  pi=13'b1011111011101;
#1 $display("%b", po);
# 1  pi=13'b1011111011110;
#1 $display("%b", po);
# 1  pi=13'b1011111011111;
#1 $display("%b", po);
# 1  pi=13'b1011111100000;
#1 $display("%b", po);
# 1  pi=13'b1011111100001;
#1 $display("%b", po);
# 1  pi=13'b1011111100010;
#1 $display("%b", po);
# 1  pi=13'b1011111100011;
#1 $display("%b", po);
# 1  pi=13'b1011111100100;
#1 $display("%b", po);
# 1  pi=13'b1011111100101;
#1 $display("%b", po);
# 1  pi=13'b1011111100110;
#1 $display("%b", po);
# 1  pi=13'b1011111100111;
#1 $display("%b", po);
# 1  pi=13'b1011111101000;
#1 $display("%b", po);
# 1  pi=13'b1011111101001;
#1 $display("%b", po);
# 1  pi=13'b1011111101010;
#1 $display("%b", po);
# 1  pi=13'b1011111101011;
#1 $display("%b", po);
# 1  pi=13'b1011111101100;
#1 $display("%b", po);
# 1  pi=13'b1011111101101;
#1 $display("%b", po);
# 1  pi=13'b1011111101110;
#1 $display("%b", po);
# 1  pi=13'b1011111101111;
#1 $display("%b", po);
# 1  pi=13'b1011111110000;
#1 $display("%b", po);
# 1  pi=13'b1011111110001;
#1 $display("%b", po);
# 1  pi=13'b1011111110010;
#1 $display("%b", po);
# 1  pi=13'b1011111110011;
#1 $display("%b", po);
# 1  pi=13'b1011111110100;
#1 $display("%b", po);
# 1  pi=13'b1011111110101;
#1 $display("%b", po);
# 1  pi=13'b1011111110110;
#1 $display("%b", po);
# 1  pi=13'b1011111110111;
#1 $display("%b", po);
# 1  pi=13'b1011111111000;
#1 $display("%b", po);
# 1  pi=13'b1011111111001;
#1 $display("%b", po);
# 1  pi=13'b1011111111010;
#1 $display("%b", po);
# 1  pi=13'b1011111111011;
#1 $display("%b", po);
# 1  pi=13'b1011111111100;
#1 $display("%b", po);
# 1  pi=13'b1011111111101;
#1 $display("%b", po);
# 1  pi=13'b1011111111110;
#1 $display("%b", po);
# 1  pi=13'b1011111111111;
#1 $display("%b", po);
# 1  pi=13'b1100000000000;
#1 $display("%b", po);
# 1  pi=13'b1100000000001;
#1 $display("%b", po);
# 1  pi=13'b1100000000010;
#1 $display("%b", po);
# 1  pi=13'b1100000000011;
#1 $display("%b", po);
# 1  pi=13'b1100000000100;
#1 $display("%b", po);
# 1  pi=13'b1100000000101;
#1 $display("%b", po);
# 1  pi=13'b1100000000110;
#1 $display("%b", po);
# 1  pi=13'b1100000000111;
#1 $display("%b", po);
# 1  pi=13'b1100000001000;
#1 $display("%b", po);
# 1  pi=13'b1100000001001;
#1 $display("%b", po);
# 1  pi=13'b1100000001010;
#1 $display("%b", po);
# 1  pi=13'b1100000001011;
#1 $display("%b", po);
# 1  pi=13'b1100000001100;
#1 $display("%b", po);
# 1  pi=13'b1100000001101;
#1 $display("%b", po);
# 1  pi=13'b1100000001110;
#1 $display("%b", po);
# 1  pi=13'b1100000001111;
#1 $display("%b", po);
# 1  pi=13'b1100000010000;
#1 $display("%b", po);
# 1  pi=13'b1100000010001;
#1 $display("%b", po);
# 1  pi=13'b1100000010010;
#1 $display("%b", po);
# 1  pi=13'b1100000010011;
#1 $display("%b", po);
# 1  pi=13'b1100000010100;
#1 $display("%b", po);
# 1  pi=13'b1100000010101;
#1 $display("%b", po);
# 1  pi=13'b1100000010110;
#1 $display("%b", po);
# 1  pi=13'b1100000010111;
#1 $display("%b", po);
# 1  pi=13'b1100000011000;
#1 $display("%b", po);
# 1  pi=13'b1100000011001;
#1 $display("%b", po);
# 1  pi=13'b1100000011010;
#1 $display("%b", po);
# 1  pi=13'b1100000011011;
#1 $display("%b", po);
# 1  pi=13'b1100000011100;
#1 $display("%b", po);
# 1  pi=13'b1100000011101;
#1 $display("%b", po);
# 1  pi=13'b1100000011110;
#1 $display("%b", po);
# 1  pi=13'b1100000011111;
#1 $display("%b", po);
# 1  pi=13'b1100000100000;
#1 $display("%b", po);
# 1  pi=13'b1100000100001;
#1 $display("%b", po);
# 1  pi=13'b1100000100010;
#1 $display("%b", po);
# 1  pi=13'b1100000100011;
#1 $display("%b", po);
# 1  pi=13'b1100000100100;
#1 $display("%b", po);
# 1  pi=13'b1100000100101;
#1 $display("%b", po);
# 1  pi=13'b1100000100110;
#1 $display("%b", po);
# 1  pi=13'b1100000100111;
#1 $display("%b", po);
# 1  pi=13'b1100000101000;
#1 $display("%b", po);
# 1  pi=13'b1100000101001;
#1 $display("%b", po);
# 1  pi=13'b1100000101010;
#1 $display("%b", po);
# 1  pi=13'b1100000101011;
#1 $display("%b", po);
# 1  pi=13'b1100000101100;
#1 $display("%b", po);
# 1  pi=13'b1100000101101;
#1 $display("%b", po);
# 1  pi=13'b1100000101110;
#1 $display("%b", po);
# 1  pi=13'b1100000101111;
#1 $display("%b", po);
# 1  pi=13'b1100000110000;
#1 $display("%b", po);
# 1  pi=13'b1100000110001;
#1 $display("%b", po);
# 1  pi=13'b1100000110010;
#1 $display("%b", po);
# 1  pi=13'b1100000110011;
#1 $display("%b", po);
# 1  pi=13'b1100000110100;
#1 $display("%b", po);
# 1  pi=13'b1100000110101;
#1 $display("%b", po);
# 1  pi=13'b1100000110110;
#1 $display("%b", po);
# 1  pi=13'b1100000110111;
#1 $display("%b", po);
# 1  pi=13'b1100000111000;
#1 $display("%b", po);
# 1  pi=13'b1100000111001;
#1 $display("%b", po);
# 1  pi=13'b1100000111010;
#1 $display("%b", po);
# 1  pi=13'b1100000111011;
#1 $display("%b", po);
# 1  pi=13'b1100000111100;
#1 $display("%b", po);
# 1  pi=13'b1100000111101;
#1 $display("%b", po);
# 1  pi=13'b1100000111110;
#1 $display("%b", po);
# 1  pi=13'b1100000111111;
#1 $display("%b", po);
# 1  pi=13'b1100001000000;
#1 $display("%b", po);
# 1  pi=13'b1100001000001;
#1 $display("%b", po);
# 1  pi=13'b1100001000010;
#1 $display("%b", po);
# 1  pi=13'b1100001000011;
#1 $display("%b", po);
# 1  pi=13'b1100001000100;
#1 $display("%b", po);
# 1  pi=13'b1100001000101;
#1 $display("%b", po);
# 1  pi=13'b1100001000110;
#1 $display("%b", po);
# 1  pi=13'b1100001000111;
#1 $display("%b", po);
# 1  pi=13'b1100001001000;
#1 $display("%b", po);
# 1  pi=13'b1100001001001;
#1 $display("%b", po);
# 1  pi=13'b1100001001010;
#1 $display("%b", po);
# 1  pi=13'b1100001001011;
#1 $display("%b", po);
# 1  pi=13'b1100001001100;
#1 $display("%b", po);
# 1  pi=13'b1100001001101;
#1 $display("%b", po);
# 1  pi=13'b1100001001110;
#1 $display("%b", po);
# 1  pi=13'b1100001001111;
#1 $display("%b", po);
# 1  pi=13'b1100001010000;
#1 $display("%b", po);
# 1  pi=13'b1100001010001;
#1 $display("%b", po);
# 1  pi=13'b1100001010010;
#1 $display("%b", po);
# 1  pi=13'b1100001010011;
#1 $display("%b", po);
# 1  pi=13'b1100001010100;
#1 $display("%b", po);
# 1  pi=13'b1100001010101;
#1 $display("%b", po);
# 1  pi=13'b1100001010110;
#1 $display("%b", po);
# 1  pi=13'b1100001010111;
#1 $display("%b", po);
# 1  pi=13'b1100001011000;
#1 $display("%b", po);
# 1  pi=13'b1100001011001;
#1 $display("%b", po);
# 1  pi=13'b1100001011010;
#1 $display("%b", po);
# 1  pi=13'b1100001011011;
#1 $display("%b", po);
# 1  pi=13'b1100001011100;
#1 $display("%b", po);
# 1  pi=13'b1100001011101;
#1 $display("%b", po);
# 1  pi=13'b1100001011110;
#1 $display("%b", po);
# 1  pi=13'b1100001011111;
#1 $display("%b", po);
# 1  pi=13'b1100001100000;
#1 $display("%b", po);
# 1  pi=13'b1100001100001;
#1 $display("%b", po);
# 1  pi=13'b1100001100010;
#1 $display("%b", po);
# 1  pi=13'b1100001100011;
#1 $display("%b", po);
# 1  pi=13'b1100001100100;
#1 $display("%b", po);
# 1  pi=13'b1100001100101;
#1 $display("%b", po);
# 1  pi=13'b1100001100110;
#1 $display("%b", po);
# 1  pi=13'b1100001100111;
#1 $display("%b", po);
# 1  pi=13'b1100001101000;
#1 $display("%b", po);
# 1  pi=13'b1100001101001;
#1 $display("%b", po);
# 1  pi=13'b1100001101010;
#1 $display("%b", po);
# 1  pi=13'b1100001101011;
#1 $display("%b", po);
# 1  pi=13'b1100001101100;
#1 $display("%b", po);
# 1  pi=13'b1100001101101;
#1 $display("%b", po);
# 1  pi=13'b1100001101110;
#1 $display("%b", po);
# 1  pi=13'b1100001101111;
#1 $display("%b", po);
# 1  pi=13'b1100001110000;
#1 $display("%b", po);
# 1  pi=13'b1100001110001;
#1 $display("%b", po);
# 1  pi=13'b1100001110010;
#1 $display("%b", po);
# 1  pi=13'b1100001110011;
#1 $display("%b", po);
# 1  pi=13'b1100001110100;
#1 $display("%b", po);
# 1  pi=13'b1100001110101;
#1 $display("%b", po);
# 1  pi=13'b1100001110110;
#1 $display("%b", po);
# 1  pi=13'b1100001110111;
#1 $display("%b", po);
# 1  pi=13'b1100001111000;
#1 $display("%b", po);
# 1  pi=13'b1100001111001;
#1 $display("%b", po);
# 1  pi=13'b1100001111010;
#1 $display("%b", po);
# 1  pi=13'b1100001111011;
#1 $display("%b", po);
# 1  pi=13'b1100001111100;
#1 $display("%b", po);
# 1  pi=13'b1100001111101;
#1 $display("%b", po);
# 1  pi=13'b1100001111110;
#1 $display("%b", po);
# 1  pi=13'b1100001111111;
#1 $display("%b", po);
# 1  pi=13'b1100010000000;
#1 $display("%b", po);
# 1  pi=13'b1100010000001;
#1 $display("%b", po);
# 1  pi=13'b1100010000010;
#1 $display("%b", po);
# 1  pi=13'b1100010000011;
#1 $display("%b", po);
# 1  pi=13'b1100010000100;
#1 $display("%b", po);
# 1  pi=13'b1100010000101;
#1 $display("%b", po);
# 1  pi=13'b1100010000110;
#1 $display("%b", po);
# 1  pi=13'b1100010000111;
#1 $display("%b", po);
# 1  pi=13'b1100010001000;
#1 $display("%b", po);
# 1  pi=13'b1100010001001;
#1 $display("%b", po);
# 1  pi=13'b1100010001010;
#1 $display("%b", po);
# 1  pi=13'b1100010001011;
#1 $display("%b", po);
# 1  pi=13'b1100010001100;
#1 $display("%b", po);
# 1  pi=13'b1100010001101;
#1 $display("%b", po);
# 1  pi=13'b1100010001110;
#1 $display("%b", po);
# 1  pi=13'b1100010001111;
#1 $display("%b", po);
# 1  pi=13'b1100010010000;
#1 $display("%b", po);
# 1  pi=13'b1100010010001;
#1 $display("%b", po);
# 1  pi=13'b1100010010010;
#1 $display("%b", po);
# 1  pi=13'b1100010010011;
#1 $display("%b", po);
# 1  pi=13'b1100010010100;
#1 $display("%b", po);
# 1  pi=13'b1100010010101;
#1 $display("%b", po);
# 1  pi=13'b1100010010110;
#1 $display("%b", po);
# 1  pi=13'b1100010010111;
#1 $display("%b", po);
# 1  pi=13'b1100010011000;
#1 $display("%b", po);
# 1  pi=13'b1100010011001;
#1 $display("%b", po);
# 1  pi=13'b1100010011010;
#1 $display("%b", po);
# 1  pi=13'b1100010011011;
#1 $display("%b", po);
# 1  pi=13'b1100010011100;
#1 $display("%b", po);
# 1  pi=13'b1100010011101;
#1 $display("%b", po);
# 1  pi=13'b1100010011110;
#1 $display("%b", po);
# 1  pi=13'b1100010011111;
#1 $display("%b", po);
# 1  pi=13'b1100010100000;
#1 $display("%b", po);
# 1  pi=13'b1100010100001;
#1 $display("%b", po);
# 1  pi=13'b1100010100010;
#1 $display("%b", po);
# 1  pi=13'b1100010100011;
#1 $display("%b", po);
# 1  pi=13'b1100010100100;
#1 $display("%b", po);
# 1  pi=13'b1100010100101;
#1 $display("%b", po);
# 1  pi=13'b1100010100110;
#1 $display("%b", po);
# 1  pi=13'b1100010100111;
#1 $display("%b", po);
# 1  pi=13'b1100010101000;
#1 $display("%b", po);
# 1  pi=13'b1100010101001;
#1 $display("%b", po);
# 1  pi=13'b1100010101010;
#1 $display("%b", po);
# 1  pi=13'b1100010101011;
#1 $display("%b", po);
# 1  pi=13'b1100010101100;
#1 $display("%b", po);
# 1  pi=13'b1100010101101;
#1 $display("%b", po);
# 1  pi=13'b1100010101110;
#1 $display("%b", po);
# 1  pi=13'b1100010101111;
#1 $display("%b", po);
# 1  pi=13'b1100010110000;
#1 $display("%b", po);
# 1  pi=13'b1100010110001;
#1 $display("%b", po);
# 1  pi=13'b1100010110010;
#1 $display("%b", po);
# 1  pi=13'b1100010110011;
#1 $display("%b", po);
# 1  pi=13'b1100010110100;
#1 $display("%b", po);
# 1  pi=13'b1100010110101;
#1 $display("%b", po);
# 1  pi=13'b1100010110110;
#1 $display("%b", po);
# 1  pi=13'b1100010110111;
#1 $display("%b", po);
# 1  pi=13'b1100010111000;
#1 $display("%b", po);
# 1  pi=13'b1100010111001;
#1 $display("%b", po);
# 1  pi=13'b1100010111010;
#1 $display("%b", po);
# 1  pi=13'b1100010111011;
#1 $display("%b", po);
# 1  pi=13'b1100010111100;
#1 $display("%b", po);
# 1  pi=13'b1100010111101;
#1 $display("%b", po);
# 1  pi=13'b1100010111110;
#1 $display("%b", po);
# 1  pi=13'b1100010111111;
#1 $display("%b", po);
# 1  pi=13'b1100011000000;
#1 $display("%b", po);
# 1  pi=13'b1100011000001;
#1 $display("%b", po);
# 1  pi=13'b1100011000010;
#1 $display("%b", po);
# 1  pi=13'b1100011000011;
#1 $display("%b", po);
# 1  pi=13'b1100011000100;
#1 $display("%b", po);
# 1  pi=13'b1100011000101;
#1 $display("%b", po);
# 1  pi=13'b1100011000110;
#1 $display("%b", po);
# 1  pi=13'b1100011000111;
#1 $display("%b", po);
# 1  pi=13'b1100011001000;
#1 $display("%b", po);
# 1  pi=13'b1100011001001;
#1 $display("%b", po);
# 1  pi=13'b1100011001010;
#1 $display("%b", po);
# 1  pi=13'b1100011001011;
#1 $display("%b", po);
# 1  pi=13'b1100011001100;
#1 $display("%b", po);
# 1  pi=13'b1100011001101;
#1 $display("%b", po);
# 1  pi=13'b1100011001110;
#1 $display("%b", po);
# 1  pi=13'b1100011001111;
#1 $display("%b", po);
# 1  pi=13'b1100011010000;
#1 $display("%b", po);
# 1  pi=13'b1100011010001;
#1 $display("%b", po);
# 1  pi=13'b1100011010010;
#1 $display("%b", po);
# 1  pi=13'b1100011010011;
#1 $display("%b", po);
# 1  pi=13'b1100011010100;
#1 $display("%b", po);
# 1  pi=13'b1100011010101;
#1 $display("%b", po);
# 1  pi=13'b1100011010110;
#1 $display("%b", po);
# 1  pi=13'b1100011010111;
#1 $display("%b", po);
# 1  pi=13'b1100011011000;
#1 $display("%b", po);
# 1  pi=13'b1100011011001;
#1 $display("%b", po);
# 1  pi=13'b1100011011010;
#1 $display("%b", po);
# 1  pi=13'b1100011011011;
#1 $display("%b", po);
# 1  pi=13'b1100011011100;
#1 $display("%b", po);
# 1  pi=13'b1100011011101;
#1 $display("%b", po);
# 1  pi=13'b1100011011110;
#1 $display("%b", po);
# 1  pi=13'b1100011011111;
#1 $display("%b", po);
# 1  pi=13'b1100011100000;
#1 $display("%b", po);
# 1  pi=13'b1100011100001;
#1 $display("%b", po);
# 1  pi=13'b1100011100010;
#1 $display("%b", po);
# 1  pi=13'b1100011100011;
#1 $display("%b", po);
# 1  pi=13'b1100011100100;
#1 $display("%b", po);
# 1  pi=13'b1100011100101;
#1 $display("%b", po);
# 1  pi=13'b1100011100110;
#1 $display("%b", po);
# 1  pi=13'b1100011100111;
#1 $display("%b", po);
# 1  pi=13'b1100011101000;
#1 $display("%b", po);
# 1  pi=13'b1100011101001;
#1 $display("%b", po);
# 1  pi=13'b1100011101010;
#1 $display("%b", po);
# 1  pi=13'b1100011101011;
#1 $display("%b", po);
# 1  pi=13'b1100011101100;
#1 $display("%b", po);
# 1  pi=13'b1100011101101;
#1 $display("%b", po);
# 1  pi=13'b1100011101110;
#1 $display("%b", po);
# 1  pi=13'b1100011101111;
#1 $display("%b", po);
# 1  pi=13'b1100011110000;
#1 $display("%b", po);
# 1  pi=13'b1100011110001;
#1 $display("%b", po);
# 1  pi=13'b1100011110010;
#1 $display("%b", po);
# 1  pi=13'b1100011110011;
#1 $display("%b", po);
# 1  pi=13'b1100011110100;
#1 $display("%b", po);
# 1  pi=13'b1100011110101;
#1 $display("%b", po);
# 1  pi=13'b1100011110110;
#1 $display("%b", po);
# 1  pi=13'b1100011110111;
#1 $display("%b", po);
# 1  pi=13'b1100011111000;
#1 $display("%b", po);
# 1  pi=13'b1100011111001;
#1 $display("%b", po);
# 1  pi=13'b1100011111010;
#1 $display("%b", po);
# 1  pi=13'b1100011111011;
#1 $display("%b", po);
# 1  pi=13'b1100011111100;
#1 $display("%b", po);
# 1  pi=13'b1100011111101;
#1 $display("%b", po);
# 1  pi=13'b1100011111110;
#1 $display("%b", po);
# 1  pi=13'b1100011111111;
#1 $display("%b", po);
# 1  pi=13'b1100100000000;
#1 $display("%b", po);
# 1  pi=13'b1100100000001;
#1 $display("%b", po);
# 1  pi=13'b1100100000010;
#1 $display("%b", po);
# 1  pi=13'b1100100000011;
#1 $display("%b", po);
# 1  pi=13'b1100100000100;
#1 $display("%b", po);
# 1  pi=13'b1100100000101;
#1 $display("%b", po);
# 1  pi=13'b1100100000110;
#1 $display("%b", po);
# 1  pi=13'b1100100000111;
#1 $display("%b", po);
# 1  pi=13'b1100100001000;
#1 $display("%b", po);
# 1  pi=13'b1100100001001;
#1 $display("%b", po);
# 1  pi=13'b1100100001010;
#1 $display("%b", po);
# 1  pi=13'b1100100001011;
#1 $display("%b", po);
# 1  pi=13'b1100100001100;
#1 $display("%b", po);
# 1  pi=13'b1100100001101;
#1 $display("%b", po);
# 1  pi=13'b1100100001110;
#1 $display("%b", po);
# 1  pi=13'b1100100001111;
#1 $display("%b", po);
# 1  pi=13'b1100100010000;
#1 $display("%b", po);
# 1  pi=13'b1100100010001;
#1 $display("%b", po);
# 1  pi=13'b1100100010010;
#1 $display("%b", po);
# 1  pi=13'b1100100010011;
#1 $display("%b", po);
# 1  pi=13'b1100100010100;
#1 $display("%b", po);
# 1  pi=13'b1100100010101;
#1 $display("%b", po);
# 1  pi=13'b1100100010110;
#1 $display("%b", po);
# 1  pi=13'b1100100010111;
#1 $display("%b", po);
# 1  pi=13'b1100100011000;
#1 $display("%b", po);
# 1  pi=13'b1100100011001;
#1 $display("%b", po);
# 1  pi=13'b1100100011010;
#1 $display("%b", po);
# 1  pi=13'b1100100011011;
#1 $display("%b", po);
# 1  pi=13'b1100100011100;
#1 $display("%b", po);
# 1  pi=13'b1100100011101;
#1 $display("%b", po);
# 1  pi=13'b1100100011110;
#1 $display("%b", po);
# 1  pi=13'b1100100011111;
#1 $display("%b", po);
# 1  pi=13'b1100100100000;
#1 $display("%b", po);
# 1  pi=13'b1100100100001;
#1 $display("%b", po);
# 1  pi=13'b1100100100010;
#1 $display("%b", po);
# 1  pi=13'b1100100100011;
#1 $display("%b", po);
# 1  pi=13'b1100100100100;
#1 $display("%b", po);
# 1  pi=13'b1100100100101;
#1 $display("%b", po);
# 1  pi=13'b1100100100110;
#1 $display("%b", po);
# 1  pi=13'b1100100100111;
#1 $display("%b", po);
# 1  pi=13'b1100100101000;
#1 $display("%b", po);
# 1  pi=13'b1100100101001;
#1 $display("%b", po);
# 1  pi=13'b1100100101010;
#1 $display("%b", po);
# 1  pi=13'b1100100101011;
#1 $display("%b", po);
# 1  pi=13'b1100100101100;
#1 $display("%b", po);
# 1  pi=13'b1100100101101;
#1 $display("%b", po);
# 1  pi=13'b1100100101110;
#1 $display("%b", po);
# 1  pi=13'b1100100101111;
#1 $display("%b", po);
# 1  pi=13'b1100100110000;
#1 $display("%b", po);
# 1  pi=13'b1100100110001;
#1 $display("%b", po);
# 1  pi=13'b1100100110010;
#1 $display("%b", po);
# 1  pi=13'b1100100110011;
#1 $display("%b", po);
# 1  pi=13'b1100100110100;
#1 $display("%b", po);
# 1  pi=13'b1100100110101;
#1 $display("%b", po);
# 1  pi=13'b1100100110110;
#1 $display("%b", po);
# 1  pi=13'b1100100110111;
#1 $display("%b", po);
# 1  pi=13'b1100100111000;
#1 $display("%b", po);
# 1  pi=13'b1100100111001;
#1 $display("%b", po);
# 1  pi=13'b1100100111010;
#1 $display("%b", po);
# 1  pi=13'b1100100111011;
#1 $display("%b", po);
# 1  pi=13'b1100100111100;
#1 $display("%b", po);
# 1  pi=13'b1100100111101;
#1 $display("%b", po);
# 1  pi=13'b1100100111110;
#1 $display("%b", po);
# 1  pi=13'b1100100111111;
#1 $display("%b", po);
# 1  pi=13'b1100101000000;
#1 $display("%b", po);
# 1  pi=13'b1100101000001;
#1 $display("%b", po);
# 1  pi=13'b1100101000010;
#1 $display("%b", po);
# 1  pi=13'b1100101000011;
#1 $display("%b", po);
# 1  pi=13'b1100101000100;
#1 $display("%b", po);
# 1  pi=13'b1100101000101;
#1 $display("%b", po);
# 1  pi=13'b1100101000110;
#1 $display("%b", po);
# 1  pi=13'b1100101000111;
#1 $display("%b", po);
# 1  pi=13'b1100101001000;
#1 $display("%b", po);
# 1  pi=13'b1100101001001;
#1 $display("%b", po);
# 1  pi=13'b1100101001010;
#1 $display("%b", po);
# 1  pi=13'b1100101001011;
#1 $display("%b", po);
# 1  pi=13'b1100101001100;
#1 $display("%b", po);
# 1  pi=13'b1100101001101;
#1 $display("%b", po);
# 1  pi=13'b1100101001110;
#1 $display("%b", po);
# 1  pi=13'b1100101001111;
#1 $display("%b", po);
# 1  pi=13'b1100101010000;
#1 $display("%b", po);
# 1  pi=13'b1100101010001;
#1 $display("%b", po);
# 1  pi=13'b1100101010010;
#1 $display("%b", po);
# 1  pi=13'b1100101010011;
#1 $display("%b", po);
# 1  pi=13'b1100101010100;
#1 $display("%b", po);
# 1  pi=13'b1100101010101;
#1 $display("%b", po);
# 1  pi=13'b1100101010110;
#1 $display("%b", po);
# 1  pi=13'b1100101010111;
#1 $display("%b", po);
# 1  pi=13'b1100101011000;
#1 $display("%b", po);
# 1  pi=13'b1100101011001;
#1 $display("%b", po);
# 1  pi=13'b1100101011010;
#1 $display("%b", po);
# 1  pi=13'b1100101011011;
#1 $display("%b", po);
# 1  pi=13'b1100101011100;
#1 $display("%b", po);
# 1  pi=13'b1100101011101;
#1 $display("%b", po);
# 1  pi=13'b1100101011110;
#1 $display("%b", po);
# 1  pi=13'b1100101011111;
#1 $display("%b", po);
# 1  pi=13'b1100101100000;
#1 $display("%b", po);
# 1  pi=13'b1100101100001;
#1 $display("%b", po);
# 1  pi=13'b1100101100010;
#1 $display("%b", po);
# 1  pi=13'b1100101100011;
#1 $display("%b", po);
# 1  pi=13'b1100101100100;
#1 $display("%b", po);
# 1  pi=13'b1100101100101;
#1 $display("%b", po);
# 1  pi=13'b1100101100110;
#1 $display("%b", po);
# 1  pi=13'b1100101100111;
#1 $display("%b", po);
# 1  pi=13'b1100101101000;
#1 $display("%b", po);
# 1  pi=13'b1100101101001;
#1 $display("%b", po);
# 1  pi=13'b1100101101010;
#1 $display("%b", po);
# 1  pi=13'b1100101101011;
#1 $display("%b", po);
# 1  pi=13'b1100101101100;
#1 $display("%b", po);
# 1  pi=13'b1100101101101;
#1 $display("%b", po);
# 1  pi=13'b1100101101110;
#1 $display("%b", po);
# 1  pi=13'b1100101101111;
#1 $display("%b", po);
# 1  pi=13'b1100101110000;
#1 $display("%b", po);
# 1  pi=13'b1100101110001;
#1 $display("%b", po);
# 1  pi=13'b1100101110010;
#1 $display("%b", po);
# 1  pi=13'b1100101110011;
#1 $display("%b", po);
# 1  pi=13'b1100101110100;
#1 $display("%b", po);
# 1  pi=13'b1100101110101;
#1 $display("%b", po);
# 1  pi=13'b1100101110110;
#1 $display("%b", po);
# 1  pi=13'b1100101110111;
#1 $display("%b", po);
# 1  pi=13'b1100101111000;
#1 $display("%b", po);
# 1  pi=13'b1100101111001;
#1 $display("%b", po);
# 1  pi=13'b1100101111010;
#1 $display("%b", po);
# 1  pi=13'b1100101111011;
#1 $display("%b", po);
# 1  pi=13'b1100101111100;
#1 $display("%b", po);
# 1  pi=13'b1100101111101;
#1 $display("%b", po);
# 1  pi=13'b1100101111110;
#1 $display("%b", po);
# 1  pi=13'b1100101111111;
#1 $display("%b", po);
# 1  pi=13'b1100110000000;
#1 $display("%b", po);
# 1  pi=13'b1100110000001;
#1 $display("%b", po);
# 1  pi=13'b1100110000010;
#1 $display("%b", po);
# 1  pi=13'b1100110000011;
#1 $display("%b", po);
# 1  pi=13'b1100110000100;
#1 $display("%b", po);
# 1  pi=13'b1100110000101;
#1 $display("%b", po);
# 1  pi=13'b1100110000110;
#1 $display("%b", po);
# 1  pi=13'b1100110000111;
#1 $display("%b", po);
# 1  pi=13'b1100110001000;
#1 $display("%b", po);
# 1  pi=13'b1100110001001;
#1 $display("%b", po);
# 1  pi=13'b1100110001010;
#1 $display("%b", po);
# 1  pi=13'b1100110001011;
#1 $display("%b", po);
# 1  pi=13'b1100110001100;
#1 $display("%b", po);
# 1  pi=13'b1100110001101;
#1 $display("%b", po);
# 1  pi=13'b1100110001110;
#1 $display("%b", po);
# 1  pi=13'b1100110001111;
#1 $display("%b", po);
# 1  pi=13'b1100110010000;
#1 $display("%b", po);
# 1  pi=13'b1100110010001;
#1 $display("%b", po);
# 1  pi=13'b1100110010010;
#1 $display("%b", po);
# 1  pi=13'b1100110010011;
#1 $display("%b", po);
# 1  pi=13'b1100110010100;
#1 $display("%b", po);
# 1  pi=13'b1100110010101;
#1 $display("%b", po);
# 1  pi=13'b1100110010110;
#1 $display("%b", po);
# 1  pi=13'b1100110010111;
#1 $display("%b", po);
# 1  pi=13'b1100110011000;
#1 $display("%b", po);
# 1  pi=13'b1100110011001;
#1 $display("%b", po);
# 1  pi=13'b1100110011010;
#1 $display("%b", po);
# 1  pi=13'b1100110011011;
#1 $display("%b", po);
# 1  pi=13'b1100110011100;
#1 $display("%b", po);
# 1  pi=13'b1100110011101;
#1 $display("%b", po);
# 1  pi=13'b1100110011110;
#1 $display("%b", po);
# 1  pi=13'b1100110011111;
#1 $display("%b", po);
# 1  pi=13'b1100110100000;
#1 $display("%b", po);
# 1  pi=13'b1100110100001;
#1 $display("%b", po);
# 1  pi=13'b1100110100010;
#1 $display("%b", po);
# 1  pi=13'b1100110100011;
#1 $display("%b", po);
# 1  pi=13'b1100110100100;
#1 $display("%b", po);
# 1  pi=13'b1100110100101;
#1 $display("%b", po);
# 1  pi=13'b1100110100110;
#1 $display("%b", po);
# 1  pi=13'b1100110100111;
#1 $display("%b", po);
# 1  pi=13'b1100110101000;
#1 $display("%b", po);
# 1  pi=13'b1100110101001;
#1 $display("%b", po);
# 1  pi=13'b1100110101010;
#1 $display("%b", po);
# 1  pi=13'b1100110101011;
#1 $display("%b", po);
# 1  pi=13'b1100110101100;
#1 $display("%b", po);
# 1  pi=13'b1100110101101;
#1 $display("%b", po);
# 1  pi=13'b1100110101110;
#1 $display("%b", po);
# 1  pi=13'b1100110101111;
#1 $display("%b", po);
# 1  pi=13'b1100110110000;
#1 $display("%b", po);
# 1  pi=13'b1100110110001;
#1 $display("%b", po);
# 1  pi=13'b1100110110010;
#1 $display("%b", po);
# 1  pi=13'b1100110110011;
#1 $display("%b", po);
# 1  pi=13'b1100110110100;
#1 $display("%b", po);
# 1  pi=13'b1100110110101;
#1 $display("%b", po);
# 1  pi=13'b1100110110110;
#1 $display("%b", po);
# 1  pi=13'b1100110110111;
#1 $display("%b", po);
# 1  pi=13'b1100110111000;
#1 $display("%b", po);
# 1  pi=13'b1100110111001;
#1 $display("%b", po);
# 1  pi=13'b1100110111010;
#1 $display("%b", po);
# 1  pi=13'b1100110111011;
#1 $display("%b", po);
# 1  pi=13'b1100110111100;
#1 $display("%b", po);
# 1  pi=13'b1100110111101;
#1 $display("%b", po);
# 1  pi=13'b1100110111110;
#1 $display("%b", po);
# 1  pi=13'b1100110111111;
#1 $display("%b", po);
# 1  pi=13'b1100111000000;
#1 $display("%b", po);
# 1  pi=13'b1100111000001;
#1 $display("%b", po);
# 1  pi=13'b1100111000010;
#1 $display("%b", po);
# 1  pi=13'b1100111000011;
#1 $display("%b", po);
# 1  pi=13'b1100111000100;
#1 $display("%b", po);
# 1  pi=13'b1100111000101;
#1 $display("%b", po);
# 1  pi=13'b1100111000110;
#1 $display("%b", po);
# 1  pi=13'b1100111000111;
#1 $display("%b", po);
# 1  pi=13'b1100111001000;
#1 $display("%b", po);
# 1  pi=13'b1100111001001;
#1 $display("%b", po);
# 1  pi=13'b1100111001010;
#1 $display("%b", po);
# 1  pi=13'b1100111001011;
#1 $display("%b", po);
# 1  pi=13'b1100111001100;
#1 $display("%b", po);
# 1  pi=13'b1100111001101;
#1 $display("%b", po);
# 1  pi=13'b1100111001110;
#1 $display("%b", po);
# 1  pi=13'b1100111001111;
#1 $display("%b", po);
# 1  pi=13'b1100111010000;
#1 $display("%b", po);
# 1  pi=13'b1100111010001;
#1 $display("%b", po);
# 1  pi=13'b1100111010010;
#1 $display("%b", po);
# 1  pi=13'b1100111010011;
#1 $display("%b", po);
# 1  pi=13'b1100111010100;
#1 $display("%b", po);
# 1  pi=13'b1100111010101;
#1 $display("%b", po);
# 1  pi=13'b1100111010110;
#1 $display("%b", po);
# 1  pi=13'b1100111010111;
#1 $display("%b", po);
# 1  pi=13'b1100111011000;
#1 $display("%b", po);
# 1  pi=13'b1100111011001;
#1 $display("%b", po);
# 1  pi=13'b1100111011010;
#1 $display("%b", po);
# 1  pi=13'b1100111011011;
#1 $display("%b", po);
# 1  pi=13'b1100111011100;
#1 $display("%b", po);
# 1  pi=13'b1100111011101;
#1 $display("%b", po);
# 1  pi=13'b1100111011110;
#1 $display("%b", po);
# 1  pi=13'b1100111011111;
#1 $display("%b", po);
# 1  pi=13'b1100111100000;
#1 $display("%b", po);
# 1  pi=13'b1100111100001;
#1 $display("%b", po);
# 1  pi=13'b1100111100010;
#1 $display("%b", po);
# 1  pi=13'b1100111100011;
#1 $display("%b", po);
# 1  pi=13'b1100111100100;
#1 $display("%b", po);
# 1  pi=13'b1100111100101;
#1 $display("%b", po);
# 1  pi=13'b1100111100110;
#1 $display("%b", po);
# 1  pi=13'b1100111100111;
#1 $display("%b", po);
# 1  pi=13'b1100111101000;
#1 $display("%b", po);
# 1  pi=13'b1100111101001;
#1 $display("%b", po);
# 1  pi=13'b1100111101010;
#1 $display("%b", po);
# 1  pi=13'b1100111101011;
#1 $display("%b", po);
# 1  pi=13'b1100111101100;
#1 $display("%b", po);
# 1  pi=13'b1100111101101;
#1 $display("%b", po);
# 1  pi=13'b1100111101110;
#1 $display("%b", po);
# 1  pi=13'b1100111101111;
#1 $display("%b", po);
# 1  pi=13'b1100111110000;
#1 $display("%b", po);
# 1  pi=13'b1100111110001;
#1 $display("%b", po);
# 1  pi=13'b1100111110010;
#1 $display("%b", po);
# 1  pi=13'b1100111110011;
#1 $display("%b", po);
# 1  pi=13'b1100111110100;
#1 $display("%b", po);
# 1  pi=13'b1100111110101;
#1 $display("%b", po);
# 1  pi=13'b1100111110110;
#1 $display("%b", po);
# 1  pi=13'b1100111110111;
#1 $display("%b", po);
# 1  pi=13'b1100111111000;
#1 $display("%b", po);
# 1  pi=13'b1100111111001;
#1 $display("%b", po);
# 1  pi=13'b1100111111010;
#1 $display("%b", po);
# 1  pi=13'b1100111111011;
#1 $display("%b", po);
# 1  pi=13'b1100111111100;
#1 $display("%b", po);
# 1  pi=13'b1100111111101;
#1 $display("%b", po);
# 1  pi=13'b1100111111110;
#1 $display("%b", po);
# 1  pi=13'b1100111111111;
#1 $display("%b", po);
# 1  pi=13'b1101000000000;
#1 $display("%b", po);
# 1  pi=13'b1101000000001;
#1 $display("%b", po);
# 1  pi=13'b1101000000010;
#1 $display("%b", po);
# 1  pi=13'b1101000000011;
#1 $display("%b", po);
# 1  pi=13'b1101000000100;
#1 $display("%b", po);
# 1  pi=13'b1101000000101;
#1 $display("%b", po);
# 1  pi=13'b1101000000110;
#1 $display("%b", po);
# 1  pi=13'b1101000000111;
#1 $display("%b", po);
# 1  pi=13'b1101000001000;
#1 $display("%b", po);
# 1  pi=13'b1101000001001;
#1 $display("%b", po);
# 1  pi=13'b1101000001010;
#1 $display("%b", po);
# 1  pi=13'b1101000001011;
#1 $display("%b", po);
# 1  pi=13'b1101000001100;
#1 $display("%b", po);
# 1  pi=13'b1101000001101;
#1 $display("%b", po);
# 1  pi=13'b1101000001110;
#1 $display("%b", po);
# 1  pi=13'b1101000001111;
#1 $display("%b", po);
# 1  pi=13'b1101000010000;
#1 $display("%b", po);
# 1  pi=13'b1101000010001;
#1 $display("%b", po);
# 1  pi=13'b1101000010010;
#1 $display("%b", po);
# 1  pi=13'b1101000010011;
#1 $display("%b", po);
# 1  pi=13'b1101000010100;
#1 $display("%b", po);
# 1  pi=13'b1101000010101;
#1 $display("%b", po);
# 1  pi=13'b1101000010110;
#1 $display("%b", po);
# 1  pi=13'b1101000010111;
#1 $display("%b", po);
# 1  pi=13'b1101000011000;
#1 $display("%b", po);
# 1  pi=13'b1101000011001;
#1 $display("%b", po);
# 1  pi=13'b1101000011010;
#1 $display("%b", po);
# 1  pi=13'b1101000011011;
#1 $display("%b", po);
# 1  pi=13'b1101000011100;
#1 $display("%b", po);
# 1  pi=13'b1101000011101;
#1 $display("%b", po);
# 1  pi=13'b1101000011110;
#1 $display("%b", po);
# 1  pi=13'b1101000011111;
#1 $display("%b", po);
# 1  pi=13'b1101000100000;
#1 $display("%b", po);
# 1  pi=13'b1101000100001;
#1 $display("%b", po);
# 1  pi=13'b1101000100010;
#1 $display("%b", po);
# 1  pi=13'b1101000100011;
#1 $display("%b", po);
# 1  pi=13'b1101000100100;
#1 $display("%b", po);
# 1  pi=13'b1101000100101;
#1 $display("%b", po);
# 1  pi=13'b1101000100110;
#1 $display("%b", po);
# 1  pi=13'b1101000100111;
#1 $display("%b", po);
# 1  pi=13'b1101000101000;
#1 $display("%b", po);
# 1  pi=13'b1101000101001;
#1 $display("%b", po);
# 1  pi=13'b1101000101010;
#1 $display("%b", po);
# 1  pi=13'b1101000101011;
#1 $display("%b", po);
# 1  pi=13'b1101000101100;
#1 $display("%b", po);
# 1  pi=13'b1101000101101;
#1 $display("%b", po);
# 1  pi=13'b1101000101110;
#1 $display("%b", po);
# 1  pi=13'b1101000101111;
#1 $display("%b", po);
# 1  pi=13'b1101000110000;
#1 $display("%b", po);
# 1  pi=13'b1101000110001;
#1 $display("%b", po);
# 1  pi=13'b1101000110010;
#1 $display("%b", po);
# 1  pi=13'b1101000110011;
#1 $display("%b", po);
# 1  pi=13'b1101000110100;
#1 $display("%b", po);
# 1  pi=13'b1101000110101;
#1 $display("%b", po);
# 1  pi=13'b1101000110110;
#1 $display("%b", po);
# 1  pi=13'b1101000110111;
#1 $display("%b", po);
# 1  pi=13'b1101000111000;
#1 $display("%b", po);
# 1  pi=13'b1101000111001;
#1 $display("%b", po);
# 1  pi=13'b1101000111010;
#1 $display("%b", po);
# 1  pi=13'b1101000111011;
#1 $display("%b", po);
# 1  pi=13'b1101000111100;
#1 $display("%b", po);
# 1  pi=13'b1101000111101;
#1 $display("%b", po);
# 1  pi=13'b1101000111110;
#1 $display("%b", po);
# 1  pi=13'b1101000111111;
#1 $display("%b", po);
# 1  pi=13'b1101001000000;
#1 $display("%b", po);
# 1  pi=13'b1101001000001;
#1 $display("%b", po);
# 1  pi=13'b1101001000010;
#1 $display("%b", po);
# 1  pi=13'b1101001000011;
#1 $display("%b", po);
# 1  pi=13'b1101001000100;
#1 $display("%b", po);
# 1  pi=13'b1101001000101;
#1 $display("%b", po);
# 1  pi=13'b1101001000110;
#1 $display("%b", po);
# 1  pi=13'b1101001000111;
#1 $display("%b", po);
# 1  pi=13'b1101001001000;
#1 $display("%b", po);
# 1  pi=13'b1101001001001;
#1 $display("%b", po);
# 1  pi=13'b1101001001010;
#1 $display("%b", po);
# 1  pi=13'b1101001001011;
#1 $display("%b", po);
# 1  pi=13'b1101001001100;
#1 $display("%b", po);
# 1  pi=13'b1101001001101;
#1 $display("%b", po);
# 1  pi=13'b1101001001110;
#1 $display("%b", po);
# 1  pi=13'b1101001001111;
#1 $display("%b", po);
# 1  pi=13'b1101001010000;
#1 $display("%b", po);
# 1  pi=13'b1101001010001;
#1 $display("%b", po);
# 1  pi=13'b1101001010010;
#1 $display("%b", po);
# 1  pi=13'b1101001010011;
#1 $display("%b", po);
# 1  pi=13'b1101001010100;
#1 $display("%b", po);
# 1  pi=13'b1101001010101;
#1 $display("%b", po);
# 1  pi=13'b1101001010110;
#1 $display("%b", po);
# 1  pi=13'b1101001010111;
#1 $display("%b", po);
# 1  pi=13'b1101001011000;
#1 $display("%b", po);
# 1  pi=13'b1101001011001;
#1 $display("%b", po);
# 1  pi=13'b1101001011010;
#1 $display("%b", po);
# 1  pi=13'b1101001011011;
#1 $display("%b", po);
# 1  pi=13'b1101001011100;
#1 $display("%b", po);
# 1  pi=13'b1101001011101;
#1 $display("%b", po);
# 1  pi=13'b1101001011110;
#1 $display("%b", po);
# 1  pi=13'b1101001011111;
#1 $display("%b", po);
# 1  pi=13'b1101001100000;
#1 $display("%b", po);
# 1  pi=13'b1101001100001;
#1 $display("%b", po);
# 1  pi=13'b1101001100010;
#1 $display("%b", po);
# 1  pi=13'b1101001100011;
#1 $display("%b", po);
# 1  pi=13'b1101001100100;
#1 $display("%b", po);
# 1  pi=13'b1101001100101;
#1 $display("%b", po);
# 1  pi=13'b1101001100110;
#1 $display("%b", po);
# 1  pi=13'b1101001100111;
#1 $display("%b", po);
# 1  pi=13'b1101001101000;
#1 $display("%b", po);
# 1  pi=13'b1101001101001;
#1 $display("%b", po);
# 1  pi=13'b1101001101010;
#1 $display("%b", po);
# 1  pi=13'b1101001101011;
#1 $display("%b", po);
# 1  pi=13'b1101001101100;
#1 $display("%b", po);
# 1  pi=13'b1101001101101;
#1 $display("%b", po);
# 1  pi=13'b1101001101110;
#1 $display("%b", po);
# 1  pi=13'b1101001101111;
#1 $display("%b", po);
# 1  pi=13'b1101001110000;
#1 $display("%b", po);
# 1  pi=13'b1101001110001;
#1 $display("%b", po);
# 1  pi=13'b1101001110010;
#1 $display("%b", po);
# 1  pi=13'b1101001110011;
#1 $display("%b", po);
# 1  pi=13'b1101001110100;
#1 $display("%b", po);
# 1  pi=13'b1101001110101;
#1 $display("%b", po);
# 1  pi=13'b1101001110110;
#1 $display("%b", po);
# 1  pi=13'b1101001110111;
#1 $display("%b", po);
# 1  pi=13'b1101001111000;
#1 $display("%b", po);
# 1  pi=13'b1101001111001;
#1 $display("%b", po);
# 1  pi=13'b1101001111010;
#1 $display("%b", po);
# 1  pi=13'b1101001111011;
#1 $display("%b", po);
# 1  pi=13'b1101001111100;
#1 $display("%b", po);
# 1  pi=13'b1101001111101;
#1 $display("%b", po);
# 1  pi=13'b1101001111110;
#1 $display("%b", po);
# 1  pi=13'b1101001111111;
#1 $display("%b", po);
# 1  pi=13'b1101010000000;
#1 $display("%b", po);
# 1  pi=13'b1101010000001;
#1 $display("%b", po);
# 1  pi=13'b1101010000010;
#1 $display("%b", po);
# 1  pi=13'b1101010000011;
#1 $display("%b", po);
# 1  pi=13'b1101010000100;
#1 $display("%b", po);
# 1  pi=13'b1101010000101;
#1 $display("%b", po);
# 1  pi=13'b1101010000110;
#1 $display("%b", po);
# 1  pi=13'b1101010000111;
#1 $display("%b", po);
# 1  pi=13'b1101010001000;
#1 $display("%b", po);
# 1  pi=13'b1101010001001;
#1 $display("%b", po);
# 1  pi=13'b1101010001010;
#1 $display("%b", po);
# 1  pi=13'b1101010001011;
#1 $display("%b", po);
# 1  pi=13'b1101010001100;
#1 $display("%b", po);
# 1  pi=13'b1101010001101;
#1 $display("%b", po);
# 1  pi=13'b1101010001110;
#1 $display("%b", po);
# 1  pi=13'b1101010001111;
#1 $display("%b", po);
# 1  pi=13'b1101010010000;
#1 $display("%b", po);
# 1  pi=13'b1101010010001;
#1 $display("%b", po);
# 1  pi=13'b1101010010010;
#1 $display("%b", po);
# 1  pi=13'b1101010010011;
#1 $display("%b", po);
# 1  pi=13'b1101010010100;
#1 $display("%b", po);
# 1  pi=13'b1101010010101;
#1 $display("%b", po);
# 1  pi=13'b1101010010110;
#1 $display("%b", po);
# 1  pi=13'b1101010010111;
#1 $display("%b", po);
# 1  pi=13'b1101010011000;
#1 $display("%b", po);
# 1  pi=13'b1101010011001;
#1 $display("%b", po);
# 1  pi=13'b1101010011010;
#1 $display("%b", po);
# 1  pi=13'b1101010011011;
#1 $display("%b", po);
# 1  pi=13'b1101010011100;
#1 $display("%b", po);
# 1  pi=13'b1101010011101;
#1 $display("%b", po);
# 1  pi=13'b1101010011110;
#1 $display("%b", po);
# 1  pi=13'b1101010011111;
#1 $display("%b", po);
# 1  pi=13'b1101010100000;
#1 $display("%b", po);
# 1  pi=13'b1101010100001;
#1 $display("%b", po);
# 1  pi=13'b1101010100010;
#1 $display("%b", po);
# 1  pi=13'b1101010100011;
#1 $display("%b", po);
# 1  pi=13'b1101010100100;
#1 $display("%b", po);
# 1  pi=13'b1101010100101;
#1 $display("%b", po);
# 1  pi=13'b1101010100110;
#1 $display("%b", po);
# 1  pi=13'b1101010100111;
#1 $display("%b", po);
# 1  pi=13'b1101010101000;
#1 $display("%b", po);
# 1  pi=13'b1101010101001;
#1 $display("%b", po);
# 1  pi=13'b1101010101010;
#1 $display("%b", po);
# 1  pi=13'b1101010101011;
#1 $display("%b", po);
# 1  pi=13'b1101010101100;
#1 $display("%b", po);
# 1  pi=13'b1101010101101;
#1 $display("%b", po);
# 1  pi=13'b1101010101110;
#1 $display("%b", po);
# 1  pi=13'b1101010101111;
#1 $display("%b", po);
# 1  pi=13'b1101010110000;
#1 $display("%b", po);
# 1  pi=13'b1101010110001;
#1 $display("%b", po);
# 1  pi=13'b1101010110010;
#1 $display("%b", po);
# 1  pi=13'b1101010110011;
#1 $display("%b", po);
# 1  pi=13'b1101010110100;
#1 $display("%b", po);
# 1  pi=13'b1101010110101;
#1 $display("%b", po);
# 1  pi=13'b1101010110110;
#1 $display("%b", po);
# 1  pi=13'b1101010110111;
#1 $display("%b", po);
# 1  pi=13'b1101010111000;
#1 $display("%b", po);
# 1  pi=13'b1101010111001;
#1 $display("%b", po);
# 1  pi=13'b1101010111010;
#1 $display("%b", po);
# 1  pi=13'b1101010111011;
#1 $display("%b", po);
# 1  pi=13'b1101010111100;
#1 $display("%b", po);
# 1  pi=13'b1101010111101;
#1 $display("%b", po);
# 1  pi=13'b1101010111110;
#1 $display("%b", po);
# 1  pi=13'b1101010111111;
#1 $display("%b", po);
# 1  pi=13'b1101011000000;
#1 $display("%b", po);
# 1  pi=13'b1101011000001;
#1 $display("%b", po);
# 1  pi=13'b1101011000010;
#1 $display("%b", po);
# 1  pi=13'b1101011000011;
#1 $display("%b", po);
# 1  pi=13'b1101011000100;
#1 $display("%b", po);
# 1  pi=13'b1101011000101;
#1 $display("%b", po);
# 1  pi=13'b1101011000110;
#1 $display("%b", po);
# 1  pi=13'b1101011000111;
#1 $display("%b", po);
# 1  pi=13'b1101011001000;
#1 $display("%b", po);
# 1  pi=13'b1101011001001;
#1 $display("%b", po);
# 1  pi=13'b1101011001010;
#1 $display("%b", po);
# 1  pi=13'b1101011001011;
#1 $display("%b", po);
# 1  pi=13'b1101011001100;
#1 $display("%b", po);
# 1  pi=13'b1101011001101;
#1 $display("%b", po);
# 1  pi=13'b1101011001110;
#1 $display("%b", po);
# 1  pi=13'b1101011001111;
#1 $display("%b", po);
# 1  pi=13'b1101011010000;
#1 $display("%b", po);
# 1  pi=13'b1101011010001;
#1 $display("%b", po);
# 1  pi=13'b1101011010010;
#1 $display("%b", po);
# 1  pi=13'b1101011010011;
#1 $display("%b", po);
# 1  pi=13'b1101011010100;
#1 $display("%b", po);
# 1  pi=13'b1101011010101;
#1 $display("%b", po);
# 1  pi=13'b1101011010110;
#1 $display("%b", po);
# 1  pi=13'b1101011010111;
#1 $display("%b", po);
# 1  pi=13'b1101011011000;
#1 $display("%b", po);
# 1  pi=13'b1101011011001;
#1 $display("%b", po);
# 1  pi=13'b1101011011010;
#1 $display("%b", po);
# 1  pi=13'b1101011011011;
#1 $display("%b", po);
# 1  pi=13'b1101011011100;
#1 $display("%b", po);
# 1  pi=13'b1101011011101;
#1 $display("%b", po);
# 1  pi=13'b1101011011110;
#1 $display("%b", po);
# 1  pi=13'b1101011011111;
#1 $display("%b", po);
# 1  pi=13'b1101011100000;
#1 $display("%b", po);
# 1  pi=13'b1101011100001;
#1 $display("%b", po);
# 1  pi=13'b1101011100010;
#1 $display("%b", po);
# 1  pi=13'b1101011100011;
#1 $display("%b", po);
# 1  pi=13'b1101011100100;
#1 $display("%b", po);
# 1  pi=13'b1101011100101;
#1 $display("%b", po);
# 1  pi=13'b1101011100110;
#1 $display("%b", po);
# 1  pi=13'b1101011100111;
#1 $display("%b", po);
# 1  pi=13'b1101011101000;
#1 $display("%b", po);
# 1  pi=13'b1101011101001;
#1 $display("%b", po);
# 1  pi=13'b1101011101010;
#1 $display("%b", po);
# 1  pi=13'b1101011101011;
#1 $display("%b", po);
# 1  pi=13'b1101011101100;
#1 $display("%b", po);
# 1  pi=13'b1101011101101;
#1 $display("%b", po);
# 1  pi=13'b1101011101110;
#1 $display("%b", po);
# 1  pi=13'b1101011101111;
#1 $display("%b", po);
# 1  pi=13'b1101011110000;
#1 $display("%b", po);
# 1  pi=13'b1101011110001;
#1 $display("%b", po);
# 1  pi=13'b1101011110010;
#1 $display("%b", po);
# 1  pi=13'b1101011110011;
#1 $display("%b", po);
# 1  pi=13'b1101011110100;
#1 $display("%b", po);
# 1  pi=13'b1101011110101;
#1 $display("%b", po);
# 1  pi=13'b1101011110110;
#1 $display("%b", po);
# 1  pi=13'b1101011110111;
#1 $display("%b", po);
# 1  pi=13'b1101011111000;
#1 $display("%b", po);
# 1  pi=13'b1101011111001;
#1 $display("%b", po);
# 1  pi=13'b1101011111010;
#1 $display("%b", po);
# 1  pi=13'b1101011111011;
#1 $display("%b", po);
# 1  pi=13'b1101011111100;
#1 $display("%b", po);
# 1  pi=13'b1101011111101;
#1 $display("%b", po);
# 1  pi=13'b1101011111110;
#1 $display("%b", po);
# 1  pi=13'b1101011111111;
#1 $display("%b", po);
# 1  pi=13'b1101100000000;
#1 $display("%b", po);
# 1  pi=13'b1101100000001;
#1 $display("%b", po);
# 1  pi=13'b1101100000010;
#1 $display("%b", po);
# 1  pi=13'b1101100000011;
#1 $display("%b", po);
# 1  pi=13'b1101100000100;
#1 $display("%b", po);
# 1  pi=13'b1101100000101;
#1 $display("%b", po);
# 1  pi=13'b1101100000110;
#1 $display("%b", po);
# 1  pi=13'b1101100000111;
#1 $display("%b", po);
# 1  pi=13'b1101100001000;
#1 $display("%b", po);
# 1  pi=13'b1101100001001;
#1 $display("%b", po);
# 1  pi=13'b1101100001010;
#1 $display("%b", po);
# 1  pi=13'b1101100001011;
#1 $display("%b", po);
# 1  pi=13'b1101100001100;
#1 $display("%b", po);
# 1  pi=13'b1101100001101;
#1 $display("%b", po);
# 1  pi=13'b1101100001110;
#1 $display("%b", po);
# 1  pi=13'b1101100001111;
#1 $display("%b", po);
# 1  pi=13'b1101100010000;
#1 $display("%b", po);
# 1  pi=13'b1101100010001;
#1 $display("%b", po);
# 1  pi=13'b1101100010010;
#1 $display("%b", po);
# 1  pi=13'b1101100010011;
#1 $display("%b", po);
# 1  pi=13'b1101100010100;
#1 $display("%b", po);
# 1  pi=13'b1101100010101;
#1 $display("%b", po);
# 1  pi=13'b1101100010110;
#1 $display("%b", po);
# 1  pi=13'b1101100010111;
#1 $display("%b", po);
# 1  pi=13'b1101100011000;
#1 $display("%b", po);
# 1  pi=13'b1101100011001;
#1 $display("%b", po);
# 1  pi=13'b1101100011010;
#1 $display("%b", po);
# 1  pi=13'b1101100011011;
#1 $display("%b", po);
# 1  pi=13'b1101100011100;
#1 $display("%b", po);
# 1  pi=13'b1101100011101;
#1 $display("%b", po);
# 1  pi=13'b1101100011110;
#1 $display("%b", po);
# 1  pi=13'b1101100011111;
#1 $display("%b", po);
# 1  pi=13'b1101100100000;
#1 $display("%b", po);
# 1  pi=13'b1101100100001;
#1 $display("%b", po);
# 1  pi=13'b1101100100010;
#1 $display("%b", po);
# 1  pi=13'b1101100100011;
#1 $display("%b", po);
# 1  pi=13'b1101100100100;
#1 $display("%b", po);
# 1  pi=13'b1101100100101;
#1 $display("%b", po);
# 1  pi=13'b1101100100110;
#1 $display("%b", po);
# 1  pi=13'b1101100100111;
#1 $display("%b", po);
# 1  pi=13'b1101100101000;
#1 $display("%b", po);
# 1  pi=13'b1101100101001;
#1 $display("%b", po);
# 1  pi=13'b1101100101010;
#1 $display("%b", po);
# 1  pi=13'b1101100101011;
#1 $display("%b", po);
# 1  pi=13'b1101100101100;
#1 $display("%b", po);
# 1  pi=13'b1101100101101;
#1 $display("%b", po);
# 1  pi=13'b1101100101110;
#1 $display("%b", po);
# 1  pi=13'b1101100101111;
#1 $display("%b", po);
# 1  pi=13'b1101100110000;
#1 $display("%b", po);
# 1  pi=13'b1101100110001;
#1 $display("%b", po);
# 1  pi=13'b1101100110010;
#1 $display("%b", po);
# 1  pi=13'b1101100110011;
#1 $display("%b", po);
# 1  pi=13'b1101100110100;
#1 $display("%b", po);
# 1  pi=13'b1101100110101;
#1 $display("%b", po);
# 1  pi=13'b1101100110110;
#1 $display("%b", po);
# 1  pi=13'b1101100110111;
#1 $display("%b", po);
# 1  pi=13'b1101100111000;
#1 $display("%b", po);
# 1  pi=13'b1101100111001;
#1 $display("%b", po);
# 1  pi=13'b1101100111010;
#1 $display("%b", po);
# 1  pi=13'b1101100111011;
#1 $display("%b", po);
# 1  pi=13'b1101100111100;
#1 $display("%b", po);
# 1  pi=13'b1101100111101;
#1 $display("%b", po);
# 1  pi=13'b1101100111110;
#1 $display("%b", po);
# 1  pi=13'b1101100111111;
#1 $display("%b", po);
# 1  pi=13'b1101101000000;
#1 $display("%b", po);
# 1  pi=13'b1101101000001;
#1 $display("%b", po);
# 1  pi=13'b1101101000010;
#1 $display("%b", po);
# 1  pi=13'b1101101000011;
#1 $display("%b", po);
# 1  pi=13'b1101101000100;
#1 $display("%b", po);
# 1  pi=13'b1101101000101;
#1 $display("%b", po);
# 1  pi=13'b1101101000110;
#1 $display("%b", po);
# 1  pi=13'b1101101000111;
#1 $display("%b", po);
# 1  pi=13'b1101101001000;
#1 $display("%b", po);
# 1  pi=13'b1101101001001;
#1 $display("%b", po);
# 1  pi=13'b1101101001010;
#1 $display("%b", po);
# 1  pi=13'b1101101001011;
#1 $display("%b", po);
# 1  pi=13'b1101101001100;
#1 $display("%b", po);
# 1  pi=13'b1101101001101;
#1 $display("%b", po);
# 1  pi=13'b1101101001110;
#1 $display("%b", po);
# 1  pi=13'b1101101001111;
#1 $display("%b", po);
# 1  pi=13'b1101101010000;
#1 $display("%b", po);
# 1  pi=13'b1101101010001;
#1 $display("%b", po);
# 1  pi=13'b1101101010010;
#1 $display("%b", po);
# 1  pi=13'b1101101010011;
#1 $display("%b", po);
# 1  pi=13'b1101101010100;
#1 $display("%b", po);
# 1  pi=13'b1101101010101;
#1 $display("%b", po);
# 1  pi=13'b1101101010110;
#1 $display("%b", po);
# 1  pi=13'b1101101010111;
#1 $display("%b", po);
# 1  pi=13'b1101101011000;
#1 $display("%b", po);
# 1  pi=13'b1101101011001;
#1 $display("%b", po);
# 1  pi=13'b1101101011010;
#1 $display("%b", po);
# 1  pi=13'b1101101011011;
#1 $display("%b", po);
# 1  pi=13'b1101101011100;
#1 $display("%b", po);
# 1  pi=13'b1101101011101;
#1 $display("%b", po);
# 1  pi=13'b1101101011110;
#1 $display("%b", po);
# 1  pi=13'b1101101011111;
#1 $display("%b", po);
# 1  pi=13'b1101101100000;
#1 $display("%b", po);
# 1  pi=13'b1101101100001;
#1 $display("%b", po);
# 1  pi=13'b1101101100010;
#1 $display("%b", po);
# 1  pi=13'b1101101100011;
#1 $display("%b", po);
# 1  pi=13'b1101101100100;
#1 $display("%b", po);
# 1  pi=13'b1101101100101;
#1 $display("%b", po);
# 1  pi=13'b1101101100110;
#1 $display("%b", po);
# 1  pi=13'b1101101100111;
#1 $display("%b", po);
# 1  pi=13'b1101101101000;
#1 $display("%b", po);
# 1  pi=13'b1101101101001;
#1 $display("%b", po);
# 1  pi=13'b1101101101010;
#1 $display("%b", po);
# 1  pi=13'b1101101101011;
#1 $display("%b", po);
# 1  pi=13'b1101101101100;
#1 $display("%b", po);
# 1  pi=13'b1101101101101;
#1 $display("%b", po);
# 1  pi=13'b1101101101110;
#1 $display("%b", po);
# 1  pi=13'b1101101101111;
#1 $display("%b", po);
# 1  pi=13'b1101101110000;
#1 $display("%b", po);
# 1  pi=13'b1101101110001;
#1 $display("%b", po);
# 1  pi=13'b1101101110010;
#1 $display("%b", po);
# 1  pi=13'b1101101110011;
#1 $display("%b", po);
# 1  pi=13'b1101101110100;
#1 $display("%b", po);
# 1  pi=13'b1101101110101;
#1 $display("%b", po);
# 1  pi=13'b1101101110110;
#1 $display("%b", po);
# 1  pi=13'b1101101110111;
#1 $display("%b", po);
# 1  pi=13'b1101101111000;
#1 $display("%b", po);
# 1  pi=13'b1101101111001;
#1 $display("%b", po);
# 1  pi=13'b1101101111010;
#1 $display("%b", po);
# 1  pi=13'b1101101111011;
#1 $display("%b", po);
# 1  pi=13'b1101101111100;
#1 $display("%b", po);
# 1  pi=13'b1101101111101;
#1 $display("%b", po);
# 1  pi=13'b1101101111110;
#1 $display("%b", po);
# 1  pi=13'b1101101111111;
#1 $display("%b", po);
# 1  pi=13'b1101110000000;
#1 $display("%b", po);
# 1  pi=13'b1101110000001;
#1 $display("%b", po);
# 1  pi=13'b1101110000010;
#1 $display("%b", po);
# 1  pi=13'b1101110000011;
#1 $display("%b", po);
# 1  pi=13'b1101110000100;
#1 $display("%b", po);
# 1  pi=13'b1101110000101;
#1 $display("%b", po);
# 1  pi=13'b1101110000110;
#1 $display("%b", po);
# 1  pi=13'b1101110000111;
#1 $display("%b", po);
# 1  pi=13'b1101110001000;
#1 $display("%b", po);
# 1  pi=13'b1101110001001;
#1 $display("%b", po);
# 1  pi=13'b1101110001010;
#1 $display("%b", po);
# 1  pi=13'b1101110001011;
#1 $display("%b", po);
# 1  pi=13'b1101110001100;
#1 $display("%b", po);
# 1  pi=13'b1101110001101;
#1 $display("%b", po);
# 1  pi=13'b1101110001110;
#1 $display("%b", po);
# 1  pi=13'b1101110001111;
#1 $display("%b", po);
# 1  pi=13'b1101110010000;
#1 $display("%b", po);
# 1  pi=13'b1101110010001;
#1 $display("%b", po);
# 1  pi=13'b1101110010010;
#1 $display("%b", po);
# 1  pi=13'b1101110010011;
#1 $display("%b", po);
# 1  pi=13'b1101110010100;
#1 $display("%b", po);
# 1  pi=13'b1101110010101;
#1 $display("%b", po);
# 1  pi=13'b1101110010110;
#1 $display("%b", po);
# 1  pi=13'b1101110010111;
#1 $display("%b", po);
# 1  pi=13'b1101110011000;
#1 $display("%b", po);
# 1  pi=13'b1101110011001;
#1 $display("%b", po);
# 1  pi=13'b1101110011010;
#1 $display("%b", po);
# 1  pi=13'b1101110011011;
#1 $display("%b", po);
# 1  pi=13'b1101110011100;
#1 $display("%b", po);
# 1  pi=13'b1101110011101;
#1 $display("%b", po);
# 1  pi=13'b1101110011110;
#1 $display("%b", po);
# 1  pi=13'b1101110011111;
#1 $display("%b", po);
# 1  pi=13'b1101110100000;
#1 $display("%b", po);
# 1  pi=13'b1101110100001;
#1 $display("%b", po);
# 1  pi=13'b1101110100010;
#1 $display("%b", po);
# 1  pi=13'b1101110100011;
#1 $display("%b", po);
# 1  pi=13'b1101110100100;
#1 $display("%b", po);
# 1  pi=13'b1101110100101;
#1 $display("%b", po);
# 1  pi=13'b1101110100110;
#1 $display("%b", po);
# 1  pi=13'b1101110100111;
#1 $display("%b", po);
# 1  pi=13'b1101110101000;
#1 $display("%b", po);
# 1  pi=13'b1101110101001;
#1 $display("%b", po);
# 1  pi=13'b1101110101010;
#1 $display("%b", po);
# 1  pi=13'b1101110101011;
#1 $display("%b", po);
# 1  pi=13'b1101110101100;
#1 $display("%b", po);
# 1  pi=13'b1101110101101;
#1 $display("%b", po);
# 1  pi=13'b1101110101110;
#1 $display("%b", po);
# 1  pi=13'b1101110101111;
#1 $display("%b", po);
# 1  pi=13'b1101110110000;
#1 $display("%b", po);
# 1  pi=13'b1101110110001;
#1 $display("%b", po);
# 1  pi=13'b1101110110010;
#1 $display("%b", po);
# 1  pi=13'b1101110110011;
#1 $display("%b", po);
# 1  pi=13'b1101110110100;
#1 $display("%b", po);
# 1  pi=13'b1101110110101;
#1 $display("%b", po);
# 1  pi=13'b1101110110110;
#1 $display("%b", po);
# 1  pi=13'b1101110110111;
#1 $display("%b", po);
# 1  pi=13'b1101110111000;
#1 $display("%b", po);
# 1  pi=13'b1101110111001;
#1 $display("%b", po);
# 1  pi=13'b1101110111010;
#1 $display("%b", po);
# 1  pi=13'b1101110111011;
#1 $display("%b", po);
# 1  pi=13'b1101110111100;
#1 $display("%b", po);
# 1  pi=13'b1101110111101;
#1 $display("%b", po);
# 1  pi=13'b1101110111110;
#1 $display("%b", po);
# 1  pi=13'b1101110111111;
#1 $display("%b", po);
# 1  pi=13'b1101111000000;
#1 $display("%b", po);
# 1  pi=13'b1101111000001;
#1 $display("%b", po);
# 1  pi=13'b1101111000010;
#1 $display("%b", po);
# 1  pi=13'b1101111000011;
#1 $display("%b", po);
# 1  pi=13'b1101111000100;
#1 $display("%b", po);
# 1  pi=13'b1101111000101;
#1 $display("%b", po);
# 1  pi=13'b1101111000110;
#1 $display("%b", po);
# 1  pi=13'b1101111000111;
#1 $display("%b", po);
# 1  pi=13'b1101111001000;
#1 $display("%b", po);
# 1  pi=13'b1101111001001;
#1 $display("%b", po);
# 1  pi=13'b1101111001010;
#1 $display("%b", po);
# 1  pi=13'b1101111001011;
#1 $display("%b", po);
# 1  pi=13'b1101111001100;
#1 $display("%b", po);
# 1  pi=13'b1101111001101;
#1 $display("%b", po);
# 1  pi=13'b1101111001110;
#1 $display("%b", po);
# 1  pi=13'b1101111001111;
#1 $display("%b", po);
# 1  pi=13'b1101111010000;
#1 $display("%b", po);
# 1  pi=13'b1101111010001;
#1 $display("%b", po);
# 1  pi=13'b1101111010010;
#1 $display("%b", po);
# 1  pi=13'b1101111010011;
#1 $display("%b", po);
# 1  pi=13'b1101111010100;
#1 $display("%b", po);
# 1  pi=13'b1101111010101;
#1 $display("%b", po);
# 1  pi=13'b1101111010110;
#1 $display("%b", po);
# 1  pi=13'b1101111010111;
#1 $display("%b", po);
# 1  pi=13'b1101111011000;
#1 $display("%b", po);
# 1  pi=13'b1101111011001;
#1 $display("%b", po);
# 1  pi=13'b1101111011010;
#1 $display("%b", po);
# 1  pi=13'b1101111011011;
#1 $display("%b", po);
# 1  pi=13'b1101111011100;
#1 $display("%b", po);
# 1  pi=13'b1101111011101;
#1 $display("%b", po);
# 1  pi=13'b1101111011110;
#1 $display("%b", po);
# 1  pi=13'b1101111011111;
#1 $display("%b", po);
# 1  pi=13'b1101111100000;
#1 $display("%b", po);
# 1  pi=13'b1101111100001;
#1 $display("%b", po);
# 1  pi=13'b1101111100010;
#1 $display("%b", po);
# 1  pi=13'b1101111100011;
#1 $display("%b", po);
# 1  pi=13'b1101111100100;
#1 $display("%b", po);
# 1  pi=13'b1101111100101;
#1 $display("%b", po);
# 1  pi=13'b1101111100110;
#1 $display("%b", po);
# 1  pi=13'b1101111100111;
#1 $display("%b", po);
# 1  pi=13'b1101111101000;
#1 $display("%b", po);
# 1  pi=13'b1101111101001;
#1 $display("%b", po);
# 1  pi=13'b1101111101010;
#1 $display("%b", po);
# 1  pi=13'b1101111101011;
#1 $display("%b", po);
# 1  pi=13'b1101111101100;
#1 $display("%b", po);
# 1  pi=13'b1101111101101;
#1 $display("%b", po);
# 1  pi=13'b1101111101110;
#1 $display("%b", po);
# 1  pi=13'b1101111101111;
#1 $display("%b", po);
# 1  pi=13'b1101111110000;
#1 $display("%b", po);
# 1  pi=13'b1101111110001;
#1 $display("%b", po);
# 1  pi=13'b1101111110010;
#1 $display("%b", po);
# 1  pi=13'b1101111110011;
#1 $display("%b", po);
# 1  pi=13'b1101111110100;
#1 $display("%b", po);
# 1  pi=13'b1101111110101;
#1 $display("%b", po);
# 1  pi=13'b1101111110110;
#1 $display("%b", po);
# 1  pi=13'b1101111110111;
#1 $display("%b", po);
# 1  pi=13'b1101111111000;
#1 $display("%b", po);
# 1  pi=13'b1101111111001;
#1 $display("%b", po);
# 1  pi=13'b1101111111010;
#1 $display("%b", po);
# 1  pi=13'b1101111111011;
#1 $display("%b", po);
# 1  pi=13'b1101111111100;
#1 $display("%b", po);
# 1  pi=13'b1101111111101;
#1 $display("%b", po);
# 1  pi=13'b1101111111110;
#1 $display("%b", po);
# 1  pi=13'b1101111111111;
#1 $display("%b", po);
# 1  pi=13'b1110000000000;
#1 $display("%b", po);
# 1  pi=13'b1110000000001;
#1 $display("%b", po);
# 1  pi=13'b1110000000010;
#1 $display("%b", po);
# 1  pi=13'b1110000000011;
#1 $display("%b", po);
# 1  pi=13'b1110000000100;
#1 $display("%b", po);
# 1  pi=13'b1110000000101;
#1 $display("%b", po);
# 1  pi=13'b1110000000110;
#1 $display("%b", po);
# 1  pi=13'b1110000000111;
#1 $display("%b", po);
# 1  pi=13'b1110000001000;
#1 $display("%b", po);
# 1  pi=13'b1110000001001;
#1 $display("%b", po);
# 1  pi=13'b1110000001010;
#1 $display("%b", po);
# 1  pi=13'b1110000001011;
#1 $display("%b", po);
# 1  pi=13'b1110000001100;
#1 $display("%b", po);
# 1  pi=13'b1110000001101;
#1 $display("%b", po);
# 1  pi=13'b1110000001110;
#1 $display("%b", po);
# 1  pi=13'b1110000001111;
#1 $display("%b", po);
# 1  pi=13'b1110000010000;
#1 $display("%b", po);
# 1  pi=13'b1110000010001;
#1 $display("%b", po);
# 1  pi=13'b1110000010010;
#1 $display("%b", po);
# 1  pi=13'b1110000010011;
#1 $display("%b", po);
# 1  pi=13'b1110000010100;
#1 $display("%b", po);
# 1  pi=13'b1110000010101;
#1 $display("%b", po);
# 1  pi=13'b1110000010110;
#1 $display("%b", po);
# 1  pi=13'b1110000010111;
#1 $display("%b", po);
# 1  pi=13'b1110000011000;
#1 $display("%b", po);
# 1  pi=13'b1110000011001;
#1 $display("%b", po);
# 1  pi=13'b1110000011010;
#1 $display("%b", po);
# 1  pi=13'b1110000011011;
#1 $display("%b", po);
# 1  pi=13'b1110000011100;
#1 $display("%b", po);
# 1  pi=13'b1110000011101;
#1 $display("%b", po);
# 1  pi=13'b1110000011110;
#1 $display("%b", po);
# 1  pi=13'b1110000011111;
#1 $display("%b", po);
# 1  pi=13'b1110000100000;
#1 $display("%b", po);
# 1  pi=13'b1110000100001;
#1 $display("%b", po);
# 1  pi=13'b1110000100010;
#1 $display("%b", po);
# 1  pi=13'b1110000100011;
#1 $display("%b", po);
# 1  pi=13'b1110000100100;
#1 $display("%b", po);
# 1  pi=13'b1110000100101;
#1 $display("%b", po);
# 1  pi=13'b1110000100110;
#1 $display("%b", po);
# 1  pi=13'b1110000100111;
#1 $display("%b", po);
# 1  pi=13'b1110000101000;
#1 $display("%b", po);
# 1  pi=13'b1110000101001;
#1 $display("%b", po);
# 1  pi=13'b1110000101010;
#1 $display("%b", po);
# 1  pi=13'b1110000101011;
#1 $display("%b", po);
# 1  pi=13'b1110000101100;
#1 $display("%b", po);
# 1  pi=13'b1110000101101;
#1 $display("%b", po);
# 1  pi=13'b1110000101110;
#1 $display("%b", po);
# 1  pi=13'b1110000101111;
#1 $display("%b", po);
# 1  pi=13'b1110000110000;
#1 $display("%b", po);
# 1  pi=13'b1110000110001;
#1 $display("%b", po);
# 1  pi=13'b1110000110010;
#1 $display("%b", po);
# 1  pi=13'b1110000110011;
#1 $display("%b", po);
# 1  pi=13'b1110000110100;
#1 $display("%b", po);
# 1  pi=13'b1110000110101;
#1 $display("%b", po);
# 1  pi=13'b1110000110110;
#1 $display("%b", po);
# 1  pi=13'b1110000110111;
#1 $display("%b", po);
# 1  pi=13'b1110000111000;
#1 $display("%b", po);
# 1  pi=13'b1110000111001;
#1 $display("%b", po);
# 1  pi=13'b1110000111010;
#1 $display("%b", po);
# 1  pi=13'b1110000111011;
#1 $display("%b", po);
# 1  pi=13'b1110000111100;
#1 $display("%b", po);
# 1  pi=13'b1110000111101;
#1 $display("%b", po);
# 1  pi=13'b1110000111110;
#1 $display("%b", po);
# 1  pi=13'b1110000111111;
#1 $display("%b", po);
# 1  pi=13'b1110001000000;
#1 $display("%b", po);
# 1  pi=13'b1110001000001;
#1 $display("%b", po);
# 1  pi=13'b1110001000010;
#1 $display("%b", po);
# 1  pi=13'b1110001000011;
#1 $display("%b", po);
# 1  pi=13'b1110001000100;
#1 $display("%b", po);
# 1  pi=13'b1110001000101;
#1 $display("%b", po);
# 1  pi=13'b1110001000110;
#1 $display("%b", po);
# 1  pi=13'b1110001000111;
#1 $display("%b", po);
# 1  pi=13'b1110001001000;
#1 $display("%b", po);
# 1  pi=13'b1110001001001;
#1 $display("%b", po);
# 1  pi=13'b1110001001010;
#1 $display("%b", po);
# 1  pi=13'b1110001001011;
#1 $display("%b", po);
# 1  pi=13'b1110001001100;
#1 $display("%b", po);
# 1  pi=13'b1110001001101;
#1 $display("%b", po);
# 1  pi=13'b1110001001110;
#1 $display("%b", po);
# 1  pi=13'b1110001001111;
#1 $display("%b", po);
# 1  pi=13'b1110001010000;
#1 $display("%b", po);
# 1  pi=13'b1110001010001;
#1 $display("%b", po);
# 1  pi=13'b1110001010010;
#1 $display("%b", po);
# 1  pi=13'b1110001010011;
#1 $display("%b", po);
# 1  pi=13'b1110001010100;
#1 $display("%b", po);
# 1  pi=13'b1110001010101;
#1 $display("%b", po);
# 1  pi=13'b1110001010110;
#1 $display("%b", po);
# 1  pi=13'b1110001010111;
#1 $display("%b", po);
# 1  pi=13'b1110001011000;
#1 $display("%b", po);
# 1  pi=13'b1110001011001;
#1 $display("%b", po);
# 1  pi=13'b1110001011010;
#1 $display("%b", po);
# 1  pi=13'b1110001011011;
#1 $display("%b", po);
# 1  pi=13'b1110001011100;
#1 $display("%b", po);
# 1  pi=13'b1110001011101;
#1 $display("%b", po);
# 1  pi=13'b1110001011110;
#1 $display("%b", po);
# 1  pi=13'b1110001011111;
#1 $display("%b", po);
# 1  pi=13'b1110001100000;
#1 $display("%b", po);
# 1  pi=13'b1110001100001;
#1 $display("%b", po);
# 1  pi=13'b1110001100010;
#1 $display("%b", po);
# 1  pi=13'b1110001100011;
#1 $display("%b", po);
# 1  pi=13'b1110001100100;
#1 $display("%b", po);
# 1  pi=13'b1110001100101;
#1 $display("%b", po);
# 1  pi=13'b1110001100110;
#1 $display("%b", po);
# 1  pi=13'b1110001100111;
#1 $display("%b", po);
# 1  pi=13'b1110001101000;
#1 $display("%b", po);
# 1  pi=13'b1110001101001;
#1 $display("%b", po);
# 1  pi=13'b1110001101010;
#1 $display("%b", po);
# 1  pi=13'b1110001101011;
#1 $display("%b", po);
# 1  pi=13'b1110001101100;
#1 $display("%b", po);
# 1  pi=13'b1110001101101;
#1 $display("%b", po);
# 1  pi=13'b1110001101110;
#1 $display("%b", po);
# 1  pi=13'b1110001101111;
#1 $display("%b", po);
# 1  pi=13'b1110001110000;
#1 $display("%b", po);
# 1  pi=13'b1110001110001;
#1 $display("%b", po);
# 1  pi=13'b1110001110010;
#1 $display("%b", po);
# 1  pi=13'b1110001110011;
#1 $display("%b", po);
# 1  pi=13'b1110001110100;
#1 $display("%b", po);
# 1  pi=13'b1110001110101;
#1 $display("%b", po);
# 1  pi=13'b1110001110110;
#1 $display("%b", po);
# 1  pi=13'b1110001110111;
#1 $display("%b", po);
# 1  pi=13'b1110001111000;
#1 $display("%b", po);
# 1  pi=13'b1110001111001;
#1 $display("%b", po);
# 1  pi=13'b1110001111010;
#1 $display("%b", po);
# 1  pi=13'b1110001111011;
#1 $display("%b", po);
# 1  pi=13'b1110001111100;
#1 $display("%b", po);
# 1  pi=13'b1110001111101;
#1 $display("%b", po);
# 1  pi=13'b1110001111110;
#1 $display("%b", po);
# 1  pi=13'b1110001111111;
#1 $display("%b", po);
# 1  pi=13'b1110010000000;
#1 $display("%b", po);
# 1  pi=13'b1110010000001;
#1 $display("%b", po);
# 1  pi=13'b1110010000010;
#1 $display("%b", po);
# 1  pi=13'b1110010000011;
#1 $display("%b", po);
# 1  pi=13'b1110010000100;
#1 $display("%b", po);
# 1  pi=13'b1110010000101;
#1 $display("%b", po);
# 1  pi=13'b1110010000110;
#1 $display("%b", po);
# 1  pi=13'b1110010000111;
#1 $display("%b", po);
# 1  pi=13'b1110010001000;
#1 $display("%b", po);
# 1  pi=13'b1110010001001;
#1 $display("%b", po);
# 1  pi=13'b1110010001010;
#1 $display("%b", po);
# 1  pi=13'b1110010001011;
#1 $display("%b", po);
# 1  pi=13'b1110010001100;
#1 $display("%b", po);
# 1  pi=13'b1110010001101;
#1 $display("%b", po);
# 1  pi=13'b1110010001110;
#1 $display("%b", po);
# 1  pi=13'b1110010001111;
#1 $display("%b", po);
# 1  pi=13'b1110010010000;
#1 $display("%b", po);
# 1  pi=13'b1110010010001;
#1 $display("%b", po);
# 1  pi=13'b1110010010010;
#1 $display("%b", po);
# 1  pi=13'b1110010010011;
#1 $display("%b", po);
# 1  pi=13'b1110010010100;
#1 $display("%b", po);
# 1  pi=13'b1110010010101;
#1 $display("%b", po);
# 1  pi=13'b1110010010110;
#1 $display("%b", po);
# 1  pi=13'b1110010010111;
#1 $display("%b", po);
# 1  pi=13'b1110010011000;
#1 $display("%b", po);
# 1  pi=13'b1110010011001;
#1 $display("%b", po);
# 1  pi=13'b1110010011010;
#1 $display("%b", po);
# 1  pi=13'b1110010011011;
#1 $display("%b", po);
# 1  pi=13'b1110010011100;
#1 $display("%b", po);
# 1  pi=13'b1110010011101;
#1 $display("%b", po);
# 1  pi=13'b1110010011110;
#1 $display("%b", po);
# 1  pi=13'b1110010011111;
#1 $display("%b", po);
# 1  pi=13'b1110010100000;
#1 $display("%b", po);
# 1  pi=13'b1110010100001;
#1 $display("%b", po);
# 1  pi=13'b1110010100010;
#1 $display("%b", po);
# 1  pi=13'b1110010100011;
#1 $display("%b", po);
# 1  pi=13'b1110010100100;
#1 $display("%b", po);
# 1  pi=13'b1110010100101;
#1 $display("%b", po);
# 1  pi=13'b1110010100110;
#1 $display("%b", po);
# 1  pi=13'b1110010100111;
#1 $display("%b", po);
# 1  pi=13'b1110010101000;
#1 $display("%b", po);
# 1  pi=13'b1110010101001;
#1 $display("%b", po);
# 1  pi=13'b1110010101010;
#1 $display("%b", po);
# 1  pi=13'b1110010101011;
#1 $display("%b", po);
# 1  pi=13'b1110010101100;
#1 $display("%b", po);
# 1  pi=13'b1110010101101;
#1 $display("%b", po);
# 1  pi=13'b1110010101110;
#1 $display("%b", po);
# 1  pi=13'b1110010101111;
#1 $display("%b", po);
# 1  pi=13'b1110010110000;
#1 $display("%b", po);
# 1  pi=13'b1110010110001;
#1 $display("%b", po);
# 1  pi=13'b1110010110010;
#1 $display("%b", po);
# 1  pi=13'b1110010110011;
#1 $display("%b", po);
# 1  pi=13'b1110010110100;
#1 $display("%b", po);
# 1  pi=13'b1110010110101;
#1 $display("%b", po);
# 1  pi=13'b1110010110110;
#1 $display("%b", po);
# 1  pi=13'b1110010110111;
#1 $display("%b", po);
# 1  pi=13'b1110010111000;
#1 $display("%b", po);
# 1  pi=13'b1110010111001;
#1 $display("%b", po);
# 1  pi=13'b1110010111010;
#1 $display("%b", po);
# 1  pi=13'b1110010111011;
#1 $display("%b", po);
# 1  pi=13'b1110010111100;
#1 $display("%b", po);
# 1  pi=13'b1110010111101;
#1 $display("%b", po);
# 1  pi=13'b1110010111110;
#1 $display("%b", po);
# 1  pi=13'b1110010111111;
#1 $display("%b", po);
# 1  pi=13'b1110011000000;
#1 $display("%b", po);
# 1  pi=13'b1110011000001;
#1 $display("%b", po);
# 1  pi=13'b1110011000010;
#1 $display("%b", po);
# 1  pi=13'b1110011000011;
#1 $display("%b", po);
# 1  pi=13'b1110011000100;
#1 $display("%b", po);
# 1  pi=13'b1110011000101;
#1 $display("%b", po);
# 1  pi=13'b1110011000110;
#1 $display("%b", po);
# 1  pi=13'b1110011000111;
#1 $display("%b", po);
# 1  pi=13'b1110011001000;
#1 $display("%b", po);
# 1  pi=13'b1110011001001;
#1 $display("%b", po);
# 1  pi=13'b1110011001010;
#1 $display("%b", po);
# 1  pi=13'b1110011001011;
#1 $display("%b", po);
# 1  pi=13'b1110011001100;
#1 $display("%b", po);
# 1  pi=13'b1110011001101;
#1 $display("%b", po);
# 1  pi=13'b1110011001110;
#1 $display("%b", po);
# 1  pi=13'b1110011001111;
#1 $display("%b", po);
# 1  pi=13'b1110011010000;
#1 $display("%b", po);
# 1  pi=13'b1110011010001;
#1 $display("%b", po);
# 1  pi=13'b1110011010010;
#1 $display("%b", po);
# 1  pi=13'b1110011010011;
#1 $display("%b", po);
# 1  pi=13'b1110011010100;
#1 $display("%b", po);
# 1  pi=13'b1110011010101;
#1 $display("%b", po);
# 1  pi=13'b1110011010110;
#1 $display("%b", po);
# 1  pi=13'b1110011010111;
#1 $display("%b", po);
# 1  pi=13'b1110011011000;
#1 $display("%b", po);
# 1  pi=13'b1110011011001;
#1 $display("%b", po);
# 1  pi=13'b1110011011010;
#1 $display("%b", po);
# 1  pi=13'b1110011011011;
#1 $display("%b", po);
# 1  pi=13'b1110011011100;
#1 $display("%b", po);
# 1  pi=13'b1110011011101;
#1 $display("%b", po);
# 1  pi=13'b1110011011110;
#1 $display("%b", po);
# 1  pi=13'b1110011011111;
#1 $display("%b", po);
# 1  pi=13'b1110011100000;
#1 $display("%b", po);
# 1  pi=13'b1110011100001;
#1 $display("%b", po);
# 1  pi=13'b1110011100010;
#1 $display("%b", po);
# 1  pi=13'b1110011100011;
#1 $display("%b", po);
# 1  pi=13'b1110011100100;
#1 $display("%b", po);
# 1  pi=13'b1110011100101;
#1 $display("%b", po);
# 1  pi=13'b1110011100110;
#1 $display("%b", po);
# 1  pi=13'b1110011100111;
#1 $display("%b", po);
# 1  pi=13'b1110011101000;
#1 $display("%b", po);
# 1  pi=13'b1110011101001;
#1 $display("%b", po);
# 1  pi=13'b1110011101010;
#1 $display("%b", po);
# 1  pi=13'b1110011101011;
#1 $display("%b", po);
# 1  pi=13'b1110011101100;
#1 $display("%b", po);
# 1  pi=13'b1110011101101;
#1 $display("%b", po);
# 1  pi=13'b1110011101110;
#1 $display("%b", po);
# 1  pi=13'b1110011101111;
#1 $display("%b", po);
# 1  pi=13'b1110011110000;
#1 $display("%b", po);
# 1  pi=13'b1110011110001;
#1 $display("%b", po);
# 1  pi=13'b1110011110010;
#1 $display("%b", po);
# 1  pi=13'b1110011110011;
#1 $display("%b", po);
# 1  pi=13'b1110011110100;
#1 $display("%b", po);
# 1  pi=13'b1110011110101;
#1 $display("%b", po);
# 1  pi=13'b1110011110110;
#1 $display("%b", po);
# 1  pi=13'b1110011110111;
#1 $display("%b", po);
# 1  pi=13'b1110011111000;
#1 $display("%b", po);
# 1  pi=13'b1110011111001;
#1 $display("%b", po);
# 1  pi=13'b1110011111010;
#1 $display("%b", po);
# 1  pi=13'b1110011111011;
#1 $display("%b", po);
# 1  pi=13'b1110011111100;
#1 $display("%b", po);
# 1  pi=13'b1110011111101;
#1 $display("%b", po);
# 1  pi=13'b1110011111110;
#1 $display("%b", po);
# 1  pi=13'b1110011111111;
#1 $display("%b", po);
# 1  pi=13'b1110100000000;
#1 $display("%b", po);
# 1  pi=13'b1110100000001;
#1 $display("%b", po);
# 1  pi=13'b1110100000010;
#1 $display("%b", po);
# 1  pi=13'b1110100000011;
#1 $display("%b", po);
# 1  pi=13'b1110100000100;
#1 $display("%b", po);
# 1  pi=13'b1110100000101;
#1 $display("%b", po);
# 1  pi=13'b1110100000110;
#1 $display("%b", po);
# 1  pi=13'b1110100000111;
#1 $display("%b", po);
# 1  pi=13'b1110100001000;
#1 $display("%b", po);
# 1  pi=13'b1110100001001;
#1 $display("%b", po);
# 1  pi=13'b1110100001010;
#1 $display("%b", po);
# 1  pi=13'b1110100001011;
#1 $display("%b", po);
# 1  pi=13'b1110100001100;
#1 $display("%b", po);
# 1  pi=13'b1110100001101;
#1 $display("%b", po);
# 1  pi=13'b1110100001110;
#1 $display("%b", po);
# 1  pi=13'b1110100001111;
#1 $display("%b", po);
# 1  pi=13'b1110100010000;
#1 $display("%b", po);
# 1  pi=13'b1110100010001;
#1 $display("%b", po);
# 1  pi=13'b1110100010010;
#1 $display("%b", po);
# 1  pi=13'b1110100010011;
#1 $display("%b", po);
# 1  pi=13'b1110100010100;
#1 $display("%b", po);
# 1  pi=13'b1110100010101;
#1 $display("%b", po);
# 1  pi=13'b1110100010110;
#1 $display("%b", po);
# 1  pi=13'b1110100010111;
#1 $display("%b", po);
# 1  pi=13'b1110100011000;
#1 $display("%b", po);
# 1  pi=13'b1110100011001;
#1 $display("%b", po);
# 1  pi=13'b1110100011010;
#1 $display("%b", po);
# 1  pi=13'b1110100011011;
#1 $display("%b", po);
# 1  pi=13'b1110100011100;
#1 $display("%b", po);
# 1  pi=13'b1110100011101;
#1 $display("%b", po);
# 1  pi=13'b1110100011110;
#1 $display("%b", po);
# 1  pi=13'b1110100011111;
#1 $display("%b", po);
# 1  pi=13'b1110100100000;
#1 $display("%b", po);
# 1  pi=13'b1110100100001;
#1 $display("%b", po);
# 1  pi=13'b1110100100010;
#1 $display("%b", po);
# 1  pi=13'b1110100100011;
#1 $display("%b", po);
# 1  pi=13'b1110100100100;
#1 $display("%b", po);
# 1  pi=13'b1110100100101;
#1 $display("%b", po);
# 1  pi=13'b1110100100110;
#1 $display("%b", po);
# 1  pi=13'b1110100100111;
#1 $display("%b", po);
# 1  pi=13'b1110100101000;
#1 $display("%b", po);
# 1  pi=13'b1110100101001;
#1 $display("%b", po);
# 1  pi=13'b1110100101010;
#1 $display("%b", po);
# 1  pi=13'b1110100101011;
#1 $display("%b", po);
# 1  pi=13'b1110100101100;
#1 $display("%b", po);
# 1  pi=13'b1110100101101;
#1 $display("%b", po);
# 1  pi=13'b1110100101110;
#1 $display("%b", po);
# 1  pi=13'b1110100101111;
#1 $display("%b", po);
# 1  pi=13'b1110100110000;
#1 $display("%b", po);
# 1  pi=13'b1110100110001;
#1 $display("%b", po);
# 1  pi=13'b1110100110010;
#1 $display("%b", po);
# 1  pi=13'b1110100110011;
#1 $display("%b", po);
# 1  pi=13'b1110100110100;
#1 $display("%b", po);
# 1  pi=13'b1110100110101;
#1 $display("%b", po);
# 1  pi=13'b1110100110110;
#1 $display("%b", po);
# 1  pi=13'b1110100110111;
#1 $display("%b", po);
# 1  pi=13'b1110100111000;
#1 $display("%b", po);
# 1  pi=13'b1110100111001;
#1 $display("%b", po);
# 1  pi=13'b1110100111010;
#1 $display("%b", po);
# 1  pi=13'b1110100111011;
#1 $display("%b", po);
# 1  pi=13'b1110100111100;
#1 $display("%b", po);
# 1  pi=13'b1110100111101;
#1 $display("%b", po);
# 1  pi=13'b1110100111110;
#1 $display("%b", po);
# 1  pi=13'b1110100111111;
#1 $display("%b", po);
# 1  pi=13'b1110101000000;
#1 $display("%b", po);
# 1  pi=13'b1110101000001;
#1 $display("%b", po);
# 1  pi=13'b1110101000010;
#1 $display("%b", po);
# 1  pi=13'b1110101000011;
#1 $display("%b", po);
# 1  pi=13'b1110101000100;
#1 $display("%b", po);
# 1  pi=13'b1110101000101;
#1 $display("%b", po);
# 1  pi=13'b1110101000110;
#1 $display("%b", po);
# 1  pi=13'b1110101000111;
#1 $display("%b", po);
# 1  pi=13'b1110101001000;
#1 $display("%b", po);
# 1  pi=13'b1110101001001;
#1 $display("%b", po);
# 1  pi=13'b1110101001010;
#1 $display("%b", po);
# 1  pi=13'b1110101001011;
#1 $display("%b", po);
# 1  pi=13'b1110101001100;
#1 $display("%b", po);
# 1  pi=13'b1110101001101;
#1 $display("%b", po);
# 1  pi=13'b1110101001110;
#1 $display("%b", po);
# 1  pi=13'b1110101001111;
#1 $display("%b", po);
# 1  pi=13'b1110101010000;
#1 $display("%b", po);
# 1  pi=13'b1110101010001;
#1 $display("%b", po);
# 1  pi=13'b1110101010010;
#1 $display("%b", po);
# 1  pi=13'b1110101010011;
#1 $display("%b", po);
# 1  pi=13'b1110101010100;
#1 $display("%b", po);
# 1  pi=13'b1110101010101;
#1 $display("%b", po);
# 1  pi=13'b1110101010110;
#1 $display("%b", po);
# 1  pi=13'b1110101010111;
#1 $display("%b", po);
# 1  pi=13'b1110101011000;
#1 $display("%b", po);
# 1  pi=13'b1110101011001;
#1 $display("%b", po);
# 1  pi=13'b1110101011010;
#1 $display("%b", po);
# 1  pi=13'b1110101011011;
#1 $display("%b", po);
# 1  pi=13'b1110101011100;
#1 $display("%b", po);
# 1  pi=13'b1110101011101;
#1 $display("%b", po);
# 1  pi=13'b1110101011110;
#1 $display("%b", po);
# 1  pi=13'b1110101011111;
#1 $display("%b", po);
# 1  pi=13'b1110101100000;
#1 $display("%b", po);
# 1  pi=13'b1110101100001;
#1 $display("%b", po);
# 1  pi=13'b1110101100010;
#1 $display("%b", po);
# 1  pi=13'b1110101100011;
#1 $display("%b", po);
# 1  pi=13'b1110101100100;
#1 $display("%b", po);
# 1  pi=13'b1110101100101;
#1 $display("%b", po);
# 1  pi=13'b1110101100110;
#1 $display("%b", po);
# 1  pi=13'b1110101100111;
#1 $display("%b", po);
# 1  pi=13'b1110101101000;
#1 $display("%b", po);
# 1  pi=13'b1110101101001;
#1 $display("%b", po);
# 1  pi=13'b1110101101010;
#1 $display("%b", po);
# 1  pi=13'b1110101101011;
#1 $display("%b", po);
# 1  pi=13'b1110101101100;
#1 $display("%b", po);
# 1  pi=13'b1110101101101;
#1 $display("%b", po);
# 1  pi=13'b1110101101110;
#1 $display("%b", po);
# 1  pi=13'b1110101101111;
#1 $display("%b", po);
# 1  pi=13'b1110101110000;
#1 $display("%b", po);
# 1  pi=13'b1110101110001;
#1 $display("%b", po);
# 1  pi=13'b1110101110010;
#1 $display("%b", po);
# 1  pi=13'b1110101110011;
#1 $display("%b", po);
# 1  pi=13'b1110101110100;
#1 $display("%b", po);
# 1  pi=13'b1110101110101;
#1 $display("%b", po);
# 1  pi=13'b1110101110110;
#1 $display("%b", po);
# 1  pi=13'b1110101110111;
#1 $display("%b", po);
# 1  pi=13'b1110101111000;
#1 $display("%b", po);
# 1  pi=13'b1110101111001;
#1 $display("%b", po);
# 1  pi=13'b1110101111010;
#1 $display("%b", po);
# 1  pi=13'b1110101111011;
#1 $display("%b", po);
# 1  pi=13'b1110101111100;
#1 $display("%b", po);
# 1  pi=13'b1110101111101;
#1 $display("%b", po);
# 1  pi=13'b1110101111110;
#1 $display("%b", po);
# 1  pi=13'b1110101111111;
#1 $display("%b", po);
# 1  pi=13'b1110110000000;
#1 $display("%b", po);
# 1  pi=13'b1110110000001;
#1 $display("%b", po);
# 1  pi=13'b1110110000010;
#1 $display("%b", po);
# 1  pi=13'b1110110000011;
#1 $display("%b", po);
# 1  pi=13'b1110110000100;
#1 $display("%b", po);
# 1  pi=13'b1110110000101;
#1 $display("%b", po);
# 1  pi=13'b1110110000110;
#1 $display("%b", po);
# 1  pi=13'b1110110000111;
#1 $display("%b", po);
# 1  pi=13'b1110110001000;
#1 $display("%b", po);
# 1  pi=13'b1110110001001;
#1 $display("%b", po);
# 1  pi=13'b1110110001010;
#1 $display("%b", po);
# 1  pi=13'b1110110001011;
#1 $display("%b", po);
# 1  pi=13'b1110110001100;
#1 $display("%b", po);
# 1  pi=13'b1110110001101;
#1 $display("%b", po);
# 1  pi=13'b1110110001110;
#1 $display("%b", po);
# 1  pi=13'b1110110001111;
#1 $display("%b", po);
# 1  pi=13'b1110110010000;
#1 $display("%b", po);
# 1  pi=13'b1110110010001;
#1 $display("%b", po);
# 1  pi=13'b1110110010010;
#1 $display("%b", po);
# 1  pi=13'b1110110010011;
#1 $display("%b", po);
# 1  pi=13'b1110110010100;
#1 $display("%b", po);
# 1  pi=13'b1110110010101;
#1 $display("%b", po);
# 1  pi=13'b1110110010110;
#1 $display("%b", po);
# 1  pi=13'b1110110010111;
#1 $display("%b", po);
# 1  pi=13'b1110110011000;
#1 $display("%b", po);
# 1  pi=13'b1110110011001;
#1 $display("%b", po);
# 1  pi=13'b1110110011010;
#1 $display("%b", po);
# 1  pi=13'b1110110011011;
#1 $display("%b", po);
# 1  pi=13'b1110110011100;
#1 $display("%b", po);
# 1  pi=13'b1110110011101;
#1 $display("%b", po);
# 1  pi=13'b1110110011110;
#1 $display("%b", po);
# 1  pi=13'b1110110011111;
#1 $display("%b", po);
# 1  pi=13'b1110110100000;
#1 $display("%b", po);
# 1  pi=13'b1110110100001;
#1 $display("%b", po);
# 1  pi=13'b1110110100010;
#1 $display("%b", po);
# 1  pi=13'b1110110100011;
#1 $display("%b", po);
# 1  pi=13'b1110110100100;
#1 $display("%b", po);
# 1  pi=13'b1110110100101;
#1 $display("%b", po);
# 1  pi=13'b1110110100110;
#1 $display("%b", po);
# 1  pi=13'b1110110100111;
#1 $display("%b", po);
# 1  pi=13'b1110110101000;
#1 $display("%b", po);
# 1  pi=13'b1110110101001;
#1 $display("%b", po);
# 1  pi=13'b1110110101010;
#1 $display("%b", po);
# 1  pi=13'b1110110101011;
#1 $display("%b", po);
# 1  pi=13'b1110110101100;
#1 $display("%b", po);
# 1  pi=13'b1110110101101;
#1 $display("%b", po);
# 1  pi=13'b1110110101110;
#1 $display("%b", po);
# 1  pi=13'b1110110101111;
#1 $display("%b", po);
# 1  pi=13'b1110110110000;
#1 $display("%b", po);
# 1  pi=13'b1110110110001;
#1 $display("%b", po);
# 1  pi=13'b1110110110010;
#1 $display("%b", po);
# 1  pi=13'b1110110110011;
#1 $display("%b", po);
# 1  pi=13'b1110110110100;
#1 $display("%b", po);
# 1  pi=13'b1110110110101;
#1 $display("%b", po);
# 1  pi=13'b1110110110110;
#1 $display("%b", po);
# 1  pi=13'b1110110110111;
#1 $display("%b", po);
# 1  pi=13'b1110110111000;
#1 $display("%b", po);
# 1  pi=13'b1110110111001;
#1 $display("%b", po);
# 1  pi=13'b1110110111010;
#1 $display("%b", po);
# 1  pi=13'b1110110111011;
#1 $display("%b", po);
# 1  pi=13'b1110110111100;
#1 $display("%b", po);
# 1  pi=13'b1110110111101;
#1 $display("%b", po);
# 1  pi=13'b1110110111110;
#1 $display("%b", po);
# 1  pi=13'b1110110111111;
#1 $display("%b", po);
# 1  pi=13'b1110111000000;
#1 $display("%b", po);
# 1  pi=13'b1110111000001;
#1 $display("%b", po);
# 1  pi=13'b1110111000010;
#1 $display("%b", po);
# 1  pi=13'b1110111000011;
#1 $display("%b", po);
# 1  pi=13'b1110111000100;
#1 $display("%b", po);
# 1  pi=13'b1110111000101;
#1 $display("%b", po);
# 1  pi=13'b1110111000110;
#1 $display("%b", po);
# 1  pi=13'b1110111000111;
#1 $display("%b", po);
# 1  pi=13'b1110111001000;
#1 $display("%b", po);
# 1  pi=13'b1110111001001;
#1 $display("%b", po);
# 1  pi=13'b1110111001010;
#1 $display("%b", po);
# 1  pi=13'b1110111001011;
#1 $display("%b", po);
# 1  pi=13'b1110111001100;
#1 $display("%b", po);
# 1  pi=13'b1110111001101;
#1 $display("%b", po);
# 1  pi=13'b1110111001110;
#1 $display("%b", po);
# 1  pi=13'b1110111001111;
#1 $display("%b", po);
# 1  pi=13'b1110111010000;
#1 $display("%b", po);
# 1  pi=13'b1110111010001;
#1 $display("%b", po);
# 1  pi=13'b1110111010010;
#1 $display("%b", po);
# 1  pi=13'b1110111010011;
#1 $display("%b", po);
# 1  pi=13'b1110111010100;
#1 $display("%b", po);
# 1  pi=13'b1110111010101;
#1 $display("%b", po);
# 1  pi=13'b1110111010110;
#1 $display("%b", po);
# 1  pi=13'b1110111010111;
#1 $display("%b", po);
# 1  pi=13'b1110111011000;
#1 $display("%b", po);
# 1  pi=13'b1110111011001;
#1 $display("%b", po);
# 1  pi=13'b1110111011010;
#1 $display("%b", po);
# 1  pi=13'b1110111011011;
#1 $display("%b", po);
# 1  pi=13'b1110111011100;
#1 $display("%b", po);
# 1  pi=13'b1110111011101;
#1 $display("%b", po);
# 1  pi=13'b1110111011110;
#1 $display("%b", po);
# 1  pi=13'b1110111011111;
#1 $display("%b", po);
# 1  pi=13'b1110111100000;
#1 $display("%b", po);
# 1  pi=13'b1110111100001;
#1 $display("%b", po);
# 1  pi=13'b1110111100010;
#1 $display("%b", po);
# 1  pi=13'b1110111100011;
#1 $display("%b", po);
# 1  pi=13'b1110111100100;
#1 $display("%b", po);
# 1  pi=13'b1110111100101;
#1 $display("%b", po);
# 1  pi=13'b1110111100110;
#1 $display("%b", po);
# 1  pi=13'b1110111100111;
#1 $display("%b", po);
# 1  pi=13'b1110111101000;
#1 $display("%b", po);
# 1  pi=13'b1110111101001;
#1 $display("%b", po);
# 1  pi=13'b1110111101010;
#1 $display("%b", po);
# 1  pi=13'b1110111101011;
#1 $display("%b", po);
# 1  pi=13'b1110111101100;
#1 $display("%b", po);
# 1  pi=13'b1110111101101;
#1 $display("%b", po);
# 1  pi=13'b1110111101110;
#1 $display("%b", po);
# 1  pi=13'b1110111101111;
#1 $display("%b", po);
# 1  pi=13'b1110111110000;
#1 $display("%b", po);
# 1  pi=13'b1110111110001;
#1 $display("%b", po);
# 1  pi=13'b1110111110010;
#1 $display("%b", po);
# 1  pi=13'b1110111110011;
#1 $display("%b", po);
# 1  pi=13'b1110111110100;
#1 $display("%b", po);
# 1  pi=13'b1110111110101;
#1 $display("%b", po);
# 1  pi=13'b1110111110110;
#1 $display("%b", po);
# 1  pi=13'b1110111110111;
#1 $display("%b", po);
# 1  pi=13'b1110111111000;
#1 $display("%b", po);
# 1  pi=13'b1110111111001;
#1 $display("%b", po);
# 1  pi=13'b1110111111010;
#1 $display("%b", po);
# 1  pi=13'b1110111111011;
#1 $display("%b", po);
# 1  pi=13'b1110111111100;
#1 $display("%b", po);
# 1  pi=13'b1110111111101;
#1 $display("%b", po);
# 1  pi=13'b1110111111110;
#1 $display("%b", po);
# 1  pi=13'b1110111111111;
#1 $display("%b", po);
# 1  pi=13'b1111000000000;
#1 $display("%b", po);
# 1  pi=13'b1111000000001;
#1 $display("%b", po);
# 1  pi=13'b1111000000010;
#1 $display("%b", po);
# 1  pi=13'b1111000000011;
#1 $display("%b", po);
# 1  pi=13'b1111000000100;
#1 $display("%b", po);
# 1  pi=13'b1111000000101;
#1 $display("%b", po);
# 1  pi=13'b1111000000110;
#1 $display("%b", po);
# 1  pi=13'b1111000000111;
#1 $display("%b", po);
# 1  pi=13'b1111000001000;
#1 $display("%b", po);
# 1  pi=13'b1111000001001;
#1 $display("%b", po);
# 1  pi=13'b1111000001010;
#1 $display("%b", po);
# 1  pi=13'b1111000001011;
#1 $display("%b", po);
# 1  pi=13'b1111000001100;
#1 $display("%b", po);
# 1  pi=13'b1111000001101;
#1 $display("%b", po);
# 1  pi=13'b1111000001110;
#1 $display("%b", po);
# 1  pi=13'b1111000001111;
#1 $display("%b", po);
# 1  pi=13'b1111000010000;
#1 $display("%b", po);
# 1  pi=13'b1111000010001;
#1 $display("%b", po);
# 1  pi=13'b1111000010010;
#1 $display("%b", po);
# 1  pi=13'b1111000010011;
#1 $display("%b", po);
# 1  pi=13'b1111000010100;
#1 $display("%b", po);
# 1  pi=13'b1111000010101;
#1 $display("%b", po);
# 1  pi=13'b1111000010110;
#1 $display("%b", po);
# 1  pi=13'b1111000010111;
#1 $display("%b", po);
# 1  pi=13'b1111000011000;
#1 $display("%b", po);
# 1  pi=13'b1111000011001;
#1 $display("%b", po);
# 1  pi=13'b1111000011010;
#1 $display("%b", po);
# 1  pi=13'b1111000011011;
#1 $display("%b", po);
# 1  pi=13'b1111000011100;
#1 $display("%b", po);
# 1  pi=13'b1111000011101;
#1 $display("%b", po);
# 1  pi=13'b1111000011110;
#1 $display("%b", po);
# 1  pi=13'b1111000011111;
#1 $display("%b", po);
# 1  pi=13'b1111000100000;
#1 $display("%b", po);
# 1  pi=13'b1111000100001;
#1 $display("%b", po);
# 1  pi=13'b1111000100010;
#1 $display("%b", po);
# 1  pi=13'b1111000100011;
#1 $display("%b", po);
# 1  pi=13'b1111000100100;
#1 $display("%b", po);
# 1  pi=13'b1111000100101;
#1 $display("%b", po);
# 1  pi=13'b1111000100110;
#1 $display("%b", po);
# 1  pi=13'b1111000100111;
#1 $display("%b", po);
# 1  pi=13'b1111000101000;
#1 $display("%b", po);
# 1  pi=13'b1111000101001;
#1 $display("%b", po);
# 1  pi=13'b1111000101010;
#1 $display("%b", po);
# 1  pi=13'b1111000101011;
#1 $display("%b", po);
# 1  pi=13'b1111000101100;
#1 $display("%b", po);
# 1  pi=13'b1111000101101;
#1 $display("%b", po);
# 1  pi=13'b1111000101110;
#1 $display("%b", po);
# 1  pi=13'b1111000101111;
#1 $display("%b", po);
# 1  pi=13'b1111000110000;
#1 $display("%b", po);
# 1  pi=13'b1111000110001;
#1 $display("%b", po);
# 1  pi=13'b1111000110010;
#1 $display("%b", po);
# 1  pi=13'b1111000110011;
#1 $display("%b", po);
# 1  pi=13'b1111000110100;
#1 $display("%b", po);
# 1  pi=13'b1111000110101;
#1 $display("%b", po);
# 1  pi=13'b1111000110110;
#1 $display("%b", po);
# 1  pi=13'b1111000110111;
#1 $display("%b", po);
# 1  pi=13'b1111000111000;
#1 $display("%b", po);
# 1  pi=13'b1111000111001;
#1 $display("%b", po);
# 1  pi=13'b1111000111010;
#1 $display("%b", po);
# 1  pi=13'b1111000111011;
#1 $display("%b", po);
# 1  pi=13'b1111000111100;
#1 $display("%b", po);
# 1  pi=13'b1111000111101;
#1 $display("%b", po);
# 1  pi=13'b1111000111110;
#1 $display("%b", po);
# 1  pi=13'b1111000111111;
#1 $display("%b", po);
# 1  pi=13'b1111001000000;
#1 $display("%b", po);
# 1  pi=13'b1111001000001;
#1 $display("%b", po);
# 1  pi=13'b1111001000010;
#1 $display("%b", po);
# 1  pi=13'b1111001000011;
#1 $display("%b", po);
# 1  pi=13'b1111001000100;
#1 $display("%b", po);
# 1  pi=13'b1111001000101;
#1 $display("%b", po);
# 1  pi=13'b1111001000110;
#1 $display("%b", po);
# 1  pi=13'b1111001000111;
#1 $display("%b", po);
# 1  pi=13'b1111001001000;
#1 $display("%b", po);
# 1  pi=13'b1111001001001;
#1 $display("%b", po);
# 1  pi=13'b1111001001010;
#1 $display("%b", po);
# 1  pi=13'b1111001001011;
#1 $display("%b", po);
# 1  pi=13'b1111001001100;
#1 $display("%b", po);
# 1  pi=13'b1111001001101;
#1 $display("%b", po);
# 1  pi=13'b1111001001110;
#1 $display("%b", po);
# 1  pi=13'b1111001001111;
#1 $display("%b", po);
# 1  pi=13'b1111001010000;
#1 $display("%b", po);
# 1  pi=13'b1111001010001;
#1 $display("%b", po);
# 1  pi=13'b1111001010010;
#1 $display("%b", po);
# 1  pi=13'b1111001010011;
#1 $display("%b", po);
# 1  pi=13'b1111001010100;
#1 $display("%b", po);
# 1  pi=13'b1111001010101;
#1 $display("%b", po);
# 1  pi=13'b1111001010110;
#1 $display("%b", po);
# 1  pi=13'b1111001010111;
#1 $display("%b", po);
# 1  pi=13'b1111001011000;
#1 $display("%b", po);
# 1  pi=13'b1111001011001;
#1 $display("%b", po);
# 1  pi=13'b1111001011010;
#1 $display("%b", po);
# 1  pi=13'b1111001011011;
#1 $display("%b", po);
# 1  pi=13'b1111001011100;
#1 $display("%b", po);
# 1  pi=13'b1111001011101;
#1 $display("%b", po);
# 1  pi=13'b1111001011110;
#1 $display("%b", po);
# 1  pi=13'b1111001011111;
#1 $display("%b", po);
# 1  pi=13'b1111001100000;
#1 $display("%b", po);
# 1  pi=13'b1111001100001;
#1 $display("%b", po);
# 1  pi=13'b1111001100010;
#1 $display("%b", po);
# 1  pi=13'b1111001100011;
#1 $display("%b", po);
# 1  pi=13'b1111001100100;
#1 $display("%b", po);
# 1  pi=13'b1111001100101;
#1 $display("%b", po);
# 1  pi=13'b1111001100110;
#1 $display("%b", po);
# 1  pi=13'b1111001100111;
#1 $display("%b", po);
# 1  pi=13'b1111001101000;
#1 $display("%b", po);
# 1  pi=13'b1111001101001;
#1 $display("%b", po);
# 1  pi=13'b1111001101010;
#1 $display("%b", po);
# 1  pi=13'b1111001101011;
#1 $display("%b", po);
# 1  pi=13'b1111001101100;
#1 $display("%b", po);
# 1  pi=13'b1111001101101;
#1 $display("%b", po);
# 1  pi=13'b1111001101110;
#1 $display("%b", po);
# 1  pi=13'b1111001101111;
#1 $display("%b", po);
# 1  pi=13'b1111001110000;
#1 $display("%b", po);
# 1  pi=13'b1111001110001;
#1 $display("%b", po);
# 1  pi=13'b1111001110010;
#1 $display("%b", po);
# 1  pi=13'b1111001110011;
#1 $display("%b", po);
# 1  pi=13'b1111001110100;
#1 $display("%b", po);
# 1  pi=13'b1111001110101;
#1 $display("%b", po);
# 1  pi=13'b1111001110110;
#1 $display("%b", po);
# 1  pi=13'b1111001110111;
#1 $display("%b", po);
# 1  pi=13'b1111001111000;
#1 $display("%b", po);
# 1  pi=13'b1111001111001;
#1 $display("%b", po);
# 1  pi=13'b1111001111010;
#1 $display("%b", po);
# 1  pi=13'b1111001111011;
#1 $display("%b", po);
# 1  pi=13'b1111001111100;
#1 $display("%b", po);
# 1  pi=13'b1111001111101;
#1 $display("%b", po);
# 1  pi=13'b1111001111110;
#1 $display("%b", po);
# 1  pi=13'b1111001111111;
#1 $display("%b", po);
# 1  pi=13'b1111010000000;
#1 $display("%b", po);
# 1  pi=13'b1111010000001;
#1 $display("%b", po);
# 1  pi=13'b1111010000010;
#1 $display("%b", po);
# 1  pi=13'b1111010000011;
#1 $display("%b", po);
# 1  pi=13'b1111010000100;
#1 $display("%b", po);
# 1  pi=13'b1111010000101;
#1 $display("%b", po);
# 1  pi=13'b1111010000110;
#1 $display("%b", po);
# 1  pi=13'b1111010000111;
#1 $display("%b", po);
# 1  pi=13'b1111010001000;
#1 $display("%b", po);
# 1  pi=13'b1111010001001;
#1 $display("%b", po);
# 1  pi=13'b1111010001010;
#1 $display("%b", po);
# 1  pi=13'b1111010001011;
#1 $display("%b", po);
# 1  pi=13'b1111010001100;
#1 $display("%b", po);
# 1  pi=13'b1111010001101;
#1 $display("%b", po);
# 1  pi=13'b1111010001110;
#1 $display("%b", po);
# 1  pi=13'b1111010001111;
#1 $display("%b", po);
# 1  pi=13'b1111010010000;
#1 $display("%b", po);
# 1  pi=13'b1111010010001;
#1 $display("%b", po);
# 1  pi=13'b1111010010010;
#1 $display("%b", po);
# 1  pi=13'b1111010010011;
#1 $display("%b", po);
# 1  pi=13'b1111010010100;
#1 $display("%b", po);
# 1  pi=13'b1111010010101;
#1 $display("%b", po);
# 1  pi=13'b1111010010110;
#1 $display("%b", po);
# 1  pi=13'b1111010010111;
#1 $display("%b", po);
# 1  pi=13'b1111010011000;
#1 $display("%b", po);
# 1  pi=13'b1111010011001;
#1 $display("%b", po);
# 1  pi=13'b1111010011010;
#1 $display("%b", po);
# 1  pi=13'b1111010011011;
#1 $display("%b", po);
# 1  pi=13'b1111010011100;
#1 $display("%b", po);
# 1  pi=13'b1111010011101;
#1 $display("%b", po);
# 1  pi=13'b1111010011110;
#1 $display("%b", po);
# 1  pi=13'b1111010011111;
#1 $display("%b", po);
# 1  pi=13'b1111010100000;
#1 $display("%b", po);
# 1  pi=13'b1111010100001;
#1 $display("%b", po);
# 1  pi=13'b1111010100010;
#1 $display("%b", po);
# 1  pi=13'b1111010100011;
#1 $display("%b", po);
# 1  pi=13'b1111010100100;
#1 $display("%b", po);
# 1  pi=13'b1111010100101;
#1 $display("%b", po);
# 1  pi=13'b1111010100110;
#1 $display("%b", po);
# 1  pi=13'b1111010100111;
#1 $display("%b", po);
# 1  pi=13'b1111010101000;
#1 $display("%b", po);
# 1  pi=13'b1111010101001;
#1 $display("%b", po);
# 1  pi=13'b1111010101010;
#1 $display("%b", po);
# 1  pi=13'b1111010101011;
#1 $display("%b", po);
# 1  pi=13'b1111010101100;
#1 $display("%b", po);
# 1  pi=13'b1111010101101;
#1 $display("%b", po);
# 1  pi=13'b1111010101110;
#1 $display("%b", po);
# 1  pi=13'b1111010101111;
#1 $display("%b", po);
# 1  pi=13'b1111010110000;
#1 $display("%b", po);
# 1  pi=13'b1111010110001;
#1 $display("%b", po);
# 1  pi=13'b1111010110010;
#1 $display("%b", po);
# 1  pi=13'b1111010110011;
#1 $display("%b", po);
# 1  pi=13'b1111010110100;
#1 $display("%b", po);
# 1  pi=13'b1111010110101;
#1 $display("%b", po);
# 1  pi=13'b1111010110110;
#1 $display("%b", po);
# 1  pi=13'b1111010110111;
#1 $display("%b", po);
# 1  pi=13'b1111010111000;
#1 $display("%b", po);
# 1  pi=13'b1111010111001;
#1 $display("%b", po);
# 1  pi=13'b1111010111010;
#1 $display("%b", po);
# 1  pi=13'b1111010111011;
#1 $display("%b", po);
# 1  pi=13'b1111010111100;
#1 $display("%b", po);
# 1  pi=13'b1111010111101;
#1 $display("%b", po);
# 1  pi=13'b1111010111110;
#1 $display("%b", po);
# 1  pi=13'b1111010111111;
#1 $display("%b", po);
# 1  pi=13'b1111011000000;
#1 $display("%b", po);
# 1  pi=13'b1111011000001;
#1 $display("%b", po);
# 1  pi=13'b1111011000010;
#1 $display("%b", po);
# 1  pi=13'b1111011000011;
#1 $display("%b", po);
# 1  pi=13'b1111011000100;
#1 $display("%b", po);
# 1  pi=13'b1111011000101;
#1 $display("%b", po);
# 1  pi=13'b1111011000110;
#1 $display("%b", po);
# 1  pi=13'b1111011000111;
#1 $display("%b", po);
# 1  pi=13'b1111011001000;
#1 $display("%b", po);
# 1  pi=13'b1111011001001;
#1 $display("%b", po);
# 1  pi=13'b1111011001010;
#1 $display("%b", po);
# 1  pi=13'b1111011001011;
#1 $display("%b", po);
# 1  pi=13'b1111011001100;
#1 $display("%b", po);
# 1  pi=13'b1111011001101;
#1 $display("%b", po);
# 1  pi=13'b1111011001110;
#1 $display("%b", po);
# 1  pi=13'b1111011001111;
#1 $display("%b", po);
# 1  pi=13'b1111011010000;
#1 $display("%b", po);
# 1  pi=13'b1111011010001;
#1 $display("%b", po);
# 1  pi=13'b1111011010010;
#1 $display("%b", po);
# 1  pi=13'b1111011010011;
#1 $display("%b", po);
# 1  pi=13'b1111011010100;
#1 $display("%b", po);
# 1  pi=13'b1111011010101;
#1 $display("%b", po);
# 1  pi=13'b1111011010110;
#1 $display("%b", po);
# 1  pi=13'b1111011010111;
#1 $display("%b", po);
# 1  pi=13'b1111011011000;
#1 $display("%b", po);
# 1  pi=13'b1111011011001;
#1 $display("%b", po);
# 1  pi=13'b1111011011010;
#1 $display("%b", po);
# 1  pi=13'b1111011011011;
#1 $display("%b", po);
# 1  pi=13'b1111011011100;
#1 $display("%b", po);
# 1  pi=13'b1111011011101;
#1 $display("%b", po);
# 1  pi=13'b1111011011110;
#1 $display("%b", po);
# 1  pi=13'b1111011011111;
#1 $display("%b", po);
# 1  pi=13'b1111011100000;
#1 $display("%b", po);
# 1  pi=13'b1111011100001;
#1 $display("%b", po);
# 1  pi=13'b1111011100010;
#1 $display("%b", po);
# 1  pi=13'b1111011100011;
#1 $display("%b", po);
# 1  pi=13'b1111011100100;
#1 $display("%b", po);
# 1  pi=13'b1111011100101;
#1 $display("%b", po);
# 1  pi=13'b1111011100110;
#1 $display("%b", po);
# 1  pi=13'b1111011100111;
#1 $display("%b", po);
# 1  pi=13'b1111011101000;
#1 $display("%b", po);
# 1  pi=13'b1111011101001;
#1 $display("%b", po);
# 1  pi=13'b1111011101010;
#1 $display("%b", po);
# 1  pi=13'b1111011101011;
#1 $display("%b", po);
# 1  pi=13'b1111011101100;
#1 $display("%b", po);
# 1  pi=13'b1111011101101;
#1 $display("%b", po);
# 1  pi=13'b1111011101110;
#1 $display("%b", po);
# 1  pi=13'b1111011101111;
#1 $display("%b", po);
# 1  pi=13'b1111011110000;
#1 $display("%b", po);
# 1  pi=13'b1111011110001;
#1 $display("%b", po);
# 1  pi=13'b1111011110010;
#1 $display("%b", po);
# 1  pi=13'b1111011110011;
#1 $display("%b", po);
# 1  pi=13'b1111011110100;
#1 $display("%b", po);
# 1  pi=13'b1111011110101;
#1 $display("%b", po);
# 1  pi=13'b1111011110110;
#1 $display("%b", po);
# 1  pi=13'b1111011110111;
#1 $display("%b", po);
# 1  pi=13'b1111011111000;
#1 $display("%b", po);
# 1  pi=13'b1111011111001;
#1 $display("%b", po);
# 1  pi=13'b1111011111010;
#1 $display("%b", po);
# 1  pi=13'b1111011111011;
#1 $display("%b", po);
# 1  pi=13'b1111011111100;
#1 $display("%b", po);
# 1  pi=13'b1111011111101;
#1 $display("%b", po);
# 1  pi=13'b1111011111110;
#1 $display("%b", po);
# 1  pi=13'b1111011111111;
#1 $display("%b", po);
# 1  pi=13'b1111100000000;
#1 $display("%b", po);
# 1  pi=13'b1111100000001;
#1 $display("%b", po);
# 1  pi=13'b1111100000010;
#1 $display("%b", po);
# 1  pi=13'b1111100000011;
#1 $display("%b", po);
# 1  pi=13'b1111100000100;
#1 $display("%b", po);
# 1  pi=13'b1111100000101;
#1 $display("%b", po);
# 1  pi=13'b1111100000110;
#1 $display("%b", po);
# 1  pi=13'b1111100000111;
#1 $display("%b", po);
# 1  pi=13'b1111100001000;
#1 $display("%b", po);
# 1  pi=13'b1111100001001;
#1 $display("%b", po);
# 1  pi=13'b1111100001010;
#1 $display("%b", po);
# 1  pi=13'b1111100001011;
#1 $display("%b", po);
# 1  pi=13'b1111100001100;
#1 $display("%b", po);
# 1  pi=13'b1111100001101;
#1 $display("%b", po);
# 1  pi=13'b1111100001110;
#1 $display("%b", po);
# 1  pi=13'b1111100001111;
#1 $display("%b", po);
# 1  pi=13'b1111100010000;
#1 $display("%b", po);
# 1  pi=13'b1111100010001;
#1 $display("%b", po);
# 1  pi=13'b1111100010010;
#1 $display("%b", po);
# 1  pi=13'b1111100010011;
#1 $display("%b", po);
# 1  pi=13'b1111100010100;
#1 $display("%b", po);
# 1  pi=13'b1111100010101;
#1 $display("%b", po);
# 1  pi=13'b1111100010110;
#1 $display("%b", po);
# 1  pi=13'b1111100010111;
#1 $display("%b", po);
# 1  pi=13'b1111100011000;
#1 $display("%b", po);
# 1  pi=13'b1111100011001;
#1 $display("%b", po);
# 1  pi=13'b1111100011010;
#1 $display("%b", po);
# 1  pi=13'b1111100011011;
#1 $display("%b", po);
# 1  pi=13'b1111100011100;
#1 $display("%b", po);
# 1  pi=13'b1111100011101;
#1 $display("%b", po);
# 1  pi=13'b1111100011110;
#1 $display("%b", po);
# 1  pi=13'b1111100011111;
#1 $display("%b", po);
# 1  pi=13'b1111100100000;
#1 $display("%b", po);
# 1  pi=13'b1111100100001;
#1 $display("%b", po);
# 1  pi=13'b1111100100010;
#1 $display("%b", po);
# 1  pi=13'b1111100100011;
#1 $display("%b", po);
# 1  pi=13'b1111100100100;
#1 $display("%b", po);
# 1  pi=13'b1111100100101;
#1 $display("%b", po);
# 1  pi=13'b1111100100110;
#1 $display("%b", po);
# 1  pi=13'b1111100100111;
#1 $display("%b", po);
# 1  pi=13'b1111100101000;
#1 $display("%b", po);
# 1  pi=13'b1111100101001;
#1 $display("%b", po);
# 1  pi=13'b1111100101010;
#1 $display("%b", po);
# 1  pi=13'b1111100101011;
#1 $display("%b", po);
# 1  pi=13'b1111100101100;
#1 $display("%b", po);
# 1  pi=13'b1111100101101;
#1 $display("%b", po);
# 1  pi=13'b1111100101110;
#1 $display("%b", po);
# 1  pi=13'b1111100101111;
#1 $display("%b", po);
# 1  pi=13'b1111100110000;
#1 $display("%b", po);
# 1  pi=13'b1111100110001;
#1 $display("%b", po);
# 1  pi=13'b1111100110010;
#1 $display("%b", po);
# 1  pi=13'b1111100110011;
#1 $display("%b", po);
# 1  pi=13'b1111100110100;
#1 $display("%b", po);
# 1  pi=13'b1111100110101;
#1 $display("%b", po);
# 1  pi=13'b1111100110110;
#1 $display("%b", po);
# 1  pi=13'b1111100110111;
#1 $display("%b", po);
# 1  pi=13'b1111100111000;
#1 $display("%b", po);
# 1  pi=13'b1111100111001;
#1 $display("%b", po);
# 1  pi=13'b1111100111010;
#1 $display("%b", po);
# 1  pi=13'b1111100111011;
#1 $display("%b", po);
# 1  pi=13'b1111100111100;
#1 $display("%b", po);
# 1  pi=13'b1111100111101;
#1 $display("%b", po);
# 1  pi=13'b1111100111110;
#1 $display("%b", po);
# 1  pi=13'b1111100111111;
#1 $display("%b", po);
# 1  pi=13'b1111101000000;
#1 $display("%b", po);
# 1  pi=13'b1111101000001;
#1 $display("%b", po);
# 1  pi=13'b1111101000010;
#1 $display("%b", po);
# 1  pi=13'b1111101000011;
#1 $display("%b", po);
# 1  pi=13'b1111101000100;
#1 $display("%b", po);
# 1  pi=13'b1111101000101;
#1 $display("%b", po);
# 1  pi=13'b1111101000110;
#1 $display("%b", po);
# 1  pi=13'b1111101000111;
#1 $display("%b", po);
# 1  pi=13'b1111101001000;
#1 $display("%b", po);
# 1  pi=13'b1111101001001;
#1 $display("%b", po);
# 1  pi=13'b1111101001010;
#1 $display("%b", po);
# 1  pi=13'b1111101001011;
#1 $display("%b", po);
# 1  pi=13'b1111101001100;
#1 $display("%b", po);
# 1  pi=13'b1111101001101;
#1 $display("%b", po);
# 1  pi=13'b1111101001110;
#1 $display("%b", po);
# 1  pi=13'b1111101001111;
#1 $display("%b", po);
# 1  pi=13'b1111101010000;
#1 $display("%b", po);
# 1  pi=13'b1111101010001;
#1 $display("%b", po);
# 1  pi=13'b1111101010010;
#1 $display("%b", po);
# 1  pi=13'b1111101010011;
#1 $display("%b", po);
# 1  pi=13'b1111101010100;
#1 $display("%b", po);
# 1  pi=13'b1111101010101;
#1 $display("%b", po);
# 1  pi=13'b1111101010110;
#1 $display("%b", po);
# 1  pi=13'b1111101010111;
#1 $display("%b", po);
# 1  pi=13'b1111101011000;
#1 $display("%b", po);
# 1  pi=13'b1111101011001;
#1 $display("%b", po);
# 1  pi=13'b1111101011010;
#1 $display("%b", po);
# 1  pi=13'b1111101011011;
#1 $display("%b", po);
# 1  pi=13'b1111101011100;
#1 $display("%b", po);
# 1  pi=13'b1111101011101;
#1 $display("%b", po);
# 1  pi=13'b1111101011110;
#1 $display("%b", po);
# 1  pi=13'b1111101011111;
#1 $display("%b", po);
# 1  pi=13'b1111101100000;
#1 $display("%b", po);
# 1  pi=13'b1111101100001;
#1 $display("%b", po);
# 1  pi=13'b1111101100010;
#1 $display("%b", po);
# 1  pi=13'b1111101100011;
#1 $display("%b", po);
# 1  pi=13'b1111101100100;
#1 $display("%b", po);
# 1  pi=13'b1111101100101;
#1 $display("%b", po);
# 1  pi=13'b1111101100110;
#1 $display("%b", po);
# 1  pi=13'b1111101100111;
#1 $display("%b", po);
# 1  pi=13'b1111101101000;
#1 $display("%b", po);
# 1  pi=13'b1111101101001;
#1 $display("%b", po);
# 1  pi=13'b1111101101010;
#1 $display("%b", po);
# 1  pi=13'b1111101101011;
#1 $display("%b", po);
# 1  pi=13'b1111101101100;
#1 $display("%b", po);
# 1  pi=13'b1111101101101;
#1 $display("%b", po);
# 1  pi=13'b1111101101110;
#1 $display("%b", po);
# 1  pi=13'b1111101101111;
#1 $display("%b", po);
# 1  pi=13'b1111101110000;
#1 $display("%b", po);
# 1  pi=13'b1111101110001;
#1 $display("%b", po);
# 1  pi=13'b1111101110010;
#1 $display("%b", po);
# 1  pi=13'b1111101110011;
#1 $display("%b", po);
# 1  pi=13'b1111101110100;
#1 $display("%b", po);
# 1  pi=13'b1111101110101;
#1 $display("%b", po);
# 1  pi=13'b1111101110110;
#1 $display("%b", po);
# 1  pi=13'b1111101110111;
#1 $display("%b", po);
# 1  pi=13'b1111101111000;
#1 $display("%b", po);
# 1  pi=13'b1111101111001;
#1 $display("%b", po);
# 1  pi=13'b1111101111010;
#1 $display("%b", po);
# 1  pi=13'b1111101111011;
#1 $display("%b", po);
# 1  pi=13'b1111101111100;
#1 $display("%b", po);
# 1  pi=13'b1111101111101;
#1 $display("%b", po);
# 1  pi=13'b1111101111110;
#1 $display("%b", po);
# 1  pi=13'b1111101111111;
#1 $display("%b", po);
# 1  pi=13'b1111110000000;
#1 $display("%b", po);
# 1  pi=13'b1111110000001;
#1 $display("%b", po);
# 1  pi=13'b1111110000010;
#1 $display("%b", po);
# 1  pi=13'b1111110000011;
#1 $display("%b", po);
# 1  pi=13'b1111110000100;
#1 $display("%b", po);
# 1  pi=13'b1111110000101;
#1 $display("%b", po);
# 1  pi=13'b1111110000110;
#1 $display("%b", po);
# 1  pi=13'b1111110000111;
#1 $display("%b", po);
# 1  pi=13'b1111110001000;
#1 $display("%b", po);
# 1  pi=13'b1111110001001;
#1 $display("%b", po);
# 1  pi=13'b1111110001010;
#1 $display("%b", po);
# 1  pi=13'b1111110001011;
#1 $display("%b", po);
# 1  pi=13'b1111110001100;
#1 $display("%b", po);
# 1  pi=13'b1111110001101;
#1 $display("%b", po);
# 1  pi=13'b1111110001110;
#1 $display("%b", po);
# 1  pi=13'b1111110001111;
#1 $display("%b", po);
# 1  pi=13'b1111110010000;
#1 $display("%b", po);
# 1  pi=13'b1111110010001;
#1 $display("%b", po);
# 1  pi=13'b1111110010010;
#1 $display("%b", po);
# 1  pi=13'b1111110010011;
#1 $display("%b", po);
# 1  pi=13'b1111110010100;
#1 $display("%b", po);
# 1  pi=13'b1111110010101;
#1 $display("%b", po);
# 1  pi=13'b1111110010110;
#1 $display("%b", po);
# 1  pi=13'b1111110010111;
#1 $display("%b", po);
# 1  pi=13'b1111110011000;
#1 $display("%b", po);
# 1  pi=13'b1111110011001;
#1 $display("%b", po);
# 1  pi=13'b1111110011010;
#1 $display("%b", po);
# 1  pi=13'b1111110011011;
#1 $display("%b", po);
# 1  pi=13'b1111110011100;
#1 $display("%b", po);
# 1  pi=13'b1111110011101;
#1 $display("%b", po);
# 1  pi=13'b1111110011110;
#1 $display("%b", po);
# 1  pi=13'b1111110011111;
#1 $display("%b", po);
# 1  pi=13'b1111110100000;
#1 $display("%b", po);
# 1  pi=13'b1111110100001;
#1 $display("%b", po);
# 1  pi=13'b1111110100010;
#1 $display("%b", po);
# 1  pi=13'b1111110100011;
#1 $display("%b", po);
# 1  pi=13'b1111110100100;
#1 $display("%b", po);
# 1  pi=13'b1111110100101;
#1 $display("%b", po);
# 1  pi=13'b1111110100110;
#1 $display("%b", po);
# 1  pi=13'b1111110100111;
#1 $display("%b", po);
# 1  pi=13'b1111110101000;
#1 $display("%b", po);
# 1  pi=13'b1111110101001;
#1 $display("%b", po);
# 1  pi=13'b1111110101010;
#1 $display("%b", po);
# 1  pi=13'b1111110101011;
#1 $display("%b", po);
# 1  pi=13'b1111110101100;
#1 $display("%b", po);
# 1  pi=13'b1111110101101;
#1 $display("%b", po);
# 1  pi=13'b1111110101110;
#1 $display("%b", po);
# 1  pi=13'b1111110101111;
#1 $display("%b", po);
# 1  pi=13'b1111110110000;
#1 $display("%b", po);
# 1  pi=13'b1111110110001;
#1 $display("%b", po);
# 1  pi=13'b1111110110010;
#1 $display("%b", po);
# 1  pi=13'b1111110110011;
#1 $display("%b", po);
# 1  pi=13'b1111110110100;
#1 $display("%b", po);
# 1  pi=13'b1111110110101;
#1 $display("%b", po);
# 1  pi=13'b1111110110110;
#1 $display("%b", po);
# 1  pi=13'b1111110110111;
#1 $display("%b", po);
# 1  pi=13'b1111110111000;
#1 $display("%b", po);
# 1  pi=13'b1111110111001;
#1 $display("%b", po);
# 1  pi=13'b1111110111010;
#1 $display("%b", po);
# 1  pi=13'b1111110111011;
#1 $display("%b", po);
# 1  pi=13'b1111110111100;
#1 $display("%b", po);
# 1  pi=13'b1111110111101;
#1 $display("%b", po);
# 1  pi=13'b1111110111110;
#1 $display("%b", po);
# 1  pi=13'b1111110111111;
#1 $display("%b", po);
# 1  pi=13'b1111111000000;
#1 $display("%b", po);
# 1  pi=13'b1111111000001;
#1 $display("%b", po);
# 1  pi=13'b1111111000010;
#1 $display("%b", po);
# 1  pi=13'b1111111000011;
#1 $display("%b", po);
# 1  pi=13'b1111111000100;
#1 $display("%b", po);
# 1  pi=13'b1111111000101;
#1 $display("%b", po);
# 1  pi=13'b1111111000110;
#1 $display("%b", po);
# 1  pi=13'b1111111000111;
#1 $display("%b", po);
# 1  pi=13'b1111111001000;
#1 $display("%b", po);
# 1  pi=13'b1111111001001;
#1 $display("%b", po);
# 1  pi=13'b1111111001010;
#1 $display("%b", po);
# 1  pi=13'b1111111001011;
#1 $display("%b", po);
# 1  pi=13'b1111111001100;
#1 $display("%b", po);
# 1  pi=13'b1111111001101;
#1 $display("%b", po);
# 1  pi=13'b1111111001110;
#1 $display("%b", po);
# 1  pi=13'b1111111001111;
#1 $display("%b", po);
# 1  pi=13'b1111111010000;
#1 $display("%b", po);
# 1  pi=13'b1111111010001;
#1 $display("%b", po);
# 1  pi=13'b1111111010010;
#1 $display("%b", po);
# 1  pi=13'b1111111010011;
#1 $display("%b", po);
# 1  pi=13'b1111111010100;
#1 $display("%b", po);
# 1  pi=13'b1111111010101;
#1 $display("%b", po);
# 1  pi=13'b1111111010110;
#1 $display("%b", po);
# 1  pi=13'b1111111010111;
#1 $display("%b", po);
# 1  pi=13'b1111111011000;
#1 $display("%b", po);
# 1  pi=13'b1111111011001;
#1 $display("%b", po);
# 1  pi=13'b1111111011010;
#1 $display("%b", po);
# 1  pi=13'b1111111011011;
#1 $display("%b", po);
# 1  pi=13'b1111111011100;
#1 $display("%b", po);
# 1  pi=13'b1111111011101;
#1 $display("%b", po);
# 1  pi=13'b1111111011110;
#1 $display("%b", po);
# 1  pi=13'b1111111011111;
#1 $display("%b", po);
# 1  pi=13'b1111111100000;
#1 $display("%b", po);
# 1  pi=13'b1111111100001;
#1 $display("%b", po);
# 1  pi=13'b1111111100010;
#1 $display("%b", po);
# 1  pi=13'b1111111100011;
#1 $display("%b", po);
# 1  pi=13'b1111111100100;
#1 $display("%b", po);
# 1  pi=13'b1111111100101;
#1 $display("%b", po);
# 1  pi=13'b1111111100110;
#1 $display("%b", po);
# 1  pi=13'b1111111100111;
#1 $display("%b", po);
# 1  pi=13'b1111111101000;
#1 $display("%b", po);
# 1  pi=13'b1111111101001;
#1 $display("%b", po);
# 1  pi=13'b1111111101010;
#1 $display("%b", po);
# 1  pi=13'b1111111101011;
#1 $display("%b", po);
# 1  pi=13'b1111111101100;
#1 $display("%b", po);
# 1  pi=13'b1111111101101;
#1 $display("%b", po);
# 1  pi=13'b1111111101110;
#1 $display("%b", po);
# 1  pi=13'b1111111101111;
#1 $display("%b", po);
# 1  pi=13'b1111111110000;
#1 $display("%b", po);
# 1  pi=13'b1111111110001;
#1 $display("%b", po);
# 1  pi=13'b1111111110010;
#1 $display("%b", po);
# 1  pi=13'b1111111110011;
#1 $display("%b", po);
# 1  pi=13'b1111111110100;
#1 $display("%b", po);
# 1  pi=13'b1111111110101;
#1 $display("%b", po);
# 1  pi=13'b1111111110110;
#1 $display("%b", po);
# 1  pi=13'b1111111110111;
#1 $display("%b", po);
# 1  pi=13'b1111111111000;
#1 $display("%b", po);
# 1  pi=13'b1111111111001;
#1 $display("%b", po);
# 1  pi=13'b1111111111010;
#1 $display("%b", po);
# 1  pi=13'b1111111111011;
#1 $display("%b", po);
# 1  pi=13'b1111111111100;
#1 $display("%b", po);
# 1  pi=13'b1111111111101;
#1 $display("%b", po);
# 1  pi=13'b1111111111110;
#1 $display("%b", po);
# 1  pi=13'b1111111111111;
#1 $display("%b", po);
end
endmodule
