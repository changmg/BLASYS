module adder_1(pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 , pi11 , po0 , po1 , po2 , po3 , po4 , po5 , po6 );
  input pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 , pi11 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 ;
  wire new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36, new_n37, new_n38, new_n39, new_n40, new_n41, new_n42, new_n43, new_n44, new_n45, new_n46, new_n47, new_n48, new_n49, new_n50, new_n51, new_n52, new_n53, new_n54, new_n55, new_n56, new_n57, new_n58, new_n59, new_n60, new_n61, new_n62;
  assign new_n13 = pi00 & pi05 ;
  assign new_n14 = ~pi00 & ~pi05 ;
  assign new_n15 = ~new_n13 & ~new_n14 ;
  assign new_n16 = ~pi10 & ~new_n15 ;
  assign new_n17 = ~pi11 & new_n15 ;
  assign new_n18 = ~new_n16 & ~new_n17 ;
  assign new_n19 = ~pi10 & ~new_n14 ;
  assign new_n20 = ~new_n13 & ~new_n19 ;
  assign new_n21 = pi06 & ~new_n20 ;
  assign new_n22 = ~pi11 & ~new_n13 ;
  assign new_n23 = ~new_n14 & ~new_n22 ;
  assign new_n24 = ~pi06 & ~new_n23 ;
  assign new_n25 = ~new_n21 & ~new_n24 ;
  assign new_n26 = pi01 & ~new_n25 ;
  assign new_n27 = ~pi01 & new_n25 ;
  assign new_n28 = ~new_n26 & ~new_n27 ;
  assign new_n29 = pi02 & pi07 ;
  assign new_n30 = ~pi02 & ~pi07 ;
  assign new_n31 = ~new_n29 & ~new_n30 ;
  assign new_n32 = pi01 & ~new_n24 ;
  assign new_n33 = ~new_n21 & ~new_n32 ;
  assign new_n34 = ~new_n31 & ~new_n33 ;
  assign new_n35 = ~pi01 & ~new_n21 ;
  assign new_n36 = ~new_n24 & ~new_n35 ;
  assign new_n37 = new_n31 & ~new_n36 ;
  assign new_n38 = ~new_n34 & ~new_n37 ;
  assign new_n39 = ~new_n30 & ~new_n33 ;
  assign new_n40 = ~new_n29 & ~new_n39 ;
  assign new_n41 = pi08 & ~new_n40 ;
  assign new_n42 = ~new_n29 & ~new_n36 ;
  assign new_n43 = ~new_n30 & ~new_n42 ;
  assign new_n44 = ~pi08 & ~new_n43 ;
  assign new_n45 = ~new_n41 & ~new_n44 ;
  assign new_n46 = pi03 & ~new_n45 ;
  assign new_n47 = ~pi03 & new_n45 ;
  assign new_n48 = ~new_n46 & ~new_n47 ;
  assign new_n49 = pi03 & ~new_n44 ;
  assign new_n50 = ~new_n41 & ~new_n49 ;
  assign new_n51 = ~pi04 & ~pi09 ;
  assign new_n52 = pi04 & pi09 ;
  assign new_n53 = ~new_n51 & ~new_n52 ;
  assign new_n54 = ~new_n50 & ~new_n53 ;
  assign new_n55 = ~pi03 & ~new_n41 ;
  assign new_n56 = ~new_n44 & ~new_n55 ;
  assign new_n57 = new_n53 & ~new_n56 ;
  assign new_n58 = ~new_n54 & ~new_n57 ;
  assign new_n59 = ~new_n50 & ~new_n51 ;
  assign new_n60 = ~new_n52 & ~new_n59 ;
  assign new_n61 = ~new_n52 & ~new_n56 ;
  assign new_n62 = ~new_n51 & ~new_n61 ;
  assign po0 = new_n18 ;
  assign po1 = new_n28 ;
  assign po2 = new_n38 ;
  assign po3 = new_n48 ;
  assign po4 = new_n58 ;
  assign po5 = new_n60 ;
  assign po6 = new_n62 ;
endmodule
