// Benchmark "mult16" written by ABC on Fri Jul  1 13:52:02 2022

module mult16 ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ,
    \r[0] , \r[1] , \r[2] , \r[3] , \r[4] , \r[5] , \r[6] , \r[7] , \r[8] ,
    \r[9] , \r[10] , \r[11] , \r[12] , \r[13] , \r[14] , \r[15] , \r[16] ,
    \r[17] , \r[18] , \r[19] , \r[20] , \r[21] , \r[22] , \r[23] , \r[24] ,
    \r[25] , \r[26] , \r[27] , \r[28] , \r[29] , \r[30] , \r[31]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] ;
  output \r[0] , \r[1] , \r[2] , \r[3] , \r[4] , \r[5] , \r[6] , \r[7] ,
    \r[8] , \r[9] , \r[10] , \r[11] , \r[12] , \r[13] , \r[14] , \r[15] ,
    \r[16] , \r[17] , \r[18] , \r[19] , \r[20] , \r[21] , \r[22] , \r[23] ,
    \r[24] , \r[25] , \r[26] , \r[27] , \r[28] , \r[29] , \r[30] , \r[31] ;
  wire new_new_n66__, new_new_n67__, new_new_n68__, new_new_n69__,
    new_new_n71__, new_new_n72__, new_new_n73__, new_new_n74__,
    new_new_n75__, new_new_n76__, new_new_n77__, new_new_n78__,
    new_new_n79__, new_new_n80__, new_new_n81__, new_new_n83__,
    new_new_n84__, new_new_n85__, new_new_n86__, new_new_n87__,
    new_new_n88__, new_new_n89__, new_new_n90__, new_new_n91__,
    new_new_n92__, new_new_n93__, new_new_n94__, new_new_n95__,
    new_new_n96__, new_new_n97__, new_new_n98__, new_new_n99__,
    new_new_n101__, new_new_n102__, new_new_n103__, new_new_n104__,
    new_new_n105__, new_new_n106__, new_new_n107__, new_new_n108__,
    new_new_n109__, new_new_n110__, new_new_n111__, new_new_n112__,
    new_new_n113__, new_new_n114__, new_new_n115__, new_new_n116__,
    new_new_n117__, new_new_n118__, new_new_n119__, new_new_n120__,
    new_new_n121__, new_new_n122__, new_new_n123__, new_new_n124__,
    new_new_n125__, new_new_n126__, new_new_n127__, new_new_n128__,
    new_new_n129__, new_new_n131__, new_new_n132__, new_new_n133__,
    new_new_n134__, new_new_n135__, new_new_n136__, new_new_n137__,
    new_new_n138__, new_new_n139__, new_new_n140__, new_new_n141__,
    new_new_n142__, new_new_n143__, new_new_n144__, new_new_n145__,
    new_new_n146__, new_new_n147__, new_new_n148__, new_new_n149__,
    new_new_n150__, new_new_n151__, new_new_n152__, new_new_n153__,
    new_new_n154__, new_new_n155__, new_new_n156__, new_new_n157__,
    new_new_n158__, new_new_n159__, new_new_n160__, new_new_n161__,
    new_new_n162__, new_new_n163__, new_new_n164__, new_new_n165__,
    new_new_n167__, new_new_n168__, new_new_n169__, new_new_n170__,
    new_new_n171__, new_new_n172__, new_new_n173__, new_new_n174__,
    new_new_n175__, new_new_n176__, new_new_n177__, new_new_n178__,
    new_new_n179__, new_new_n180__, new_new_n181__, new_new_n182__,
    new_new_n183__, new_new_n184__, new_new_n185__, new_new_n186__,
    new_new_n187__, new_new_n188__, new_new_n189__, new_new_n190__,
    new_new_n191__, new_new_n192__, new_new_n193__, new_new_n194__,
    new_new_n195__, new_new_n196__, new_new_n197__, new_new_n198__,
    new_new_n199__, new_new_n200__, new_new_n201__, new_new_n202__,
    new_new_n203__, new_new_n204__, new_new_n205__, new_new_n206__,
    new_new_n207__, new_new_n208__, new_new_n209__, new_new_n210__,
    new_new_n211__, new_new_n212__, new_new_n213__, new_new_n214__,
    new_new_n216__, new_new_n217__, new_new_n218__, new_new_n219__,
    new_new_n220__, new_new_n221__, new_new_n222__, new_new_n223__,
    new_new_n224__, new_new_n225__, new_new_n226__, new_new_n227__,
    new_new_n228__, new_new_n229__, new_new_n230__, new_new_n231__,
    new_new_n232__, new_new_n233__, new_new_n234__, new_new_n235__,
    new_new_n236__, new_new_n237__, new_new_n238__, new_new_n239__,
    new_new_n240__, new_new_n241__, new_new_n242__, new_new_n243__,
    new_new_n244__, new_new_n245__, new_new_n246__, new_new_n247__,
    new_new_n248__, new_new_n249__, new_new_n250__, new_new_n251__,
    new_new_n252__, new_new_n253__, new_new_n254__, new_new_n255__,
    new_new_n256__, new_new_n257__, new_new_n258__, new_new_n259__,
    new_new_n260__, new_new_n261__, new_new_n262__, new_new_n263__,
    new_new_n264__, new_new_n265__, new_new_n266__, new_new_n267__,
    new_new_n268__, new_new_n269__, new_new_n271__, new_new_n272__,
    new_new_n273__, new_new_n274__, new_new_n275__, new_new_n276__,
    new_new_n277__, new_new_n278__, new_new_n279__, new_new_n280__,
    new_new_n281__, new_new_n282__, new_new_n283__, new_new_n284__,
    new_new_n285__, new_new_n286__, new_new_n287__, new_new_n288__,
    new_new_n289__, new_new_n290__, new_new_n291__, new_new_n292__,
    new_new_n293__, new_new_n294__, new_new_n295__, new_new_n296__,
    new_new_n297__, new_new_n298__, new_new_n299__, new_new_n300__,
    new_new_n301__, new_new_n302__, new_new_n303__, new_new_n304__,
    new_new_n305__, new_new_n306__, new_new_n307__, new_new_n308__,
    new_new_n309__, new_new_n310__, new_new_n311__, new_new_n312__,
    new_new_n313__, new_new_n314__, new_new_n315__, new_new_n316__,
    new_new_n317__, new_new_n318__, new_new_n319__, new_new_n320__,
    new_new_n321__, new_new_n322__, new_new_n323__, new_new_n324__,
    new_new_n325__, new_new_n326__, new_new_n327__, new_new_n328__,
    new_new_n329__, new_new_n330__, new_new_n331__, new_new_n332__,
    new_new_n333__, new_new_n334__, new_new_n335__, new_new_n336__,
    new_new_n337__, new_new_n338__, new_new_n339__, new_new_n341__,
    new_new_n342__, new_new_n343__, new_new_n344__, new_new_n345__,
    new_new_n346__, new_new_n347__, new_new_n348__, new_new_n349__,
    new_new_n350__, new_new_n351__, new_new_n352__, new_new_n353__,
    new_new_n354__, new_new_n355__, new_new_n356__, new_new_n357__,
    new_new_n358__, new_new_n359__, new_new_n360__, new_new_n361__,
    new_new_n362__, new_new_n363__, new_new_n364__, new_new_n365__,
    new_new_n366__, new_new_n367__, new_new_n368__, new_new_n369__,
    new_new_n370__, new_new_n371__, new_new_n372__, new_new_n373__,
    new_new_n374__, new_new_n375__, new_new_n376__, new_new_n377__,
    new_new_n378__, new_new_n379__, new_new_n380__, new_new_n381__,
    new_new_n382__, new_new_n383__, new_new_n384__, new_new_n385__,
    new_new_n386__, new_new_n387__, new_new_n388__, new_new_n389__,
    new_new_n390__, new_new_n391__, new_new_n392__, new_new_n393__,
    new_new_n394__, new_new_n395__, new_new_n396__, new_new_n397__,
    new_new_n398__, new_new_n399__, new_new_n400__, new_new_n401__,
    new_new_n402__, new_new_n403__, new_new_n404__, new_new_n405__,
    new_new_n406__, new_new_n407__, new_new_n408__, new_new_n409__,
    new_new_n410__, new_new_n411__, new_new_n412__, new_new_n413__,
    new_new_n414__, new_new_n416__, new_new_n417__, new_new_n418__,
    new_new_n419__, new_new_n420__, new_new_n421__, new_new_n422__,
    new_new_n423__, new_new_n424__, new_new_n425__, new_new_n426__,
    new_new_n427__, new_new_n428__, new_new_n429__, new_new_n430__,
    new_new_n431__, new_new_n432__, new_new_n433__, new_new_n434__,
    new_new_n435__, new_new_n436__, new_new_n437__, new_new_n438__,
    new_new_n439__, new_new_n440__, new_new_n441__, new_new_n442__,
    new_new_n443__, new_new_n444__, new_new_n445__, new_new_n446__,
    new_new_n447__, new_new_n448__, new_new_n449__, new_new_n450__,
    new_new_n451__, new_new_n452__, new_new_n453__, new_new_n454__,
    new_new_n455__, new_new_n456__, new_new_n457__, new_new_n458__,
    new_new_n459__, new_new_n460__, new_new_n461__, new_new_n462__,
    new_new_n463__, new_new_n464__, new_new_n465__, new_new_n466__,
    new_new_n467__, new_new_n468__, new_new_n469__, new_new_n470__,
    new_new_n471__, new_new_n472__, new_new_n473__, new_new_n474__,
    new_new_n475__, new_new_n476__, new_new_n477__, new_new_n478__,
    new_new_n479__, new_new_n480__, new_new_n481__, new_new_n482__,
    new_new_n483__, new_new_n484__, new_new_n485__, new_new_n486__,
    new_new_n487__, new_new_n488__, new_new_n489__, new_new_n490__,
    new_new_n491__, new_new_n492__, new_new_n493__, new_new_n494__,
    new_new_n495__, new_new_n496__, new_new_n497__, new_new_n499__,
    new_new_n500__, new_new_n501__, new_new_n502__, new_new_n503__,
    new_new_n504__, new_new_n505__, new_new_n506__, new_new_n507__,
    new_new_n508__, new_new_n509__, new_new_n510__, new_new_n511__,
    new_new_n512__, new_new_n513__, new_new_n514__, new_new_n515__,
    new_new_n516__, new_new_n517__, new_new_n518__, new_new_n519__,
    new_new_n520__, new_new_n521__, new_new_n522__, new_new_n523__,
    new_new_n524__, new_new_n525__, new_new_n526__, new_new_n527__,
    new_new_n528__, new_new_n529__, new_new_n530__, new_new_n531__,
    new_new_n532__, new_new_n533__, new_new_n534__, new_new_n535__,
    new_new_n536__, new_new_n537__, new_new_n538__, new_new_n539__,
    new_new_n540__, new_new_n541__, new_new_n542__, new_new_n543__,
    new_new_n544__, new_new_n545__, new_new_n546__, new_new_n547__,
    new_new_n548__, new_new_n549__, new_new_n550__, new_new_n551__,
    new_new_n552__, new_new_n553__, new_new_n554__, new_new_n555__,
    new_new_n556__, new_new_n557__, new_new_n558__, new_new_n559__,
    new_new_n560__, new_new_n561__, new_new_n562__, new_new_n563__,
    new_new_n564__, new_new_n565__, new_new_n566__, new_new_n567__,
    new_new_n568__, new_new_n569__, new_new_n570__, new_new_n571__,
    new_new_n572__, new_new_n573__, new_new_n574__, new_new_n575__,
    new_new_n576__, new_new_n577__, new_new_n578__, new_new_n579__,
    new_new_n580__, new_new_n581__, new_new_n582__, new_new_n583__,
    new_new_n584__, new_new_n585__, new_new_n586__, new_new_n587__,
    new_new_n588__, new_new_n589__, new_new_n591__, new_new_n592__,
    new_new_n593__, new_new_n594__, new_new_n595__, new_new_n596__,
    new_new_n597__, new_new_n598__, new_new_n599__, new_new_n600__,
    new_new_n601__, new_new_n602__, new_new_n603__, new_new_n604__,
    new_new_n605__, new_new_n606__, new_new_n607__, new_new_n608__,
    new_new_n609__, new_new_n610__, new_new_n611__, new_new_n612__,
    new_new_n613__, new_new_n614__, new_new_n615__, new_new_n616__,
    new_new_n617__, new_new_n618__, new_new_n619__, new_new_n620__,
    new_new_n621__, new_new_n622__, new_new_n623__, new_new_n624__,
    new_new_n625__, new_new_n626__, new_new_n627__, new_new_n628__,
    new_new_n629__, new_new_n630__, new_new_n631__, new_new_n632__,
    new_new_n633__, new_new_n634__, new_new_n635__, new_new_n636__,
    new_new_n637__, new_new_n638__, new_new_n639__, new_new_n640__,
    new_new_n641__, new_new_n642__, new_new_n643__, new_new_n644__,
    new_new_n645__, new_new_n646__, new_new_n647__, new_new_n648__,
    new_new_n649__, new_new_n650__, new_new_n651__, new_new_n652__,
    new_new_n653__, new_new_n654__, new_new_n655__, new_new_n656__,
    new_new_n657__, new_new_n658__, new_new_n659__, new_new_n660__,
    new_new_n661__, new_new_n662__, new_new_n663__, new_new_n664__,
    new_new_n665__, new_new_n666__, new_new_n667__, new_new_n668__,
    new_new_n669__, new_new_n670__, new_new_n671__, new_new_n672__,
    new_new_n673__, new_new_n674__, new_new_n675__, new_new_n676__,
    new_new_n677__, new_new_n678__, new_new_n679__, new_new_n680__,
    new_new_n681__, new_new_n682__, new_new_n683__, new_new_n684__,
    new_new_n685__, new_new_n686__, new_new_n687__, new_new_n688__,
    new_new_n689__, new_new_n690__, new_new_n691__, new_new_n693__,
    new_new_n694__, new_new_n695__, new_new_n696__, new_new_n697__,
    new_new_n698__, new_new_n699__, new_new_n700__, new_new_n701__,
    new_new_n702__, new_new_n703__, new_new_n704__, new_new_n705__,
    new_new_n706__, new_new_n707__, new_new_n708__, new_new_n709__,
    new_new_n710__, new_new_n711__, new_new_n712__, new_new_n713__,
    new_new_n714__, new_new_n715__, new_new_n716__, new_new_n717__,
    new_new_n718__, new_new_n719__, new_new_n720__, new_new_n721__,
    new_new_n722__, new_new_n723__, new_new_n724__, new_new_n725__,
    new_new_n726__, new_new_n727__, new_new_n728__, new_new_n729__,
    new_new_n730__, new_new_n731__, new_new_n732__, new_new_n733__,
    new_new_n734__, new_new_n735__, new_new_n736__, new_new_n737__,
    new_new_n738__, new_new_n739__, new_new_n740__, new_new_n741__,
    new_new_n742__, new_new_n743__, new_new_n744__, new_new_n745__,
    new_new_n746__, new_new_n747__, new_new_n748__, new_new_n749__,
    new_new_n750__, new_new_n751__, new_new_n752__, new_new_n753__,
    new_new_n754__, new_new_n755__, new_new_n756__, new_new_n757__,
    new_new_n758__, new_new_n759__, new_new_n760__, new_new_n761__,
    new_new_n762__, new_new_n763__, new_new_n764__, new_new_n765__,
    new_new_n766__, new_new_n767__, new_new_n768__, new_new_n769__,
    new_new_n770__, new_new_n771__, new_new_n772__, new_new_n773__,
    new_new_n774__, new_new_n775__, new_new_n776__, new_new_n777__,
    new_new_n778__, new_new_n779__, new_new_n780__, new_new_n781__,
    new_new_n782__, new_new_n783__, new_new_n784__, new_new_n785__,
    new_new_n786__, new_new_n787__, new_new_n788__, new_new_n789__,
    new_new_n790__, new_new_n791__, new_new_n792__, new_new_n793__,
    new_new_n794__, new_new_n795__, new_new_n797__, new_new_n798__,
    new_new_n799__, new_new_n800__, new_new_n801__, new_new_n802__,
    new_new_n803__, new_new_n804__, new_new_n805__, new_new_n806__,
    new_new_n807__, new_new_n808__, new_new_n809__, new_new_n810__,
    new_new_n811__, new_new_n812__, new_new_n813__, new_new_n814__,
    new_new_n815__, new_new_n816__, new_new_n817__, new_new_n818__,
    new_new_n819__, new_new_n820__, new_new_n821__, new_new_n822__,
    new_new_n823__, new_new_n824__, new_new_n825__, new_new_n826__,
    new_new_n827__, new_new_n828__, new_new_n829__, new_new_n830__,
    new_new_n831__, new_new_n832__, new_new_n833__, new_new_n834__,
    new_new_n835__, new_new_n836__, new_new_n837__, new_new_n838__,
    new_new_n839__, new_new_n840__, new_new_n841__, new_new_n842__,
    new_new_n843__, new_new_n844__, new_new_n845__, new_new_n846__,
    new_new_n847__, new_new_n848__, new_new_n849__, new_new_n850__,
    new_new_n851__, new_new_n852__, new_new_n853__, new_new_n854__,
    new_new_n855__, new_new_n856__, new_new_n857__, new_new_n858__,
    new_new_n859__, new_new_n860__, new_new_n861__, new_new_n862__,
    new_new_n863__, new_new_n864__, new_new_n865__, new_new_n866__,
    new_new_n867__, new_new_n868__, new_new_n869__, new_new_n870__,
    new_new_n871__, new_new_n872__, new_new_n873__, new_new_n874__,
    new_new_n875__, new_new_n876__, new_new_n877__, new_new_n878__,
    new_new_n879__, new_new_n880__, new_new_n881__, new_new_n882__,
    new_new_n883__, new_new_n884__, new_new_n885__, new_new_n886__,
    new_new_n887__, new_new_n888__, new_new_n889__, new_new_n890__,
    new_new_n891__, new_new_n892__, new_new_n893__, new_new_n894__,
    new_new_n895__, new_new_n896__, new_new_n897__, new_new_n898__,
    new_new_n899__, new_new_n900__, new_new_n901__, new_new_n902__,
    new_new_n903__, new_new_n904__, new_new_n905__, new_new_n906__,
    new_new_n907__, new_new_n908__, new_new_n909__, new_new_n910__,
    new_new_n912__, new_new_n913__, new_new_n914__, new_new_n915__,
    new_new_n916__, new_new_n917__, new_new_n918__, new_new_n919__,
    new_new_n920__, new_new_n921__, new_new_n922__, new_new_n923__,
    new_new_n924__, new_new_n925__, new_new_n926__, new_new_n927__,
    new_new_n928__, new_new_n929__, new_new_n930__, new_new_n931__,
    new_new_n932__, new_new_n933__, new_new_n934__, new_new_n935__,
    new_new_n936__, new_new_n937__, new_new_n938__, new_new_n939__,
    new_new_n940__, new_new_n941__, new_new_n942__, new_new_n943__,
    new_new_n944__, new_new_n945__, new_new_n946__, new_new_n947__,
    new_new_n948__, new_new_n949__, new_new_n950__, new_new_n951__,
    new_new_n952__, new_new_n953__, new_new_n954__, new_new_n955__,
    new_new_n956__, new_new_n957__, new_new_n958__, new_new_n959__,
    new_new_n960__, new_new_n961__, new_new_n962__, new_new_n963__,
    new_new_n964__, new_new_n965__, new_new_n966__, new_new_n967__,
    new_new_n968__, new_new_n969__, new_new_n970__, new_new_n971__,
    new_new_n972__, new_new_n973__, new_new_n974__, new_new_n975__,
    new_new_n976__, new_new_n977__, new_new_n978__, new_new_n979__,
    new_new_n980__, new_new_n981__, new_new_n982__, new_new_n983__,
    new_new_n984__, new_new_n985__, new_new_n986__, new_new_n987__,
    new_new_n988__, new_new_n989__, new_new_n990__, new_new_n991__,
    new_new_n992__, new_new_n993__, new_new_n994__, new_new_n995__,
    new_new_n996__, new_new_n997__, new_new_n998__, new_new_n999__,
    new_new_n1000__, new_new_n1001__, new_new_n1002__, new_new_n1003__,
    new_new_n1004__, new_new_n1005__, new_new_n1006__, new_new_n1007__,
    new_new_n1008__, new_new_n1009__, new_new_n1010__, new_new_n1011__,
    new_new_n1012__, new_new_n1013__, new_new_n1014__, new_new_n1015__,
    new_new_n1016__, new_new_n1017__, new_new_n1018__, new_new_n1019__,
    new_new_n1020__, new_new_n1021__, new_new_n1022__, new_new_n1023__,
    new_new_n1024__, new_new_n1025__, new_new_n1026__, new_new_n1027__,
    new_new_n1028__, new_new_n1029__, new_new_n1031__, new_new_n1032__,
    new_new_n1033__, new_new_n1034__, new_new_n1035__, new_new_n1036__,
    new_new_n1037__, new_new_n1038__, new_new_n1039__, new_new_n1040__,
    new_new_n1041__, new_new_n1042__, new_new_n1043__, new_new_n1044__,
    new_new_n1045__, new_new_n1046__, new_new_n1047__, new_new_n1048__,
    new_new_n1049__, new_new_n1050__, new_new_n1051__, new_new_n1052__,
    new_new_n1053__, new_new_n1054__, new_new_n1055__, new_new_n1056__,
    new_new_n1057__, new_new_n1058__, new_new_n1059__, new_new_n1060__,
    new_new_n1061__, new_new_n1062__, new_new_n1063__, new_new_n1064__,
    new_new_n1065__, new_new_n1066__, new_new_n1067__, new_new_n1068__,
    new_new_n1069__, new_new_n1070__, new_new_n1071__, new_new_n1072__,
    new_new_n1073__, new_new_n1074__, new_new_n1075__, new_new_n1076__,
    new_new_n1077__, new_new_n1078__, new_new_n1079__, new_new_n1080__,
    new_new_n1081__, new_new_n1082__, new_new_n1083__, new_new_n1084__,
    new_new_n1085__, new_new_n1086__, new_new_n1087__, new_new_n1088__,
    new_new_n1089__, new_new_n1090__, new_new_n1091__, new_new_n1092__,
    new_new_n1093__, new_new_n1094__, new_new_n1095__, new_new_n1096__,
    new_new_n1097__, new_new_n1098__, new_new_n1099__, new_new_n1100__,
    new_new_n1101__, new_new_n1102__, new_new_n1103__, new_new_n1104__,
    new_new_n1105__, new_new_n1106__, new_new_n1107__, new_new_n1108__,
    new_new_n1109__, new_new_n1110__, new_new_n1111__, new_new_n1112__,
    new_new_n1113__, new_new_n1114__, new_new_n1115__, new_new_n1116__,
    new_new_n1117__, new_new_n1118__, new_new_n1119__, new_new_n1120__,
    new_new_n1121__, new_new_n1122__, new_new_n1123__, new_new_n1124__,
    new_new_n1125__, new_new_n1126__, new_new_n1127__, new_new_n1128__,
    new_new_n1129__, new_new_n1130__, new_new_n1131__, new_new_n1132__,
    new_new_n1133__, new_new_n1134__, new_new_n1135__, new_new_n1136__,
    new_new_n1137__, new_new_n1138__, new_new_n1139__, new_new_n1140__,
    new_new_n1141__, new_new_n1142__, new_new_n1143__, new_new_n1144__,
    new_new_n1145__, new_new_n1146__, new_new_n1147__, new_new_n1148__,
    new_new_n1149__, new_new_n1150__, new_new_n1151__, new_new_n1152__,
    new_new_n1154__, new_new_n1155__, new_new_n1156__, new_new_n1157__,
    new_new_n1158__, new_new_n1159__, new_new_n1160__, new_new_n1161__,
    new_new_n1162__, new_new_n1163__, new_new_n1164__, new_new_n1165__,
    new_new_n1166__, new_new_n1167__, new_new_n1168__, new_new_n1169__,
    new_new_n1170__, new_new_n1171__, new_new_n1172__, new_new_n1173__,
    new_new_n1174__, new_new_n1175__, new_new_n1176__, new_new_n1177__,
    new_new_n1178__, new_new_n1179__, new_new_n1180__, new_new_n1181__,
    new_new_n1182__, new_new_n1183__, new_new_n1184__, new_new_n1185__,
    new_new_n1186__, new_new_n1187__, new_new_n1188__, new_new_n1189__,
    new_new_n1190__, new_new_n1191__, new_new_n1192__, new_new_n1193__,
    new_new_n1194__, new_new_n1195__, new_new_n1196__, new_new_n1197__,
    new_new_n1198__, new_new_n1199__, new_new_n1200__, new_new_n1201__,
    new_new_n1202__, new_new_n1203__, new_new_n1204__, new_new_n1205__,
    new_new_n1206__, new_new_n1207__, new_new_n1208__, new_new_n1209__,
    new_new_n1210__, new_new_n1211__, new_new_n1212__, new_new_n1213__,
    new_new_n1214__, new_new_n1215__, new_new_n1216__, new_new_n1217__,
    new_new_n1218__, new_new_n1219__, new_new_n1220__, new_new_n1221__,
    new_new_n1222__, new_new_n1223__, new_new_n1224__, new_new_n1225__,
    new_new_n1226__, new_new_n1227__, new_new_n1228__, new_new_n1229__,
    new_new_n1230__, new_new_n1231__, new_new_n1232__, new_new_n1233__,
    new_new_n1234__, new_new_n1235__, new_new_n1236__, new_new_n1237__,
    new_new_n1238__, new_new_n1239__, new_new_n1240__, new_new_n1241__,
    new_new_n1242__, new_new_n1243__, new_new_n1244__, new_new_n1245__,
    new_new_n1246__, new_new_n1247__, new_new_n1248__, new_new_n1249__,
    new_new_n1250__, new_new_n1251__, new_new_n1252__, new_new_n1253__,
    new_new_n1254__, new_new_n1255__, new_new_n1256__, new_new_n1257__,
    new_new_n1258__, new_new_n1259__, new_new_n1260__, new_new_n1261__,
    new_new_n1262__, new_new_n1263__, new_new_n1264__, new_new_n1266__,
    new_new_n1267__, new_new_n1268__, new_new_n1269__, new_new_n1270__,
    new_new_n1271__, new_new_n1272__, new_new_n1273__, new_new_n1274__,
    new_new_n1275__, new_new_n1276__, new_new_n1277__, new_new_n1278__,
    new_new_n1279__, new_new_n1280__, new_new_n1281__, new_new_n1282__,
    new_new_n1283__, new_new_n1284__, new_new_n1285__, new_new_n1286__,
    new_new_n1287__, new_new_n1288__, new_new_n1289__, new_new_n1290__,
    new_new_n1291__, new_new_n1292__, new_new_n1293__, new_new_n1294__,
    new_new_n1295__, new_new_n1296__, new_new_n1297__, new_new_n1298__,
    new_new_n1299__, new_new_n1300__, new_new_n1301__, new_new_n1302__,
    new_new_n1303__, new_new_n1304__, new_new_n1305__, new_new_n1306__,
    new_new_n1307__, new_new_n1308__, new_new_n1309__, new_new_n1310__,
    new_new_n1311__, new_new_n1312__, new_new_n1313__, new_new_n1314__,
    new_new_n1315__, new_new_n1316__, new_new_n1317__, new_new_n1318__,
    new_new_n1319__, new_new_n1320__, new_new_n1321__, new_new_n1322__,
    new_new_n1323__, new_new_n1324__, new_new_n1325__, new_new_n1326__,
    new_new_n1327__, new_new_n1328__, new_new_n1329__, new_new_n1330__,
    new_new_n1331__, new_new_n1332__, new_new_n1333__, new_new_n1334__,
    new_new_n1335__, new_new_n1336__, new_new_n1337__, new_new_n1338__,
    new_new_n1339__, new_new_n1340__, new_new_n1341__, new_new_n1342__,
    new_new_n1343__, new_new_n1344__, new_new_n1345__, new_new_n1346__,
    new_new_n1347__, new_new_n1348__, new_new_n1349__, new_new_n1350__,
    new_new_n1351__, new_new_n1352__, new_new_n1353__, new_new_n1354__,
    new_new_n1355__, new_new_n1356__, new_new_n1357__, new_new_n1358__,
    new_new_n1359__, new_new_n1360__, new_new_n1361__, new_new_n1362__,
    new_new_n1363__, new_new_n1364__, new_new_n1365__, new_new_n1366__,
    new_new_n1367__, new_new_n1368__, new_new_n1369__, new_new_n1370__,
    new_new_n1371__, new_new_n1372__, new_new_n1373__, new_new_n1375__,
    new_new_n1376__, new_new_n1377__, new_new_n1378__, new_new_n1379__,
    new_new_n1380__, new_new_n1381__, new_new_n1382__, new_new_n1383__,
    new_new_n1384__, new_new_n1385__, new_new_n1386__, new_new_n1387__,
    new_new_n1388__, new_new_n1389__, new_new_n1390__, new_new_n1391__,
    new_new_n1392__, new_new_n1393__, new_new_n1394__, new_new_n1395__,
    new_new_n1396__, new_new_n1397__, new_new_n1398__, new_new_n1399__,
    new_new_n1400__, new_new_n1401__, new_new_n1402__, new_new_n1403__,
    new_new_n1404__, new_new_n1405__, new_new_n1406__, new_new_n1407__,
    new_new_n1408__, new_new_n1409__, new_new_n1410__, new_new_n1411__,
    new_new_n1412__, new_new_n1413__, new_new_n1414__, new_new_n1415__,
    new_new_n1416__, new_new_n1417__, new_new_n1418__, new_new_n1419__,
    new_new_n1420__, new_new_n1421__, new_new_n1422__, new_new_n1423__,
    new_new_n1424__, new_new_n1425__, new_new_n1426__, new_new_n1427__,
    new_new_n1428__, new_new_n1429__, new_new_n1430__, new_new_n1431__,
    new_new_n1432__, new_new_n1433__, new_new_n1434__, new_new_n1435__,
    new_new_n1436__, new_new_n1437__, new_new_n1438__, new_new_n1439__,
    new_new_n1440__, new_new_n1441__, new_new_n1442__, new_new_n1443__,
    new_new_n1444__, new_new_n1445__, new_new_n1446__, new_new_n1447__,
    new_new_n1448__, new_new_n1449__, new_new_n1450__, new_new_n1451__,
    new_new_n1452__, new_new_n1453__, new_new_n1454__, new_new_n1455__,
    new_new_n1456__, new_new_n1457__, new_new_n1458__, new_new_n1459__,
    new_new_n1460__, new_new_n1461__, new_new_n1462__, new_new_n1463__,
    new_new_n1464__, new_new_n1465__, new_new_n1466__, new_new_n1467__,
    new_new_n1468__, new_new_n1469__, new_new_n1470__, new_new_n1471__,
    new_new_n1472__, new_new_n1474__, new_new_n1475__, new_new_n1476__,
    new_new_n1477__, new_new_n1478__, new_new_n1479__, new_new_n1480__,
    new_new_n1481__, new_new_n1482__, new_new_n1483__, new_new_n1484__,
    new_new_n1485__, new_new_n1486__, new_new_n1487__, new_new_n1488__,
    new_new_n1489__, new_new_n1490__, new_new_n1491__, new_new_n1492__,
    new_new_n1493__, new_new_n1494__, new_new_n1495__, new_new_n1496__,
    new_new_n1497__, new_new_n1498__, new_new_n1499__, new_new_n1500__,
    new_new_n1501__, new_new_n1502__, new_new_n1503__, new_new_n1504__,
    new_new_n1505__, new_new_n1506__, new_new_n1507__, new_new_n1508__,
    new_new_n1509__, new_new_n1510__, new_new_n1511__, new_new_n1512__,
    new_new_n1513__, new_new_n1514__, new_new_n1515__, new_new_n1516__,
    new_new_n1517__, new_new_n1518__, new_new_n1519__, new_new_n1520__,
    new_new_n1521__, new_new_n1522__, new_new_n1523__, new_new_n1524__,
    new_new_n1525__, new_new_n1526__, new_new_n1527__, new_new_n1528__,
    new_new_n1529__, new_new_n1530__, new_new_n1531__, new_new_n1532__,
    new_new_n1533__, new_new_n1534__, new_new_n1535__, new_new_n1536__,
    new_new_n1537__, new_new_n1538__, new_new_n1539__, new_new_n1540__,
    new_new_n1541__, new_new_n1542__, new_new_n1543__, new_new_n1544__,
    new_new_n1545__, new_new_n1546__, new_new_n1547__, new_new_n1548__,
    new_new_n1549__, new_new_n1550__, new_new_n1551__, new_new_n1552__,
    new_new_n1553__, new_new_n1554__, new_new_n1555__, new_new_n1556__,
    new_new_n1557__, new_new_n1558__, new_new_n1559__, new_new_n1560__,
    new_new_n1561__, new_new_n1562__, new_new_n1563__, new_new_n1564__,
    new_new_n1565__, new_new_n1566__, new_new_n1567__, new_new_n1568__,
    new_new_n1569__, new_new_n1570__, new_new_n1571__, new_new_n1573__,
    new_new_n1574__, new_new_n1575__, new_new_n1576__, new_new_n1577__,
    new_new_n1578__, new_new_n1579__, new_new_n1580__, new_new_n1581__,
    new_new_n1582__, new_new_n1583__, new_new_n1584__, new_new_n1585__,
    new_new_n1586__, new_new_n1587__, new_new_n1588__, new_new_n1589__,
    new_new_n1590__, new_new_n1591__, new_new_n1592__, new_new_n1593__,
    new_new_n1594__, new_new_n1595__, new_new_n1596__, new_new_n1597__,
    new_new_n1598__, new_new_n1599__, new_new_n1600__, new_new_n1601__,
    new_new_n1602__, new_new_n1603__, new_new_n1604__, new_new_n1605__,
    new_new_n1606__, new_new_n1607__, new_new_n1608__, new_new_n1609__,
    new_new_n1610__, new_new_n1611__, new_new_n1612__, new_new_n1613__,
    new_new_n1614__, new_new_n1615__, new_new_n1616__, new_new_n1617__,
    new_new_n1618__, new_new_n1619__, new_new_n1620__, new_new_n1621__,
    new_new_n1622__, new_new_n1623__, new_new_n1624__, new_new_n1625__,
    new_new_n1626__, new_new_n1627__, new_new_n1628__, new_new_n1629__,
    new_new_n1630__, new_new_n1631__, new_new_n1632__, new_new_n1633__,
    new_new_n1634__, new_new_n1635__, new_new_n1636__, new_new_n1637__,
    new_new_n1638__, new_new_n1639__, new_new_n1640__, new_new_n1641__,
    new_new_n1642__, new_new_n1643__, new_new_n1644__, new_new_n1645__,
    new_new_n1646__, new_new_n1647__, new_new_n1648__, new_new_n1649__,
    new_new_n1650__, new_new_n1651__, new_new_n1652__, new_new_n1653__,
    new_new_n1654__, new_new_n1655__, new_new_n1657__, new_new_n1658__,
    new_new_n1659__, new_new_n1660__, new_new_n1661__, new_new_n1662__,
    new_new_n1663__, new_new_n1664__, new_new_n1665__, new_new_n1666__,
    new_new_n1667__, new_new_n1668__, new_new_n1669__, new_new_n1670__,
    new_new_n1671__, new_new_n1672__, new_new_n1673__, new_new_n1674__,
    new_new_n1675__, new_new_n1676__, new_new_n1677__, new_new_n1678__,
    new_new_n1679__, new_new_n1680__, new_new_n1681__, new_new_n1682__,
    new_new_n1683__, new_new_n1684__, new_new_n1685__, new_new_n1686__,
    new_new_n1687__, new_new_n1688__, new_new_n1689__, new_new_n1690__,
    new_new_n1691__, new_new_n1692__, new_new_n1693__, new_new_n1694__,
    new_new_n1695__, new_new_n1696__, new_new_n1697__, new_new_n1698__,
    new_new_n1699__, new_new_n1700__, new_new_n1701__, new_new_n1702__,
    new_new_n1703__, new_new_n1704__, new_new_n1705__, new_new_n1706__,
    new_new_n1707__, new_new_n1708__, new_new_n1709__, new_new_n1710__,
    new_new_n1711__, new_new_n1712__, new_new_n1713__, new_new_n1714__,
    new_new_n1715__, new_new_n1716__, new_new_n1717__, new_new_n1718__,
    new_new_n1719__, new_new_n1720__, new_new_n1721__, new_new_n1722__,
    new_new_n1723__, new_new_n1724__, new_new_n1725__, new_new_n1726__,
    new_new_n1727__, new_new_n1728__, new_new_n1729__, new_new_n1730__,
    new_new_n1731__, new_new_n1732__, new_new_n1734__, new_new_n1735__,
    new_new_n1736__, new_new_n1737__, new_new_n1738__, new_new_n1739__,
    new_new_n1740__, new_new_n1741__, new_new_n1742__, new_new_n1743__,
    new_new_n1744__, new_new_n1745__, new_new_n1746__, new_new_n1747__,
    new_new_n1748__, new_new_n1749__, new_new_n1750__, new_new_n1751__,
    new_new_n1752__, new_new_n1753__, new_new_n1754__, new_new_n1755__,
    new_new_n1756__, new_new_n1757__, new_new_n1758__, new_new_n1759__,
    new_new_n1760__, new_new_n1761__, new_new_n1762__, new_new_n1763__,
    new_new_n1764__, new_new_n1765__, new_new_n1766__, new_new_n1767__,
    new_new_n1768__, new_new_n1769__, new_new_n1770__, new_new_n1771__,
    new_new_n1772__, new_new_n1773__, new_new_n1774__, new_new_n1775__,
    new_new_n1776__, new_new_n1777__, new_new_n1778__, new_new_n1779__,
    new_new_n1780__, new_new_n1781__, new_new_n1782__, new_new_n1783__,
    new_new_n1784__, new_new_n1785__, new_new_n1786__, new_new_n1787__,
    new_new_n1788__, new_new_n1789__, new_new_n1790__, new_new_n1791__,
    new_new_n1792__, new_new_n1793__, new_new_n1794__, new_new_n1795__,
    new_new_n1796__, new_new_n1797__, new_new_n1798__, new_new_n1799__,
    new_new_n1800__, new_new_n1802__, new_new_n1803__, new_new_n1804__,
    new_new_n1805__, new_new_n1806__, new_new_n1807__, new_new_n1808__,
    new_new_n1809__, new_new_n1810__, new_new_n1811__, new_new_n1812__,
    new_new_n1813__, new_new_n1814__, new_new_n1815__, new_new_n1816__,
    new_new_n1817__, new_new_n1818__, new_new_n1819__, new_new_n1820__,
    new_new_n1821__, new_new_n1822__, new_new_n1823__, new_new_n1824__,
    new_new_n1825__, new_new_n1826__, new_new_n1827__, new_new_n1828__,
    new_new_n1829__, new_new_n1830__, new_new_n1831__, new_new_n1832__,
    new_new_n1833__, new_new_n1834__, new_new_n1835__, new_new_n1836__,
    new_new_n1837__, new_new_n1838__, new_new_n1839__, new_new_n1840__,
    new_new_n1841__, new_new_n1842__, new_new_n1843__, new_new_n1844__,
    new_new_n1845__, new_new_n1846__, new_new_n1847__, new_new_n1848__,
    new_new_n1849__, new_new_n1850__, new_new_n1851__, new_new_n1852__,
    new_new_n1853__, new_new_n1854__, new_new_n1855__, new_new_n1856__,
    new_new_n1857__, new_new_n1858__, new_new_n1859__, new_new_n1860__,
    new_new_n1861__, new_new_n1862__, new_new_n1863__, new_new_n1864__,
    new_new_n1865__, new_new_n1866__, new_new_n1867__, new_new_n1868__,
    new_new_n1869__, new_new_n1870__, new_new_n1871__, new_new_n1872__,
    new_new_n1873__, new_new_n1874__, new_new_n1875__, new_new_n1877__,
    new_new_n1878__, new_new_n1879__, new_new_n1880__, new_new_n1881__,
    new_new_n1882__, new_new_n1883__, new_new_n1884__, new_new_n1885__,
    new_new_n1886__, new_new_n1887__, new_new_n1888__, new_new_n1889__,
    new_new_n1890__, new_new_n1891__, new_new_n1892__, new_new_n1893__,
    new_new_n1894__, new_new_n1895__, new_new_n1896__, new_new_n1897__,
    new_new_n1898__, new_new_n1899__, new_new_n1900__, new_new_n1901__,
    new_new_n1902__, new_new_n1903__, new_new_n1904__, new_new_n1905__,
    new_new_n1906__, new_new_n1907__, new_new_n1908__, new_new_n1909__,
    new_new_n1910__, new_new_n1911__, new_new_n1912__, new_new_n1913__,
    new_new_n1914__, new_new_n1915__, new_new_n1916__, new_new_n1917__,
    new_new_n1918__, new_new_n1919__, new_new_n1920__, new_new_n1921__,
    new_new_n1922__, new_new_n1923__, new_new_n1924__, new_new_n1925__,
    new_new_n1926__, new_new_n1927__, new_new_n1928__, new_new_n1930__,
    new_new_n1931__, new_new_n1932__, new_new_n1933__, new_new_n1934__,
    new_new_n1935__, new_new_n1936__, new_new_n1937__, new_new_n1938__,
    new_new_n1939__, new_new_n1940__, new_new_n1941__, new_new_n1942__,
    new_new_n1943__, new_new_n1944__, new_new_n1945__, new_new_n1946__,
    new_new_n1947__, new_new_n1948__, new_new_n1949__, new_new_n1950__,
    new_new_n1951__, new_new_n1952__, new_new_n1953__, new_new_n1954__,
    new_new_n1955__, new_new_n1956__, new_new_n1957__, new_new_n1958__,
    new_new_n1959__, new_new_n1960__, new_new_n1961__, new_new_n1962__,
    new_new_n1963__, new_new_n1964__, new_new_n1965__, new_new_n1966__,
    new_new_n1967__, new_new_n1968__, new_new_n1969__, new_new_n1970__,
    new_new_n1971__, new_new_n1972__, new_new_n1973__, new_new_n1974__,
    new_new_n1976__, new_new_n1977__, new_new_n1978__, new_new_n1979__,
    new_new_n1980__, new_new_n1981__, new_new_n1982__, new_new_n1983__,
    new_new_n1984__, new_new_n1985__, new_new_n1986__, new_new_n1987__,
    new_new_n1988__, new_new_n1989__, new_new_n1990__, new_new_n1991__,
    new_new_n1992__, new_new_n1993__, new_new_n1994__, new_new_n1995__,
    new_new_n1996__, new_new_n1997__, new_new_n1998__, new_new_n1999__,
    new_new_n2000__, new_new_n2001__, new_new_n2002__, new_new_n2003__,
    new_new_n2004__, new_new_n2005__, new_new_n2006__, new_new_n2007__,
    new_new_n2008__, new_new_n2009__, new_new_n2010__, new_new_n2011__,
    new_new_n2012__, new_new_n2013__, new_new_n2015__, new_new_n2016__,
    new_new_n2017__, new_new_n2018__, new_new_n2019__, new_new_n2020__,
    new_new_n2021__, new_new_n2022__, new_new_n2023__, new_new_n2024__,
    new_new_n2025__, new_new_n2026__, new_new_n2027__, new_new_n2028__,
    new_new_n2029__, new_new_n2030__, new_new_n2031__, new_new_n2032__,
    new_new_n2033__, new_new_n2034__, new_new_n2035__, new_new_n2036__,
    new_new_n2037__, new_new_n2038__, new_new_n2039__, new_new_n2040__,
    new_new_n2041__, new_new_n2042__, new_new_n2043__, new_new_n2044__,
    new_new_n2045__, new_new_n2046__, new_new_n2047__, new_new_n2048__,
    new_new_n2049__, new_new_n2050__, new_new_n2051__, new_new_n2052__,
    new_new_n2053__, new_new_n2055__, new_new_n2056__, new_new_n2057__,
    new_new_n2058__, new_new_n2059__, new_new_n2060__, new_new_n2061__,
    new_new_n2062__, new_new_n2063__, new_new_n2064__, new_new_n2065__,
    new_new_n2066__, new_new_n2067__, new_new_n2068__, new_new_n2069__,
    new_new_n2070__, new_new_n2071__, new_new_n2072__, new_new_n2073__,
    new_new_n2074__, new_new_n2075__, new_new_n2076__, new_new_n2077__,
    new_new_n2079__, new_new_n2080__, new_new_n2081__, new_new_n2082__,
    new_new_n2083__, new_new_n2084__, new_new_n2085__, new_new_n2086__,
    new_new_n2087__, new_new_n2088__, new_new_n2089__, new_new_n2090__,
    new_new_n2091__, new_new_n2092__, new_new_n2094__, new_new_n2095__,
    new_new_n2096__;
  assign \r[0]  = \a[0]  & \b[0] ;
  assign new_new_n66__ = \a[1]  & \b[0] ;
  assign new_new_n67__ = \a[0]  & \b[1] ;
  assign new_new_n68__ = ~new_new_n66__ & ~new_new_n67__;
  assign new_new_n69__ = new_new_n66__ & new_new_n67__;
  assign \r[1]  = ~new_new_n68__ & ~new_new_n69__;
  assign new_new_n71__ = \a[0]  & \b[2] ;
  assign new_new_n72__ = \a[1]  & \b[1] ;
  assign new_new_n73__ = \a[2]  & \b[0] ;
  assign new_new_n74__ = ~new_new_n72__ & ~new_new_n73__;
  assign new_new_n75__ = new_new_n72__ & new_new_n73__;
  assign new_new_n76__ = ~new_new_n69__ & new_new_n75__;
  assign new_new_n77__ = new_new_n69__ & ~new_new_n75__;
  assign new_new_n78__ = ~new_new_n74__ & ~new_new_n76__;
  assign new_new_n79__ = ~new_new_n77__ & new_new_n78__;
  assign new_new_n80__ = new_new_n71__ & new_new_n79__;
  assign new_new_n81__ = ~new_new_n71__ & ~new_new_n79__;
  assign \r[2]  = ~new_new_n80__ & ~new_new_n81__;
  assign new_new_n83__ = ~new_new_n77__ & ~new_new_n80__;
  assign new_new_n84__ = \a[1]  & \b[2] ;
  assign new_new_n85__ = \a[3]  & \b[0] ;
  assign new_new_n86__ = \a[0]  & \b[3] ;
  assign new_new_n87__ = ~new_new_n85__ & ~new_new_n86__;
  assign new_new_n88__ = new_new_n85__ & new_new_n86__;
  assign new_new_n89__ = ~new_new_n87__ & ~new_new_n88__;
  assign new_new_n90__ = \a[2]  & \b[1] ;
  assign new_new_n91__ = ~new_new_n66__ & new_new_n90__;
  assign new_new_n92__ = new_new_n89__ & ~new_new_n91__;
  assign new_new_n93__ = ~new_new_n89__ & new_new_n91__;
  assign new_new_n94__ = ~new_new_n92__ & ~new_new_n93__;
  assign new_new_n95__ = new_new_n84__ & ~new_new_n94__;
  assign new_new_n96__ = ~new_new_n84__ & new_new_n94__;
  assign new_new_n97__ = ~new_new_n95__ & ~new_new_n96__;
  assign new_new_n98__ = ~new_new_n83__ & new_new_n97__;
  assign new_new_n99__ = new_new_n83__ & ~new_new_n97__;
  assign \r[3]  = ~new_new_n98__ & ~new_new_n99__;
  assign new_new_n101__ = new_new_n75__ & ~new_new_n89__;
  assign new_new_n102__ = ~new_new_n95__ & ~new_new_n101__;
  assign new_new_n103__ = \a[0]  & \b[4] ;
  assign new_new_n104__ = \a[2]  & \b[2] ;
  assign new_new_n105__ = ~new_new_n103__ & ~new_new_n104__;
  assign new_new_n106__ = new_new_n103__ & new_new_n104__;
  assign new_new_n107__ = ~new_new_n105__ & ~new_new_n106__;
  assign new_new_n108__ = \a[3]  & \b[1] ;
  assign new_new_n109__ = \a[4]  & \b[0] ;
  assign new_new_n110__ = \a[1]  & \b[3] ;
  assign new_new_n111__ = ~new_new_n109__ & ~new_new_n110__;
  assign new_new_n112__ = new_new_n109__ & new_new_n110__;
  assign new_new_n113__ = ~new_new_n111__ & ~new_new_n112__;
  assign new_new_n114__ = new_new_n108__ & new_new_n113__;
  assign new_new_n115__ = ~new_new_n108__ & ~new_new_n113__;
  assign new_new_n116__ = ~new_new_n114__ & ~new_new_n115__;
  assign new_new_n117__ = ~new_new_n88__ & ~new_new_n90__;
  assign new_new_n118__ = ~new_new_n87__ & ~new_new_n117__;
  assign new_new_n119__ = new_new_n116__ & new_new_n118__;
  assign new_new_n120__ = ~new_new_n116__ & ~new_new_n118__;
  assign new_new_n121__ = ~new_new_n119__ & ~new_new_n120__;
  assign new_new_n122__ = ~new_new_n107__ & ~new_new_n121__;
  assign new_new_n123__ = new_new_n107__ & new_new_n121__;
  assign new_new_n124__ = ~new_new_n122__ & ~new_new_n123__;
  assign new_new_n125__ = new_new_n102__ & ~new_new_n124__;
  assign new_new_n126__ = ~new_new_n102__ & new_new_n124__;
  assign new_new_n127__ = ~new_new_n125__ & ~new_new_n126__;
  assign new_new_n128__ = new_new_n98__ & new_new_n127__;
  assign new_new_n129__ = ~new_new_n98__ & ~new_new_n127__;
  assign \r[4]  = ~new_new_n128__ & ~new_new_n129__;
  assign new_new_n131__ = ~new_new_n119__ & ~new_new_n123__;
  assign new_new_n132__ = \a[0]  & \b[5] ;
  assign new_new_n133__ = \a[1]  & \b[4] ;
  assign new_new_n134__ = \a[3]  & \b[2] ;
  assign new_new_n135__ = ~new_new_n133__ & ~new_new_n134__;
  assign new_new_n136__ = new_new_n133__ & new_new_n134__;
  assign new_new_n137__ = ~new_new_n135__ & ~new_new_n136__;
  assign new_new_n138__ = new_new_n132__ & new_new_n137__;
  assign new_new_n139__ = ~new_new_n132__ & ~new_new_n137__;
  assign new_new_n140__ = ~new_new_n138__ & ~new_new_n139__;
  assign new_new_n141__ = ~new_new_n112__ & ~new_new_n114__;
  assign new_new_n142__ = \a[4]  & \b[1] ;
  assign new_new_n143__ = \a[5]  & \b[0] ;
  assign new_new_n144__ = \a[2]  & \b[3] ;
  assign new_new_n145__ = ~new_new_n143__ & ~new_new_n144__;
  assign new_new_n146__ = new_new_n143__ & new_new_n144__;
  assign new_new_n147__ = ~new_new_n145__ & ~new_new_n146__;
  assign new_new_n148__ = new_new_n142__ & new_new_n147__;
  assign new_new_n149__ = ~new_new_n142__ & ~new_new_n147__;
  assign new_new_n150__ = ~new_new_n148__ & ~new_new_n149__;
  assign new_new_n151__ = ~new_new_n141__ & new_new_n150__;
  assign new_new_n152__ = new_new_n141__ & ~new_new_n150__;
  assign new_new_n153__ = ~new_new_n151__ & ~new_new_n152__;
  assign new_new_n154__ = new_new_n140__ & new_new_n153__;
  assign new_new_n155__ = ~new_new_n140__ & ~new_new_n153__;
  assign new_new_n156__ = ~new_new_n154__ & ~new_new_n155__;
  assign new_new_n157__ = ~new_new_n131__ & new_new_n156__;
  assign new_new_n158__ = new_new_n131__ & ~new_new_n156__;
  assign new_new_n159__ = ~new_new_n157__ & ~new_new_n158__;
  assign new_new_n160__ = new_new_n106__ & new_new_n159__;
  assign new_new_n161__ = ~new_new_n106__ & ~new_new_n159__;
  assign new_new_n162__ = ~new_new_n160__ & ~new_new_n161__;
  assign new_new_n163__ = ~new_new_n126__ & ~new_new_n128__;
  assign new_new_n164__ = new_new_n162__ & new_new_n163__;
  assign new_new_n165__ = ~new_new_n162__ & ~new_new_n163__;
  assign \r[5]  = new_new_n164__ | new_new_n165__;
  assign new_new_n167__ = new_new_n126__ & new_new_n162__;
  assign new_new_n168__ = ~new_new_n157__ & ~new_new_n160__;
  assign new_new_n169__ = \a[0]  & \b[6] ;
  assign new_new_n170__ = ~new_new_n136__ & ~new_new_n138__;
  assign new_new_n171__ = new_new_n169__ & ~new_new_n170__;
  assign new_new_n172__ = ~new_new_n169__ & new_new_n170__;
  assign new_new_n173__ = ~new_new_n171__ & ~new_new_n172__;
  assign new_new_n174__ = ~new_new_n151__ & ~new_new_n154__;
  assign new_new_n175__ = \a[1]  & \b[5] ;
  assign new_new_n176__ = \a[2]  & \b[4] ;
  assign new_new_n177__ = \a[4]  & \b[2] ;
  assign new_new_n178__ = ~new_new_n176__ & ~new_new_n177__;
  assign new_new_n179__ = new_new_n176__ & new_new_n177__;
  assign new_new_n180__ = ~new_new_n178__ & ~new_new_n179__;
  assign new_new_n181__ = new_new_n175__ & new_new_n180__;
  assign new_new_n182__ = ~new_new_n175__ & ~new_new_n180__;
  assign new_new_n183__ = ~new_new_n181__ & ~new_new_n182__;
  assign new_new_n184__ = ~new_new_n146__ & ~new_new_n148__;
  assign new_new_n185__ = \a[5]  & \b[1] ;
  assign new_new_n186__ = \a[3]  & \b[3] ;
  assign new_new_n187__ = \a[6]  & \b[0] ;
  assign new_new_n188__ = ~new_new_n186__ & ~new_new_n187__;
  assign new_new_n189__ = new_new_n186__ & new_new_n187__;
  assign new_new_n190__ = ~new_new_n188__ & ~new_new_n189__;
  assign new_new_n191__ = new_new_n185__ & new_new_n190__;
  assign new_new_n192__ = ~new_new_n185__ & ~new_new_n190__;
  assign new_new_n193__ = ~new_new_n191__ & ~new_new_n192__;
  assign new_new_n194__ = ~new_new_n184__ & new_new_n193__;
  assign new_new_n195__ = new_new_n184__ & ~new_new_n193__;
  assign new_new_n196__ = ~new_new_n194__ & ~new_new_n195__;
  assign new_new_n197__ = new_new_n183__ & new_new_n196__;
  assign new_new_n198__ = ~new_new_n183__ & ~new_new_n196__;
  assign new_new_n199__ = ~new_new_n197__ & ~new_new_n198__;
  assign new_new_n200__ = ~new_new_n174__ & new_new_n199__;
  assign new_new_n201__ = new_new_n174__ & ~new_new_n199__;
  assign new_new_n202__ = ~new_new_n200__ & ~new_new_n201__;
  assign new_new_n203__ = new_new_n173__ & new_new_n202__;
  assign new_new_n204__ = ~new_new_n173__ & ~new_new_n202__;
  assign new_new_n205__ = ~new_new_n203__ & ~new_new_n204__;
  assign new_new_n206__ = new_new_n168__ & ~new_new_n205__;
  assign new_new_n207__ = ~new_new_n168__ & new_new_n205__;
  assign new_new_n208__ = ~new_new_n206__ & ~new_new_n207__;
  assign new_new_n209__ = ~new_new_n167__ & ~new_new_n208__;
  assign new_new_n210__ = new_new_n167__ & new_new_n208__;
  assign new_new_n211__ = ~new_new_n209__ & ~new_new_n210__;
  assign new_new_n212__ = new_new_n128__ & new_new_n162__;
  assign new_new_n213__ = new_new_n211__ & new_new_n212__;
  assign new_new_n214__ = ~new_new_n211__ & ~new_new_n212__;
  assign \r[6]  = ~new_new_n213__ & ~new_new_n214__;
  assign new_new_n216__ = ~new_new_n200__ & ~new_new_n203__;
  assign new_new_n217__ = ~new_new_n194__ & ~new_new_n197__;
  assign new_new_n218__ = ~new_new_n189__ & ~new_new_n191__;
  assign new_new_n219__ = \a[4]  & \b[3] ;
  assign new_new_n220__ = \a[7]  & \b[0] ;
  assign new_new_n221__ = ~new_new_n219__ & ~new_new_n220__;
  assign new_new_n222__ = new_new_n219__ & new_new_n220__;
  assign new_new_n223__ = ~new_new_n221__ & ~new_new_n222__;
  assign new_new_n224__ = \a[6]  & \b[1] ;
  assign new_new_n225__ = new_new_n223__ & new_new_n224__;
  assign new_new_n226__ = ~new_new_n223__ & ~new_new_n224__;
  assign new_new_n227__ = ~new_new_n225__ & ~new_new_n226__;
  assign new_new_n228__ = new_new_n218__ & ~new_new_n227__;
  assign new_new_n229__ = ~new_new_n218__ & new_new_n227__;
  assign new_new_n230__ = ~new_new_n228__ & ~new_new_n229__;
  assign new_new_n231__ = \a[2]  & \b[5] ;
  assign new_new_n232__ = \a[3]  & \b[4] ;
  assign new_new_n233__ = \a[5]  & \b[2] ;
  assign new_new_n234__ = ~new_new_n232__ & ~new_new_n233__;
  assign new_new_n235__ = new_new_n232__ & new_new_n233__;
  assign new_new_n236__ = ~new_new_n234__ & ~new_new_n235__;
  assign new_new_n237__ = ~new_new_n231__ & ~new_new_n236__;
  assign new_new_n238__ = new_new_n231__ & new_new_n236__;
  assign new_new_n239__ = ~new_new_n237__ & ~new_new_n238__;
  assign new_new_n240__ = new_new_n230__ & new_new_n239__;
  assign new_new_n241__ = ~new_new_n230__ & ~new_new_n239__;
  assign new_new_n242__ = ~new_new_n240__ & ~new_new_n241__;
  assign new_new_n243__ = new_new_n217__ & ~new_new_n242__;
  assign new_new_n244__ = ~new_new_n217__ & new_new_n242__;
  assign new_new_n245__ = ~new_new_n243__ & ~new_new_n244__;
  assign new_new_n246__ = \a[0]  & \b[7] ;
  assign new_new_n247__ = \a[1]  & \b[6] ;
  assign new_new_n248__ = ~new_new_n246__ & ~new_new_n247__;
  assign new_new_n249__ = new_new_n246__ & new_new_n247__;
  assign new_new_n250__ = ~new_new_n248__ & ~new_new_n249__;
  assign new_new_n251__ = ~new_new_n179__ & ~new_new_n181__;
  assign new_new_n252__ = ~new_new_n250__ & new_new_n251__;
  assign new_new_n253__ = new_new_n250__ & ~new_new_n251__;
  assign new_new_n254__ = ~new_new_n252__ & ~new_new_n253__;
  assign new_new_n255__ = new_new_n245__ & new_new_n254__;
  assign new_new_n256__ = ~new_new_n245__ & ~new_new_n254__;
  assign new_new_n257__ = ~new_new_n255__ & ~new_new_n256__;
  assign new_new_n258__ = new_new_n216__ & ~new_new_n257__;
  assign new_new_n259__ = ~new_new_n216__ & new_new_n257__;
  assign new_new_n260__ = ~new_new_n258__ & ~new_new_n259__;
  assign new_new_n261__ = new_new_n171__ & new_new_n260__;
  assign new_new_n262__ = ~new_new_n171__ & ~new_new_n260__;
  assign new_new_n263__ = ~new_new_n261__ & ~new_new_n262__;
  assign new_new_n264__ = ~new_new_n207__ & ~new_new_n210__;
  assign new_new_n265__ = new_new_n263__ & new_new_n264__;
  assign new_new_n266__ = ~new_new_n263__ & ~new_new_n264__;
  assign new_new_n267__ = ~new_new_n265__ & ~new_new_n266__;
  assign new_new_n268__ = new_new_n213__ & ~new_new_n267__;
  assign new_new_n269__ = ~new_new_n213__ & new_new_n267__;
  assign \r[7]  = ~new_new_n268__ & ~new_new_n269__;
  assign new_new_n271__ = new_new_n207__ & new_new_n263__;
  assign new_new_n272__ = ~new_new_n259__ & ~new_new_n261__;
  assign new_new_n273__ = ~new_new_n244__ & ~new_new_n255__;
  assign new_new_n274__ = \a[0]  & \b[8] ;
  assign new_new_n275__ = \a[1]  & \b[7] ;
  assign new_new_n276__ = \a[2]  & \b[6] ;
  assign new_new_n277__ = ~new_new_n275__ & ~new_new_n276__;
  assign new_new_n278__ = new_new_n275__ & new_new_n276__;
  assign new_new_n279__ = ~new_new_n277__ & ~new_new_n278__;
  assign new_new_n280__ = new_new_n274__ & new_new_n279__;
  assign new_new_n281__ = ~new_new_n274__ & ~new_new_n279__;
  assign new_new_n282__ = ~new_new_n280__ & ~new_new_n281__;
  assign new_new_n283__ = ~new_new_n235__ & ~new_new_n238__;
  assign new_new_n284__ = new_new_n282__ & ~new_new_n283__;
  assign new_new_n285__ = ~new_new_n282__ & new_new_n283__;
  assign new_new_n286__ = ~new_new_n284__ & ~new_new_n285__;
  assign new_new_n287__ = new_new_n249__ & new_new_n286__;
  assign new_new_n288__ = ~new_new_n249__ & ~new_new_n286__;
  assign new_new_n289__ = ~new_new_n287__ & ~new_new_n288__;
  assign new_new_n290__ = ~new_new_n229__ & ~new_new_n240__;
  assign new_new_n291__ = \a[3]  & \b[5] ;
  assign new_new_n292__ = \a[4]  & \b[4] ;
  assign new_new_n293__ = \a[6]  & \b[2] ;
  assign new_new_n294__ = ~new_new_n292__ & ~new_new_n293__;
  assign new_new_n295__ = new_new_n292__ & new_new_n293__;
  assign new_new_n296__ = ~new_new_n294__ & ~new_new_n295__;
  assign new_new_n297__ = new_new_n291__ & new_new_n296__;
  assign new_new_n298__ = ~new_new_n291__ & ~new_new_n296__;
  assign new_new_n299__ = ~new_new_n297__ & ~new_new_n298__;
  assign new_new_n300__ = ~new_new_n222__ & ~new_new_n225__;
  assign new_new_n301__ = \a[7]  & \b[1] ;
  assign new_new_n302__ = \a[5]  & \b[3] ;
  assign new_new_n303__ = \a[8]  & \b[0] ;
  assign new_new_n304__ = ~new_new_n302__ & ~new_new_n303__;
  assign new_new_n305__ = new_new_n302__ & new_new_n303__;
  assign new_new_n306__ = ~new_new_n304__ & ~new_new_n305__;
  assign new_new_n307__ = new_new_n301__ & new_new_n306__;
  assign new_new_n308__ = ~new_new_n301__ & ~new_new_n306__;
  assign new_new_n309__ = ~new_new_n307__ & ~new_new_n308__;
  assign new_new_n310__ = ~new_new_n300__ & new_new_n309__;
  assign new_new_n311__ = new_new_n300__ & ~new_new_n309__;
  assign new_new_n312__ = ~new_new_n310__ & ~new_new_n311__;
  assign new_new_n313__ = new_new_n299__ & new_new_n312__;
  assign new_new_n314__ = ~new_new_n299__ & ~new_new_n312__;
  assign new_new_n315__ = ~new_new_n313__ & ~new_new_n314__;
  assign new_new_n316__ = ~new_new_n290__ & new_new_n315__;
  assign new_new_n317__ = new_new_n290__ & ~new_new_n315__;
  assign new_new_n318__ = ~new_new_n316__ & ~new_new_n317__;
  assign new_new_n319__ = new_new_n289__ & new_new_n318__;
  assign new_new_n320__ = ~new_new_n289__ & ~new_new_n318__;
  assign new_new_n321__ = ~new_new_n319__ & ~new_new_n320__;
  assign new_new_n322__ = ~new_new_n273__ & new_new_n321__;
  assign new_new_n323__ = new_new_n273__ & ~new_new_n321__;
  assign new_new_n324__ = ~new_new_n322__ & ~new_new_n323__;
  assign new_new_n325__ = new_new_n253__ & new_new_n324__;
  assign new_new_n326__ = ~new_new_n253__ & ~new_new_n324__;
  assign new_new_n327__ = ~new_new_n325__ & ~new_new_n326__;
  assign new_new_n328__ = new_new_n272__ & ~new_new_n327__;
  assign new_new_n329__ = ~new_new_n272__ & new_new_n327__;
  assign new_new_n330__ = ~new_new_n328__ & ~new_new_n329__;
  assign new_new_n331__ = new_new_n271__ & new_new_n330__;
  assign new_new_n332__ = ~new_new_n271__ & ~new_new_n330__;
  assign new_new_n333__ = ~new_new_n331__ & ~new_new_n332__;
  assign new_new_n334__ = new_new_n210__ & new_new_n263__;
  assign new_new_n335__ = new_new_n333__ & new_new_n334__;
  assign new_new_n336__ = ~new_new_n333__ & ~new_new_n334__;
  assign new_new_n337__ = ~new_new_n335__ & ~new_new_n336__;
  assign new_new_n338__ = new_new_n268__ & new_new_n337__;
  assign new_new_n339__ = ~new_new_n268__ & ~new_new_n337__;
  assign \r[8]  = ~new_new_n338__ & ~new_new_n339__;
  assign new_new_n341__ = ~new_new_n322__ & ~new_new_n325__;
  assign new_new_n342__ = \a[0]  & \b[9] ;
  assign new_new_n343__ = ~new_new_n284__ & ~new_new_n287__;
  assign new_new_n344__ = new_new_n342__ & ~new_new_n343__;
  assign new_new_n345__ = ~new_new_n342__ & new_new_n343__;
  assign new_new_n346__ = ~new_new_n344__ & ~new_new_n345__;
  assign new_new_n347__ = ~new_new_n316__ & ~new_new_n319__;
  assign new_new_n348__ = ~new_new_n278__ & ~new_new_n280__;
  assign new_new_n349__ = \a[1]  & \b[8] ;
  assign new_new_n350__ = \a[2]  & \b[7] ;
  assign new_new_n351__ = \a[3]  & \b[6] ;
  assign new_new_n352__ = ~new_new_n350__ & ~new_new_n351__;
  assign new_new_n353__ = new_new_n350__ & new_new_n351__;
  assign new_new_n354__ = ~new_new_n352__ & ~new_new_n353__;
  assign new_new_n355__ = new_new_n349__ & new_new_n354__;
  assign new_new_n356__ = ~new_new_n349__ & ~new_new_n354__;
  assign new_new_n357__ = ~new_new_n355__ & ~new_new_n356__;
  assign new_new_n358__ = ~new_new_n295__ & ~new_new_n297__;
  assign new_new_n359__ = new_new_n357__ & ~new_new_n358__;
  assign new_new_n360__ = ~new_new_n357__ & new_new_n358__;
  assign new_new_n361__ = ~new_new_n359__ & ~new_new_n360__;
  assign new_new_n362__ = ~new_new_n348__ & new_new_n361__;
  assign new_new_n363__ = new_new_n348__ & ~new_new_n361__;
  assign new_new_n364__ = ~new_new_n362__ & ~new_new_n363__;
  assign new_new_n365__ = ~new_new_n310__ & ~new_new_n313__;
  assign new_new_n366__ = \a[4]  & \b[5] ;
  assign new_new_n367__ = \a[5]  & \b[4] ;
  assign new_new_n368__ = \a[7]  & \b[2] ;
  assign new_new_n369__ = ~new_new_n367__ & ~new_new_n368__;
  assign new_new_n370__ = new_new_n367__ & new_new_n368__;
  assign new_new_n371__ = ~new_new_n369__ & ~new_new_n370__;
  assign new_new_n372__ = new_new_n366__ & new_new_n371__;
  assign new_new_n373__ = ~new_new_n366__ & ~new_new_n371__;
  assign new_new_n374__ = ~new_new_n372__ & ~new_new_n373__;
  assign new_new_n375__ = ~new_new_n305__ & ~new_new_n307__;
  assign new_new_n376__ = \a[8]  & \b[1] ;
  assign new_new_n377__ = \a[6]  & \b[3] ;
  assign new_new_n378__ = \a[9]  & \b[0] ;
  assign new_new_n379__ = ~new_new_n377__ & ~new_new_n378__;
  assign new_new_n380__ = new_new_n377__ & new_new_n378__;
  assign new_new_n381__ = ~new_new_n379__ & ~new_new_n380__;
  assign new_new_n382__ = new_new_n376__ & new_new_n381__;
  assign new_new_n383__ = ~new_new_n376__ & ~new_new_n381__;
  assign new_new_n384__ = ~new_new_n382__ & ~new_new_n383__;
  assign new_new_n385__ = ~new_new_n375__ & new_new_n384__;
  assign new_new_n386__ = new_new_n375__ & ~new_new_n384__;
  assign new_new_n387__ = ~new_new_n385__ & ~new_new_n386__;
  assign new_new_n388__ = new_new_n374__ & new_new_n387__;
  assign new_new_n389__ = ~new_new_n374__ & ~new_new_n387__;
  assign new_new_n390__ = ~new_new_n388__ & ~new_new_n389__;
  assign new_new_n391__ = ~new_new_n365__ & new_new_n390__;
  assign new_new_n392__ = new_new_n365__ & ~new_new_n390__;
  assign new_new_n393__ = ~new_new_n391__ & ~new_new_n392__;
  assign new_new_n394__ = new_new_n364__ & new_new_n393__;
  assign new_new_n395__ = ~new_new_n364__ & ~new_new_n393__;
  assign new_new_n396__ = ~new_new_n394__ & ~new_new_n395__;
  assign new_new_n397__ = ~new_new_n347__ & new_new_n396__;
  assign new_new_n398__ = new_new_n347__ & ~new_new_n396__;
  assign new_new_n399__ = ~new_new_n397__ & ~new_new_n398__;
  assign new_new_n400__ = new_new_n346__ & new_new_n399__;
  assign new_new_n401__ = ~new_new_n346__ & ~new_new_n399__;
  assign new_new_n402__ = ~new_new_n400__ & ~new_new_n401__;
  assign new_new_n403__ = ~new_new_n341__ & new_new_n402__;
  assign new_new_n404__ = new_new_n341__ & ~new_new_n402__;
  assign new_new_n405__ = ~new_new_n403__ & ~new_new_n404__;
  assign new_new_n406__ = ~new_new_n329__ & ~new_new_n331__;
  assign new_new_n407__ = new_new_n405__ & new_new_n406__;
  assign new_new_n408__ = ~new_new_n405__ & ~new_new_n406__;
  assign new_new_n409__ = ~new_new_n407__ & ~new_new_n408__;
  assign new_new_n410__ = new_new_n335__ & ~new_new_n409__;
  assign new_new_n411__ = ~new_new_n335__ & new_new_n409__;
  assign new_new_n412__ = ~new_new_n338__ & new_new_n411__;
  assign new_new_n413__ = new_new_n338__ & ~new_new_n409__;
  assign new_new_n414__ = ~new_new_n410__ & ~new_new_n412__;
  assign \r[9]  = ~new_new_n413__ & new_new_n414__;
  assign new_new_n416__ = new_new_n331__ & new_new_n405__;
  assign new_new_n417__ = ~new_new_n410__ & ~new_new_n416__;
  assign new_new_n418__ = ~new_new_n413__ & new_new_n417__;
  assign new_new_n419__ = ~new_new_n397__ & ~new_new_n400__;
  assign new_new_n420__ = \a[0]  & \b[10] ;
  assign new_new_n421__ = \a[1]  & \b[9] ;
  assign new_new_n422__ = ~new_new_n420__ & ~new_new_n421__;
  assign new_new_n423__ = new_new_n420__ & new_new_n421__;
  assign new_new_n424__ = ~new_new_n422__ & ~new_new_n423__;
  assign new_new_n425__ = ~new_new_n359__ & ~new_new_n362__;
  assign new_new_n426__ = new_new_n424__ & ~new_new_n425__;
  assign new_new_n427__ = ~new_new_n424__ & new_new_n425__;
  assign new_new_n428__ = ~new_new_n426__ & ~new_new_n427__;
  assign new_new_n429__ = ~new_new_n391__ & ~new_new_n394__;
  assign new_new_n430__ = ~new_new_n353__ & ~new_new_n355__;
  assign new_new_n431__ = \a[2]  & \b[8] ;
  assign new_new_n432__ = \a[3]  & \b[7] ;
  assign new_new_n433__ = \a[4]  & \b[6] ;
  assign new_new_n434__ = ~new_new_n432__ & ~new_new_n433__;
  assign new_new_n435__ = new_new_n432__ & new_new_n433__;
  assign new_new_n436__ = ~new_new_n434__ & ~new_new_n435__;
  assign new_new_n437__ = ~new_new_n431__ & ~new_new_n436__;
  assign new_new_n438__ = new_new_n431__ & new_new_n436__;
  assign new_new_n439__ = ~new_new_n437__ & ~new_new_n438__;
  assign new_new_n440__ = ~new_new_n370__ & ~new_new_n372__;
  assign new_new_n441__ = new_new_n439__ & ~new_new_n440__;
  assign new_new_n442__ = ~new_new_n439__ & new_new_n440__;
  assign new_new_n443__ = ~new_new_n441__ & ~new_new_n442__;
  assign new_new_n444__ = ~new_new_n430__ & new_new_n443__;
  assign new_new_n445__ = new_new_n430__ & ~new_new_n443__;
  assign new_new_n446__ = ~new_new_n444__ & ~new_new_n445__;
  assign new_new_n447__ = ~new_new_n385__ & ~new_new_n388__;
  assign new_new_n448__ = \a[5]  & \b[5] ;
  assign new_new_n449__ = \a[6]  & \b[4] ;
  assign new_new_n450__ = \a[8]  & \b[2] ;
  assign new_new_n451__ = ~new_new_n449__ & ~new_new_n450__;
  assign new_new_n452__ = new_new_n449__ & new_new_n450__;
  assign new_new_n453__ = ~new_new_n451__ & ~new_new_n452__;
  assign new_new_n454__ = new_new_n448__ & new_new_n453__;
  assign new_new_n455__ = ~new_new_n448__ & ~new_new_n453__;
  assign new_new_n456__ = ~new_new_n454__ & ~new_new_n455__;
  assign new_new_n457__ = ~new_new_n380__ & ~new_new_n382__;
  assign new_new_n458__ = \a[9]  & \b[1] ;
  assign new_new_n459__ = \a[7]  & \b[3] ;
  assign new_new_n460__ = \a[10]  & \b[0] ;
  assign new_new_n461__ = ~new_new_n459__ & ~new_new_n460__;
  assign new_new_n462__ = new_new_n459__ & new_new_n460__;
  assign new_new_n463__ = ~new_new_n461__ & ~new_new_n462__;
  assign new_new_n464__ = new_new_n458__ & new_new_n463__;
  assign new_new_n465__ = ~new_new_n458__ & ~new_new_n463__;
  assign new_new_n466__ = ~new_new_n464__ & ~new_new_n465__;
  assign new_new_n467__ = ~new_new_n457__ & new_new_n466__;
  assign new_new_n468__ = new_new_n457__ & ~new_new_n466__;
  assign new_new_n469__ = ~new_new_n467__ & ~new_new_n468__;
  assign new_new_n470__ = new_new_n456__ & new_new_n469__;
  assign new_new_n471__ = ~new_new_n456__ & ~new_new_n469__;
  assign new_new_n472__ = ~new_new_n470__ & ~new_new_n471__;
  assign new_new_n473__ = ~new_new_n447__ & new_new_n472__;
  assign new_new_n474__ = new_new_n447__ & ~new_new_n472__;
  assign new_new_n475__ = ~new_new_n473__ & ~new_new_n474__;
  assign new_new_n476__ = new_new_n446__ & new_new_n475__;
  assign new_new_n477__ = ~new_new_n446__ & ~new_new_n475__;
  assign new_new_n478__ = ~new_new_n476__ & ~new_new_n477__;
  assign new_new_n479__ = ~new_new_n429__ & new_new_n478__;
  assign new_new_n480__ = new_new_n429__ & ~new_new_n478__;
  assign new_new_n481__ = ~new_new_n479__ & ~new_new_n480__;
  assign new_new_n482__ = new_new_n428__ & new_new_n481__;
  assign new_new_n483__ = ~new_new_n428__ & ~new_new_n481__;
  assign new_new_n484__ = ~new_new_n482__ & ~new_new_n483__;
  assign new_new_n485__ = ~new_new_n419__ & new_new_n484__;
  assign new_new_n486__ = new_new_n419__ & ~new_new_n484__;
  assign new_new_n487__ = ~new_new_n485__ & ~new_new_n486__;
  assign new_new_n488__ = new_new_n344__ & new_new_n487__;
  assign new_new_n489__ = ~new_new_n344__ & ~new_new_n487__;
  assign new_new_n490__ = ~new_new_n488__ & ~new_new_n489__;
  assign new_new_n491__ = new_new_n329__ & new_new_n405__;
  assign new_new_n492__ = ~new_new_n403__ & ~new_new_n491__;
  assign new_new_n493__ = new_new_n490__ & new_new_n492__;
  assign new_new_n494__ = ~new_new_n490__ & ~new_new_n492__;
  assign new_new_n495__ = ~new_new_n493__ & ~new_new_n494__;
  assign new_new_n496__ = ~new_new_n418__ & ~new_new_n495__;
  assign new_new_n497__ = new_new_n418__ & new_new_n495__;
  assign \r[10]  = ~new_new_n496__ & ~new_new_n497__;
  assign new_new_n499__ = new_new_n490__ & new_new_n491__;
  assign new_new_n500__ = ~new_new_n496__ & ~new_new_n499__;
  assign new_new_n501__ = new_new_n403__ & new_new_n490__;
  assign new_new_n502__ = ~new_new_n485__ & ~new_new_n488__;
  assign new_new_n503__ = ~new_new_n479__ & ~new_new_n482__;
  assign new_new_n504__ = \a[0]  & \b[11] ;
  assign new_new_n505__ = \a[1]  & \b[10] ;
  assign new_new_n506__ = \a[2]  & \b[9] ;
  assign new_new_n507__ = ~new_new_n505__ & ~new_new_n506__;
  assign new_new_n508__ = new_new_n505__ & new_new_n506__;
  assign new_new_n509__ = ~new_new_n507__ & ~new_new_n508__;
  assign new_new_n510__ = new_new_n504__ & new_new_n509__;
  assign new_new_n511__ = ~new_new_n504__ & ~new_new_n509__;
  assign new_new_n512__ = ~new_new_n510__ & ~new_new_n511__;
  assign new_new_n513__ = new_new_n423__ & new_new_n512__;
  assign new_new_n514__ = ~new_new_n423__ & ~new_new_n512__;
  assign new_new_n515__ = ~new_new_n513__ & ~new_new_n514__;
  assign new_new_n516__ = ~new_new_n441__ & ~new_new_n444__;
  assign new_new_n517__ = new_new_n515__ & ~new_new_n516__;
  assign new_new_n518__ = ~new_new_n515__ & new_new_n516__;
  assign new_new_n519__ = ~new_new_n517__ & ~new_new_n518__;
  assign new_new_n520__ = ~new_new_n473__ & ~new_new_n476__;
  assign new_new_n521__ = ~new_new_n435__ & ~new_new_n438__;
  assign new_new_n522__ = \a[3]  & \b[8] ;
  assign new_new_n523__ = \a[4]  & \b[7] ;
  assign new_new_n524__ = \a[5]  & \b[6] ;
  assign new_new_n525__ = ~new_new_n523__ & ~new_new_n524__;
  assign new_new_n526__ = new_new_n523__ & new_new_n524__;
  assign new_new_n527__ = ~new_new_n525__ & ~new_new_n526__;
  assign new_new_n528__ = ~new_new_n522__ & ~new_new_n527__;
  assign new_new_n529__ = new_new_n522__ & new_new_n527__;
  assign new_new_n530__ = ~new_new_n528__ & ~new_new_n529__;
  assign new_new_n531__ = ~new_new_n452__ & ~new_new_n454__;
  assign new_new_n532__ = new_new_n530__ & ~new_new_n531__;
  assign new_new_n533__ = ~new_new_n530__ & new_new_n531__;
  assign new_new_n534__ = ~new_new_n532__ & ~new_new_n533__;
  assign new_new_n535__ = ~new_new_n521__ & new_new_n534__;
  assign new_new_n536__ = new_new_n521__ & ~new_new_n534__;
  assign new_new_n537__ = ~new_new_n535__ & ~new_new_n536__;
  assign new_new_n538__ = ~new_new_n467__ & ~new_new_n470__;
  assign new_new_n539__ = \a[6]  & \b[5] ;
  assign new_new_n540__ = \a[7]  & \b[4] ;
  assign new_new_n541__ = \a[9]  & \b[2] ;
  assign new_new_n542__ = ~new_new_n540__ & ~new_new_n541__;
  assign new_new_n543__ = new_new_n540__ & new_new_n541__;
  assign new_new_n544__ = ~new_new_n542__ & ~new_new_n543__;
  assign new_new_n545__ = new_new_n539__ & new_new_n544__;
  assign new_new_n546__ = ~new_new_n539__ & ~new_new_n544__;
  assign new_new_n547__ = ~new_new_n545__ & ~new_new_n546__;
  assign new_new_n548__ = ~new_new_n462__ & ~new_new_n464__;
  assign new_new_n549__ = \a[10]  & \b[1] ;
  assign new_new_n550__ = \a[8]  & \b[3] ;
  assign new_new_n551__ = \a[11]  & \b[0] ;
  assign new_new_n552__ = ~new_new_n550__ & ~new_new_n551__;
  assign new_new_n553__ = new_new_n550__ & new_new_n551__;
  assign new_new_n554__ = ~new_new_n552__ & ~new_new_n553__;
  assign new_new_n555__ = new_new_n549__ & new_new_n554__;
  assign new_new_n556__ = ~new_new_n549__ & ~new_new_n554__;
  assign new_new_n557__ = ~new_new_n555__ & ~new_new_n556__;
  assign new_new_n558__ = ~new_new_n548__ & new_new_n557__;
  assign new_new_n559__ = new_new_n548__ & ~new_new_n557__;
  assign new_new_n560__ = ~new_new_n558__ & ~new_new_n559__;
  assign new_new_n561__ = new_new_n547__ & new_new_n560__;
  assign new_new_n562__ = ~new_new_n547__ & ~new_new_n560__;
  assign new_new_n563__ = ~new_new_n561__ & ~new_new_n562__;
  assign new_new_n564__ = ~new_new_n538__ & new_new_n563__;
  assign new_new_n565__ = new_new_n538__ & ~new_new_n563__;
  assign new_new_n566__ = ~new_new_n564__ & ~new_new_n565__;
  assign new_new_n567__ = new_new_n537__ & new_new_n566__;
  assign new_new_n568__ = ~new_new_n537__ & ~new_new_n566__;
  assign new_new_n569__ = ~new_new_n567__ & ~new_new_n568__;
  assign new_new_n570__ = ~new_new_n520__ & new_new_n569__;
  assign new_new_n571__ = new_new_n520__ & ~new_new_n569__;
  assign new_new_n572__ = ~new_new_n570__ & ~new_new_n571__;
  assign new_new_n573__ = new_new_n519__ & new_new_n572__;
  assign new_new_n574__ = ~new_new_n519__ & ~new_new_n572__;
  assign new_new_n575__ = ~new_new_n573__ & ~new_new_n574__;
  assign new_new_n576__ = ~new_new_n503__ & new_new_n575__;
  assign new_new_n577__ = new_new_n503__ & ~new_new_n575__;
  assign new_new_n578__ = ~new_new_n576__ & ~new_new_n577__;
  assign new_new_n579__ = new_new_n426__ & new_new_n578__;
  assign new_new_n580__ = ~new_new_n426__ & ~new_new_n578__;
  assign new_new_n581__ = ~new_new_n579__ & ~new_new_n580__;
  assign new_new_n582__ = new_new_n502__ & ~new_new_n581__;
  assign new_new_n583__ = ~new_new_n502__ & new_new_n581__;
  assign new_new_n584__ = ~new_new_n582__ & ~new_new_n583__;
  assign new_new_n585__ = new_new_n501__ & new_new_n584__;
  assign new_new_n586__ = ~new_new_n501__ & ~new_new_n584__;
  assign new_new_n587__ = ~new_new_n585__ & ~new_new_n586__;
  assign new_new_n588__ = new_new_n500__ & new_new_n587__;
  assign new_new_n589__ = ~new_new_n500__ & ~new_new_n587__;
  assign \r[11]  = new_new_n588__ | new_new_n589__;
  assign new_new_n591__ = ~new_new_n576__ & ~new_new_n579__;
  assign new_new_n592__ = ~new_new_n570__ & ~new_new_n573__;
  assign new_new_n593__ = \a[0]  & \b[12] ;
  assign new_new_n594__ = ~new_new_n508__ & ~new_new_n510__;
  assign new_new_n595__ = \a[1]  & \b[11] ;
  assign new_new_n596__ = \a[2]  & \b[10] ;
  assign new_new_n597__ = \a[3]  & \b[9] ;
  assign new_new_n598__ = ~new_new_n596__ & ~new_new_n597__;
  assign new_new_n599__ = new_new_n596__ & new_new_n597__;
  assign new_new_n600__ = ~new_new_n598__ & ~new_new_n599__;
  assign new_new_n601__ = new_new_n595__ & new_new_n600__;
  assign new_new_n602__ = ~new_new_n595__ & ~new_new_n600__;
  assign new_new_n603__ = ~new_new_n601__ & ~new_new_n602__;
  assign new_new_n604__ = ~new_new_n594__ & new_new_n603__;
  assign new_new_n605__ = new_new_n594__ & ~new_new_n603__;
  assign new_new_n606__ = ~new_new_n604__ & ~new_new_n605__;
  assign new_new_n607__ = ~new_new_n593__ & ~new_new_n606__;
  assign new_new_n608__ = new_new_n593__ & new_new_n606__;
  assign new_new_n609__ = ~new_new_n607__ & ~new_new_n608__;
  assign new_new_n610__ = ~new_new_n532__ & ~new_new_n535__;
  assign new_new_n611__ = new_new_n609__ & ~new_new_n610__;
  assign new_new_n612__ = ~new_new_n609__ & new_new_n610__;
  assign new_new_n613__ = ~new_new_n611__ & ~new_new_n612__;
  assign new_new_n614__ = new_new_n513__ & new_new_n613__;
  assign new_new_n615__ = ~new_new_n513__ & ~new_new_n613__;
  assign new_new_n616__ = ~new_new_n614__ & ~new_new_n615__;
  assign new_new_n617__ = ~new_new_n564__ & ~new_new_n567__;
  assign new_new_n618__ = ~new_new_n526__ & ~new_new_n529__;
  assign new_new_n619__ = \a[4]  & \b[8] ;
  assign new_new_n620__ = \a[5]  & \b[7] ;
  assign new_new_n621__ = \a[6]  & \b[6] ;
  assign new_new_n622__ = ~new_new_n620__ & ~new_new_n621__;
  assign new_new_n623__ = new_new_n620__ & new_new_n621__;
  assign new_new_n624__ = ~new_new_n622__ & ~new_new_n623__;
  assign new_new_n625__ = ~new_new_n619__ & ~new_new_n624__;
  assign new_new_n626__ = new_new_n619__ & new_new_n624__;
  assign new_new_n627__ = ~new_new_n625__ & ~new_new_n626__;
  assign new_new_n628__ = ~new_new_n543__ & ~new_new_n545__;
  assign new_new_n629__ = ~new_new_n627__ & new_new_n628__;
  assign new_new_n630__ = new_new_n627__ & ~new_new_n628__;
  assign new_new_n631__ = ~new_new_n629__ & ~new_new_n630__;
  assign new_new_n632__ = ~new_new_n618__ & new_new_n631__;
  assign new_new_n633__ = new_new_n618__ & ~new_new_n631__;
  assign new_new_n634__ = ~new_new_n632__ & ~new_new_n633__;
  assign new_new_n635__ = ~new_new_n558__ & ~new_new_n561__;
  assign new_new_n636__ = \a[7]  & \b[5] ;
  assign new_new_n637__ = \a[8]  & \b[4] ;
  assign new_new_n638__ = \a[10]  & \b[2] ;
  assign new_new_n639__ = ~new_new_n637__ & ~new_new_n638__;
  assign new_new_n640__ = new_new_n637__ & new_new_n638__;
  assign new_new_n641__ = ~new_new_n639__ & ~new_new_n640__;
  assign new_new_n642__ = new_new_n636__ & new_new_n641__;
  assign new_new_n643__ = ~new_new_n636__ & ~new_new_n641__;
  assign new_new_n644__ = ~new_new_n642__ & ~new_new_n643__;
  assign new_new_n645__ = ~new_new_n553__ & ~new_new_n555__;
  assign new_new_n646__ = \a[11]  & \b[1] ;
  assign new_new_n647__ = \a[9]  & \b[3] ;
  assign new_new_n648__ = \a[12]  & \b[0] ;
  assign new_new_n649__ = ~new_new_n647__ & ~new_new_n648__;
  assign new_new_n650__ = new_new_n647__ & new_new_n648__;
  assign new_new_n651__ = ~new_new_n649__ & ~new_new_n650__;
  assign new_new_n652__ = new_new_n646__ & new_new_n651__;
  assign new_new_n653__ = ~new_new_n646__ & ~new_new_n651__;
  assign new_new_n654__ = ~new_new_n652__ & ~new_new_n653__;
  assign new_new_n655__ = ~new_new_n645__ & new_new_n654__;
  assign new_new_n656__ = new_new_n645__ & ~new_new_n654__;
  assign new_new_n657__ = ~new_new_n655__ & ~new_new_n656__;
  assign new_new_n658__ = new_new_n644__ & new_new_n657__;
  assign new_new_n659__ = ~new_new_n644__ & ~new_new_n657__;
  assign new_new_n660__ = ~new_new_n658__ & ~new_new_n659__;
  assign new_new_n661__ = ~new_new_n635__ & new_new_n660__;
  assign new_new_n662__ = new_new_n635__ & ~new_new_n660__;
  assign new_new_n663__ = ~new_new_n661__ & ~new_new_n662__;
  assign new_new_n664__ = new_new_n634__ & new_new_n663__;
  assign new_new_n665__ = ~new_new_n634__ & ~new_new_n663__;
  assign new_new_n666__ = ~new_new_n664__ & ~new_new_n665__;
  assign new_new_n667__ = ~new_new_n617__ & new_new_n666__;
  assign new_new_n668__ = new_new_n617__ & ~new_new_n666__;
  assign new_new_n669__ = ~new_new_n667__ & ~new_new_n668__;
  assign new_new_n670__ = new_new_n616__ & new_new_n669__;
  assign new_new_n671__ = ~new_new_n616__ & ~new_new_n669__;
  assign new_new_n672__ = ~new_new_n670__ & ~new_new_n671__;
  assign new_new_n673__ = ~new_new_n592__ & new_new_n672__;
  assign new_new_n674__ = new_new_n592__ & ~new_new_n672__;
  assign new_new_n675__ = ~new_new_n673__ & ~new_new_n674__;
  assign new_new_n676__ = new_new_n517__ & new_new_n675__;
  assign new_new_n677__ = ~new_new_n517__ & ~new_new_n675__;
  assign new_new_n678__ = ~new_new_n676__ & ~new_new_n677__;
  assign new_new_n679__ = new_new_n591__ & ~new_new_n678__;
  assign new_new_n680__ = ~new_new_n591__ & new_new_n678__;
  assign new_new_n681__ = ~new_new_n679__ & ~new_new_n680__;
  assign new_new_n682__ = new_new_n583__ & new_new_n681__;
  assign new_new_n683__ = ~new_new_n583__ & ~new_new_n681__;
  assign new_new_n684__ = ~new_new_n682__ & ~new_new_n683__;
  assign new_new_n685__ = ~new_new_n495__ & new_new_n584__;
  assign new_new_n686__ = ~new_new_n418__ & new_new_n685__;
  assign new_new_n687__ = ~new_new_n499__ & ~new_new_n585__;
  assign new_new_n688__ = ~new_new_n586__ & ~new_new_n687__;
  assign new_new_n689__ = ~new_new_n686__ & ~new_new_n688__;
  assign new_new_n690__ = new_new_n684__ & ~new_new_n689__;
  assign new_new_n691__ = ~new_new_n684__ & new_new_n689__;
  assign \r[12]  = ~new_new_n690__ & ~new_new_n691__;
  assign new_new_n693__ = ~new_new_n682__ & ~new_new_n690__;
  assign new_new_n694__ = ~new_new_n673__ & ~new_new_n676__;
  assign new_new_n695__ = ~new_new_n611__ & ~new_new_n614__;
  assign new_new_n696__ = ~new_new_n667__ & ~new_new_n670__;
  assign new_new_n697__ = ~new_new_n604__ & ~new_new_n608__;
  assign new_new_n698__ = \a[0]  & \b[13] ;
  assign new_new_n699__ = \a[1]  & \b[12] ;
  assign new_new_n700__ = ~new_new_n698__ & ~new_new_n699__;
  assign new_new_n701__ = new_new_n698__ & new_new_n699__;
  assign new_new_n702__ = ~new_new_n700__ & ~new_new_n701__;
  assign new_new_n703__ = ~new_new_n599__ & ~new_new_n601__;
  assign new_new_n704__ = \a[2]  & \b[11] ;
  assign new_new_n705__ = \a[3]  & \b[10] ;
  assign new_new_n706__ = \a[4]  & \b[9] ;
  assign new_new_n707__ = ~new_new_n705__ & ~new_new_n706__;
  assign new_new_n708__ = new_new_n705__ & new_new_n706__;
  assign new_new_n709__ = ~new_new_n707__ & ~new_new_n708__;
  assign new_new_n710__ = new_new_n704__ & new_new_n709__;
  assign new_new_n711__ = ~new_new_n704__ & ~new_new_n709__;
  assign new_new_n712__ = ~new_new_n710__ & ~new_new_n711__;
  assign new_new_n713__ = ~new_new_n703__ & new_new_n712__;
  assign new_new_n714__ = new_new_n703__ & ~new_new_n712__;
  assign new_new_n715__ = ~new_new_n713__ & ~new_new_n714__;
  assign new_new_n716__ = ~new_new_n702__ & ~new_new_n715__;
  assign new_new_n717__ = new_new_n702__ & new_new_n715__;
  assign new_new_n718__ = ~new_new_n716__ & ~new_new_n717__;
  assign new_new_n719__ = ~new_new_n630__ & ~new_new_n632__;
  assign new_new_n720__ = new_new_n718__ & ~new_new_n719__;
  assign new_new_n721__ = ~new_new_n718__ & new_new_n719__;
  assign new_new_n722__ = ~new_new_n720__ & ~new_new_n721__;
  assign new_new_n723__ = ~new_new_n697__ & new_new_n722__;
  assign new_new_n724__ = new_new_n697__ & ~new_new_n722__;
  assign new_new_n725__ = ~new_new_n723__ & ~new_new_n724__;
  assign new_new_n726__ = ~new_new_n661__ & ~new_new_n664__;
  assign new_new_n727__ = ~new_new_n623__ & ~new_new_n626__;
  assign new_new_n728__ = \a[5]  & \b[8] ;
  assign new_new_n729__ = \a[6]  & \b[7] ;
  assign new_new_n730__ = \a[7]  & \b[6] ;
  assign new_new_n731__ = ~new_new_n729__ & ~new_new_n730__;
  assign new_new_n732__ = new_new_n729__ & new_new_n730__;
  assign new_new_n733__ = ~new_new_n731__ & ~new_new_n732__;
  assign new_new_n734__ = ~new_new_n728__ & ~new_new_n733__;
  assign new_new_n735__ = new_new_n728__ & new_new_n733__;
  assign new_new_n736__ = ~new_new_n734__ & ~new_new_n735__;
  assign new_new_n737__ = ~new_new_n640__ & ~new_new_n642__;
  assign new_new_n738__ = new_new_n736__ & ~new_new_n737__;
  assign new_new_n739__ = ~new_new_n736__ & new_new_n737__;
  assign new_new_n740__ = ~new_new_n738__ & ~new_new_n739__;
  assign new_new_n741__ = ~new_new_n727__ & new_new_n740__;
  assign new_new_n742__ = new_new_n727__ & ~new_new_n740__;
  assign new_new_n743__ = ~new_new_n741__ & ~new_new_n742__;
  assign new_new_n744__ = ~new_new_n655__ & ~new_new_n658__;
  assign new_new_n745__ = \a[8]  & \b[5] ;
  assign new_new_n746__ = \a[9]  & \b[4] ;
  assign new_new_n747__ = \a[11]  & \b[2] ;
  assign new_new_n748__ = ~new_new_n746__ & ~new_new_n747__;
  assign new_new_n749__ = new_new_n746__ & new_new_n747__;
  assign new_new_n750__ = ~new_new_n748__ & ~new_new_n749__;
  assign new_new_n751__ = new_new_n745__ & new_new_n750__;
  assign new_new_n752__ = ~new_new_n745__ & ~new_new_n750__;
  assign new_new_n753__ = ~new_new_n751__ & ~new_new_n752__;
  assign new_new_n754__ = ~new_new_n650__ & ~new_new_n652__;
  assign new_new_n755__ = \a[12]  & \b[1] ;
  assign new_new_n756__ = \a[10]  & \b[3] ;
  assign new_new_n757__ = \a[13]  & \b[0] ;
  assign new_new_n758__ = ~new_new_n756__ & ~new_new_n757__;
  assign new_new_n759__ = new_new_n756__ & new_new_n757__;
  assign new_new_n760__ = ~new_new_n758__ & ~new_new_n759__;
  assign new_new_n761__ = new_new_n755__ & new_new_n760__;
  assign new_new_n762__ = ~new_new_n755__ & ~new_new_n760__;
  assign new_new_n763__ = ~new_new_n761__ & ~new_new_n762__;
  assign new_new_n764__ = ~new_new_n754__ & new_new_n763__;
  assign new_new_n765__ = new_new_n754__ & ~new_new_n763__;
  assign new_new_n766__ = ~new_new_n764__ & ~new_new_n765__;
  assign new_new_n767__ = new_new_n753__ & new_new_n766__;
  assign new_new_n768__ = ~new_new_n753__ & ~new_new_n766__;
  assign new_new_n769__ = ~new_new_n767__ & ~new_new_n768__;
  assign new_new_n770__ = ~new_new_n744__ & new_new_n769__;
  assign new_new_n771__ = new_new_n744__ & ~new_new_n769__;
  assign new_new_n772__ = ~new_new_n770__ & ~new_new_n771__;
  assign new_new_n773__ = new_new_n743__ & new_new_n772__;
  assign new_new_n774__ = ~new_new_n743__ & ~new_new_n772__;
  assign new_new_n775__ = ~new_new_n773__ & ~new_new_n774__;
  assign new_new_n776__ = ~new_new_n726__ & new_new_n775__;
  assign new_new_n777__ = new_new_n726__ & ~new_new_n775__;
  assign new_new_n778__ = ~new_new_n776__ & ~new_new_n777__;
  assign new_new_n779__ = new_new_n725__ & new_new_n778__;
  assign new_new_n780__ = ~new_new_n725__ & ~new_new_n778__;
  assign new_new_n781__ = ~new_new_n779__ & ~new_new_n780__;
  assign new_new_n782__ = ~new_new_n696__ & new_new_n781__;
  assign new_new_n783__ = new_new_n696__ & ~new_new_n781__;
  assign new_new_n784__ = ~new_new_n782__ & ~new_new_n783__;
  assign new_new_n785__ = ~new_new_n695__ & new_new_n784__;
  assign new_new_n786__ = new_new_n695__ & ~new_new_n784__;
  assign new_new_n787__ = ~new_new_n785__ & ~new_new_n786__;
  assign new_new_n788__ = new_new_n694__ & ~new_new_n787__;
  assign new_new_n789__ = ~new_new_n694__ & new_new_n787__;
  assign new_new_n790__ = ~new_new_n788__ & ~new_new_n789__;
  assign new_new_n791__ = new_new_n680__ & new_new_n790__;
  assign new_new_n792__ = ~new_new_n680__ & ~new_new_n790__;
  assign new_new_n793__ = ~new_new_n791__ & ~new_new_n792__;
  assign new_new_n794__ = new_new_n693__ & new_new_n793__;
  assign new_new_n795__ = ~new_new_n693__ & ~new_new_n793__;
  assign \r[13]  = new_new_n794__ | new_new_n795__;
  assign new_new_n797__ = new_new_n684__ & new_new_n793__;
  assign new_new_n798__ = ~new_new_n689__ & new_new_n797__;
  assign new_new_n799__ = ~new_new_n680__ & ~new_new_n682__;
  assign new_new_n800__ = new_new_n790__ & ~new_new_n799__;
  assign new_new_n801__ = ~new_new_n798__ & ~new_new_n800__;
  assign new_new_n802__ = ~new_new_n782__ & ~new_new_n785__;
  assign new_new_n803__ = ~new_new_n720__ & ~new_new_n723__;
  assign new_new_n804__ = new_new_n701__ & ~new_new_n803__;
  assign new_new_n805__ = ~new_new_n701__ & new_new_n803__;
  assign new_new_n806__ = ~new_new_n804__ & ~new_new_n805__;
  assign new_new_n807__ = ~new_new_n776__ & ~new_new_n779__;
  assign new_new_n808__ = ~new_new_n713__ & ~new_new_n717__;
  assign new_new_n809__ = \a[0]  & \b[14] ;
  assign new_new_n810__ = \a[1]  & \b[13] ;
  assign new_new_n811__ = \a[2]  & \b[12] ;
  assign new_new_n812__ = ~new_new_n810__ & ~new_new_n811__;
  assign new_new_n813__ = new_new_n810__ & new_new_n811__;
  assign new_new_n814__ = ~new_new_n812__ & ~new_new_n813__;
  assign new_new_n815__ = new_new_n809__ & new_new_n814__;
  assign new_new_n816__ = ~new_new_n809__ & ~new_new_n814__;
  assign new_new_n817__ = ~new_new_n815__ & ~new_new_n816__;
  assign new_new_n818__ = ~new_new_n708__ & ~new_new_n710__;
  assign new_new_n819__ = \a[3]  & \b[11] ;
  assign new_new_n820__ = \a[4]  & \b[10] ;
  assign new_new_n821__ = \a[5]  & \b[9] ;
  assign new_new_n822__ = ~new_new_n820__ & ~new_new_n821__;
  assign new_new_n823__ = new_new_n820__ & new_new_n821__;
  assign new_new_n824__ = ~new_new_n822__ & ~new_new_n823__;
  assign new_new_n825__ = new_new_n819__ & new_new_n824__;
  assign new_new_n826__ = ~new_new_n819__ & ~new_new_n824__;
  assign new_new_n827__ = ~new_new_n825__ & ~new_new_n826__;
  assign new_new_n828__ = ~new_new_n818__ & new_new_n827__;
  assign new_new_n829__ = new_new_n818__ & ~new_new_n827__;
  assign new_new_n830__ = ~new_new_n828__ & ~new_new_n829__;
  assign new_new_n831__ = ~new_new_n817__ & ~new_new_n830__;
  assign new_new_n832__ = new_new_n817__ & new_new_n830__;
  assign new_new_n833__ = ~new_new_n831__ & ~new_new_n832__;
  assign new_new_n834__ = ~new_new_n738__ & ~new_new_n741__;
  assign new_new_n835__ = ~new_new_n833__ & new_new_n834__;
  assign new_new_n836__ = new_new_n833__ & ~new_new_n834__;
  assign new_new_n837__ = ~new_new_n835__ & ~new_new_n836__;
  assign new_new_n838__ = ~new_new_n808__ & new_new_n837__;
  assign new_new_n839__ = new_new_n808__ & ~new_new_n837__;
  assign new_new_n840__ = ~new_new_n838__ & ~new_new_n839__;
  assign new_new_n841__ = ~new_new_n770__ & ~new_new_n773__;
  assign new_new_n842__ = ~new_new_n732__ & ~new_new_n735__;
  assign new_new_n843__ = \a[6]  & \b[8] ;
  assign new_new_n844__ = \a[7]  & \b[7] ;
  assign new_new_n845__ = \a[8]  & \b[6] ;
  assign new_new_n846__ = ~new_new_n844__ & ~new_new_n845__;
  assign new_new_n847__ = new_new_n844__ & new_new_n845__;
  assign new_new_n848__ = ~new_new_n846__ & ~new_new_n847__;
  assign new_new_n849__ = ~new_new_n843__ & ~new_new_n848__;
  assign new_new_n850__ = new_new_n843__ & new_new_n848__;
  assign new_new_n851__ = ~new_new_n849__ & ~new_new_n850__;
  assign new_new_n852__ = ~new_new_n749__ & ~new_new_n751__;
  assign new_new_n853__ = new_new_n851__ & ~new_new_n852__;
  assign new_new_n854__ = ~new_new_n851__ & new_new_n852__;
  assign new_new_n855__ = ~new_new_n853__ & ~new_new_n854__;
  assign new_new_n856__ = ~new_new_n842__ & new_new_n855__;
  assign new_new_n857__ = new_new_n842__ & ~new_new_n855__;
  assign new_new_n858__ = ~new_new_n856__ & ~new_new_n857__;
  assign new_new_n859__ = ~new_new_n764__ & ~new_new_n767__;
  assign new_new_n860__ = \a[9]  & \b[5] ;
  assign new_new_n861__ = \a[10]  & \b[4] ;
  assign new_new_n862__ = \a[12]  & \b[2] ;
  assign new_new_n863__ = ~new_new_n861__ & ~new_new_n862__;
  assign new_new_n864__ = new_new_n861__ & new_new_n862__;
  assign new_new_n865__ = ~new_new_n863__ & ~new_new_n864__;
  assign new_new_n866__ = new_new_n860__ & new_new_n865__;
  assign new_new_n867__ = ~new_new_n860__ & ~new_new_n865__;
  assign new_new_n868__ = ~new_new_n866__ & ~new_new_n867__;
  assign new_new_n869__ = ~new_new_n759__ & ~new_new_n761__;
  assign new_new_n870__ = \a[13]  & \b[1] ;
  assign new_new_n871__ = \a[11]  & \b[3] ;
  assign new_new_n872__ = \a[14]  & \b[0] ;
  assign new_new_n873__ = ~new_new_n871__ & ~new_new_n872__;
  assign new_new_n874__ = new_new_n871__ & new_new_n872__;
  assign new_new_n875__ = ~new_new_n873__ & ~new_new_n874__;
  assign new_new_n876__ = new_new_n870__ & new_new_n875__;
  assign new_new_n877__ = ~new_new_n870__ & ~new_new_n875__;
  assign new_new_n878__ = ~new_new_n876__ & ~new_new_n877__;
  assign new_new_n879__ = ~new_new_n869__ & new_new_n878__;
  assign new_new_n880__ = new_new_n869__ & ~new_new_n878__;
  assign new_new_n881__ = ~new_new_n879__ & ~new_new_n880__;
  assign new_new_n882__ = new_new_n868__ & new_new_n881__;
  assign new_new_n883__ = ~new_new_n868__ & ~new_new_n881__;
  assign new_new_n884__ = ~new_new_n882__ & ~new_new_n883__;
  assign new_new_n885__ = ~new_new_n859__ & new_new_n884__;
  assign new_new_n886__ = new_new_n859__ & ~new_new_n884__;
  assign new_new_n887__ = ~new_new_n885__ & ~new_new_n886__;
  assign new_new_n888__ = new_new_n858__ & new_new_n887__;
  assign new_new_n889__ = ~new_new_n858__ & ~new_new_n887__;
  assign new_new_n890__ = ~new_new_n888__ & ~new_new_n889__;
  assign new_new_n891__ = ~new_new_n841__ & new_new_n890__;
  assign new_new_n892__ = new_new_n841__ & ~new_new_n890__;
  assign new_new_n893__ = ~new_new_n891__ & ~new_new_n892__;
  assign new_new_n894__ = new_new_n840__ & new_new_n893__;
  assign new_new_n895__ = ~new_new_n840__ & ~new_new_n893__;
  assign new_new_n896__ = ~new_new_n894__ & ~new_new_n895__;
  assign new_new_n897__ = ~new_new_n807__ & new_new_n896__;
  assign new_new_n898__ = new_new_n807__ & ~new_new_n896__;
  assign new_new_n899__ = ~new_new_n897__ & ~new_new_n898__;
  assign new_new_n900__ = new_new_n806__ & new_new_n899__;
  assign new_new_n901__ = ~new_new_n806__ & ~new_new_n899__;
  assign new_new_n902__ = ~new_new_n900__ & ~new_new_n901__;
  assign new_new_n903__ = new_new_n802__ & ~new_new_n902__;
  assign new_new_n904__ = ~new_new_n802__ & new_new_n902__;
  assign new_new_n905__ = ~new_new_n903__ & ~new_new_n904__;
  assign new_new_n906__ = new_new_n789__ & new_new_n905__;
  assign new_new_n907__ = ~new_new_n789__ & ~new_new_n905__;
  assign new_new_n908__ = ~new_new_n906__ & ~new_new_n907__;
  assign new_new_n909__ = ~new_new_n801__ & new_new_n908__;
  assign new_new_n910__ = new_new_n801__ & ~new_new_n908__;
  assign \r[14]  = ~new_new_n909__ & ~new_new_n910__;
  assign new_new_n912__ = ~new_new_n906__ & ~new_new_n909__;
  assign new_new_n913__ = ~new_new_n897__ & ~new_new_n900__;
  assign new_new_n914__ = \a[0]  & \b[15] ;
  assign new_new_n915__ = ~new_new_n813__ & ~new_new_n815__;
  assign new_new_n916__ = ~new_new_n836__ & ~new_new_n838__;
  assign new_new_n917__ = ~new_new_n915__ & ~new_new_n916__;
  assign new_new_n918__ = new_new_n915__ & new_new_n916__;
  assign new_new_n919__ = ~new_new_n917__ & ~new_new_n918__;
  assign new_new_n920__ = new_new_n914__ & new_new_n919__;
  assign new_new_n921__ = ~new_new_n914__ & ~new_new_n919__;
  assign new_new_n922__ = ~new_new_n920__ & ~new_new_n921__;
  assign new_new_n923__ = ~new_new_n891__ & ~new_new_n894__;
  assign new_new_n924__ = ~new_new_n828__ & ~new_new_n832__;
  assign new_new_n925__ = \a[1]  & \b[14] ;
  assign new_new_n926__ = \a[2]  & \b[13] ;
  assign new_new_n927__ = \a[3]  & \b[12] ;
  assign new_new_n928__ = ~new_new_n926__ & ~new_new_n927__;
  assign new_new_n929__ = new_new_n926__ & new_new_n927__;
  assign new_new_n930__ = ~new_new_n928__ & ~new_new_n929__;
  assign new_new_n931__ = new_new_n925__ & new_new_n930__;
  assign new_new_n932__ = ~new_new_n925__ & ~new_new_n930__;
  assign new_new_n933__ = ~new_new_n931__ & ~new_new_n932__;
  assign new_new_n934__ = ~new_new_n823__ & ~new_new_n825__;
  assign new_new_n935__ = \a[4]  & \b[11] ;
  assign new_new_n936__ = \a[5]  & \b[10] ;
  assign new_new_n937__ = \a[6]  & \b[9] ;
  assign new_new_n938__ = ~new_new_n936__ & ~new_new_n937__;
  assign new_new_n939__ = new_new_n936__ & new_new_n937__;
  assign new_new_n940__ = ~new_new_n938__ & ~new_new_n939__;
  assign new_new_n941__ = new_new_n935__ & new_new_n940__;
  assign new_new_n942__ = ~new_new_n935__ & ~new_new_n940__;
  assign new_new_n943__ = ~new_new_n941__ & ~new_new_n942__;
  assign new_new_n944__ = ~new_new_n934__ & new_new_n943__;
  assign new_new_n945__ = new_new_n934__ & ~new_new_n943__;
  assign new_new_n946__ = ~new_new_n944__ & ~new_new_n945__;
  assign new_new_n947__ = ~new_new_n933__ & ~new_new_n946__;
  assign new_new_n948__ = new_new_n933__ & new_new_n946__;
  assign new_new_n949__ = ~new_new_n947__ & ~new_new_n948__;
  assign new_new_n950__ = ~new_new_n853__ & ~new_new_n856__;
  assign new_new_n951__ = new_new_n949__ & ~new_new_n950__;
  assign new_new_n952__ = ~new_new_n949__ & new_new_n950__;
  assign new_new_n953__ = ~new_new_n951__ & ~new_new_n952__;
  assign new_new_n954__ = ~new_new_n924__ & new_new_n953__;
  assign new_new_n955__ = new_new_n924__ & ~new_new_n953__;
  assign new_new_n956__ = ~new_new_n954__ & ~new_new_n955__;
  assign new_new_n957__ = ~new_new_n885__ & ~new_new_n888__;
  assign new_new_n958__ = ~new_new_n847__ & ~new_new_n850__;
  assign new_new_n959__ = \a[7]  & \b[8] ;
  assign new_new_n960__ = \a[8]  & \b[7] ;
  assign new_new_n961__ = \a[9]  & \b[6] ;
  assign new_new_n962__ = ~new_new_n960__ & ~new_new_n961__;
  assign new_new_n963__ = new_new_n960__ & new_new_n961__;
  assign new_new_n964__ = ~new_new_n962__ & ~new_new_n963__;
  assign new_new_n965__ = ~new_new_n959__ & ~new_new_n964__;
  assign new_new_n966__ = new_new_n959__ & new_new_n964__;
  assign new_new_n967__ = ~new_new_n965__ & ~new_new_n966__;
  assign new_new_n968__ = ~new_new_n864__ & ~new_new_n866__;
  assign new_new_n969__ = new_new_n967__ & ~new_new_n968__;
  assign new_new_n970__ = ~new_new_n967__ & new_new_n968__;
  assign new_new_n971__ = ~new_new_n969__ & ~new_new_n970__;
  assign new_new_n972__ = ~new_new_n958__ & new_new_n971__;
  assign new_new_n973__ = new_new_n958__ & ~new_new_n971__;
  assign new_new_n974__ = ~new_new_n972__ & ~new_new_n973__;
  assign new_new_n975__ = ~new_new_n879__ & ~new_new_n882__;
  assign new_new_n976__ = \a[10]  & \b[5] ;
  assign new_new_n977__ = \a[11]  & \b[4] ;
  assign new_new_n978__ = \a[13]  & \b[2] ;
  assign new_new_n979__ = ~new_new_n977__ & ~new_new_n978__;
  assign new_new_n980__ = new_new_n977__ & new_new_n978__;
  assign new_new_n981__ = ~new_new_n979__ & ~new_new_n980__;
  assign new_new_n982__ = new_new_n976__ & new_new_n981__;
  assign new_new_n983__ = ~new_new_n976__ & ~new_new_n981__;
  assign new_new_n984__ = ~new_new_n982__ & ~new_new_n983__;
  assign new_new_n985__ = ~new_new_n874__ & ~new_new_n876__;
  assign new_new_n986__ = \a[14]  & \b[1] ;
  assign new_new_n987__ = \a[12]  & \b[3] ;
  assign new_new_n988__ = \a[15]  & \b[0] ;
  assign new_new_n989__ = ~new_new_n987__ & ~new_new_n988__;
  assign new_new_n990__ = new_new_n987__ & new_new_n988__;
  assign new_new_n991__ = ~new_new_n989__ & ~new_new_n990__;
  assign new_new_n992__ = new_new_n986__ & new_new_n991__;
  assign new_new_n993__ = ~new_new_n986__ & ~new_new_n991__;
  assign new_new_n994__ = ~new_new_n992__ & ~new_new_n993__;
  assign new_new_n995__ = ~new_new_n985__ & new_new_n994__;
  assign new_new_n996__ = new_new_n985__ & ~new_new_n994__;
  assign new_new_n997__ = ~new_new_n995__ & ~new_new_n996__;
  assign new_new_n998__ = new_new_n984__ & new_new_n997__;
  assign new_new_n999__ = ~new_new_n984__ & ~new_new_n997__;
  assign new_new_n1000__ = ~new_new_n998__ & ~new_new_n999__;
  assign new_new_n1001__ = ~new_new_n975__ & new_new_n1000__;
  assign new_new_n1002__ = new_new_n975__ & ~new_new_n1000__;
  assign new_new_n1003__ = ~new_new_n1001__ & ~new_new_n1002__;
  assign new_new_n1004__ = new_new_n974__ & new_new_n1003__;
  assign new_new_n1005__ = ~new_new_n974__ & ~new_new_n1003__;
  assign new_new_n1006__ = ~new_new_n1004__ & ~new_new_n1005__;
  assign new_new_n1007__ = ~new_new_n957__ & new_new_n1006__;
  assign new_new_n1008__ = new_new_n957__ & ~new_new_n1006__;
  assign new_new_n1009__ = ~new_new_n1007__ & ~new_new_n1008__;
  assign new_new_n1010__ = new_new_n956__ & new_new_n1009__;
  assign new_new_n1011__ = ~new_new_n956__ & ~new_new_n1009__;
  assign new_new_n1012__ = ~new_new_n1010__ & ~new_new_n1011__;
  assign new_new_n1013__ = ~new_new_n923__ & new_new_n1012__;
  assign new_new_n1014__ = new_new_n923__ & ~new_new_n1012__;
  assign new_new_n1015__ = ~new_new_n1013__ & ~new_new_n1014__;
  assign new_new_n1016__ = new_new_n922__ & new_new_n1015__;
  assign new_new_n1017__ = ~new_new_n922__ & ~new_new_n1015__;
  assign new_new_n1018__ = ~new_new_n1016__ & ~new_new_n1017__;
  assign new_new_n1019__ = ~new_new_n913__ & new_new_n1018__;
  assign new_new_n1020__ = new_new_n913__ & ~new_new_n1018__;
  assign new_new_n1021__ = ~new_new_n1019__ & ~new_new_n1020__;
  assign new_new_n1022__ = new_new_n804__ & new_new_n1021__;
  assign new_new_n1023__ = ~new_new_n804__ & ~new_new_n1021__;
  assign new_new_n1024__ = ~new_new_n1022__ & ~new_new_n1023__;
  assign new_new_n1025__ = new_new_n904__ & new_new_n1024__;
  assign new_new_n1026__ = ~new_new_n904__ & ~new_new_n1024__;
  assign new_new_n1027__ = ~new_new_n1025__ & ~new_new_n1026__;
  assign new_new_n1028__ = new_new_n912__ & ~new_new_n1027__;
  assign new_new_n1029__ = ~new_new_n912__ & new_new_n1027__;
  assign \r[15]  = ~new_new_n1028__ & ~new_new_n1029__;
  assign new_new_n1031__ = ~new_new_n1019__ & ~new_new_n1022__;
  assign new_new_n1032__ = ~new_new_n917__ & ~new_new_n920__;
  assign new_new_n1033__ = ~new_new_n1013__ & ~new_new_n1016__;
  assign new_new_n1034__ = \a[1]  & \b[15] ;
  assign new_new_n1035__ = ~new_new_n929__ & ~new_new_n931__;
  assign new_new_n1036__ = ~new_new_n951__ & ~new_new_n954__;
  assign new_new_n1037__ = ~new_new_n1035__ & ~new_new_n1036__;
  assign new_new_n1038__ = new_new_n1035__ & new_new_n1036__;
  assign new_new_n1039__ = ~new_new_n1037__ & ~new_new_n1038__;
  assign new_new_n1040__ = new_new_n1034__ & new_new_n1039__;
  assign new_new_n1041__ = ~new_new_n1034__ & ~new_new_n1039__;
  assign new_new_n1042__ = ~new_new_n1040__ & ~new_new_n1041__;
  assign new_new_n1043__ = ~new_new_n1007__ & ~new_new_n1010__;
  assign new_new_n1044__ = ~new_new_n1001__ & ~new_new_n1004__;
  assign new_new_n1045__ = ~new_new_n963__ & ~new_new_n966__;
  assign new_new_n1046__ = \a[8]  & \b[8] ;
  assign new_new_n1047__ = \a[9]  & \b[7] ;
  assign new_new_n1048__ = \a[10]  & \b[6] ;
  assign new_new_n1049__ = ~new_new_n1047__ & ~new_new_n1048__;
  assign new_new_n1050__ = new_new_n1047__ & new_new_n1048__;
  assign new_new_n1051__ = ~new_new_n1049__ & ~new_new_n1050__;
  assign new_new_n1052__ = ~new_new_n1046__ & ~new_new_n1051__;
  assign new_new_n1053__ = new_new_n1046__ & new_new_n1051__;
  assign new_new_n1054__ = ~new_new_n1052__ & ~new_new_n1053__;
  assign new_new_n1055__ = ~new_new_n980__ & ~new_new_n982__;
  assign new_new_n1056__ = new_new_n1054__ & ~new_new_n1055__;
  assign new_new_n1057__ = ~new_new_n1054__ & new_new_n1055__;
  assign new_new_n1058__ = ~new_new_n1056__ & ~new_new_n1057__;
  assign new_new_n1059__ = ~new_new_n1045__ & new_new_n1058__;
  assign new_new_n1060__ = new_new_n1045__ & ~new_new_n1058__;
  assign new_new_n1061__ = ~new_new_n1059__ & ~new_new_n1060__;
  assign new_new_n1062__ = ~new_new_n995__ & ~new_new_n998__;
  assign new_new_n1063__ = \a[11]  & \b[5] ;
  assign new_new_n1064__ = \a[12]  & \b[4] ;
  assign new_new_n1065__ = \a[14]  & \b[2] ;
  assign new_new_n1066__ = ~new_new_n1064__ & ~new_new_n1065__;
  assign new_new_n1067__ = new_new_n1064__ & new_new_n1065__;
  assign new_new_n1068__ = ~new_new_n1066__ & ~new_new_n1067__;
  assign new_new_n1069__ = new_new_n1063__ & new_new_n1068__;
  assign new_new_n1070__ = ~new_new_n1063__ & ~new_new_n1068__;
  assign new_new_n1071__ = ~new_new_n1069__ & ~new_new_n1070__;
  assign new_new_n1072__ = ~new_new_n990__ & ~new_new_n992__;
  assign new_new_n1073__ = \a[13]  & \b[3] ;
  assign new_new_n1074__ = \a[15]  & \b[1] ;
  assign new_new_n1075__ = ~new_new_n1073__ & ~new_new_n1074__;
  assign new_new_n1076__ = new_new_n1073__ & new_new_n1074__;
  assign new_new_n1077__ = ~new_new_n1075__ & ~new_new_n1076__;
  assign new_new_n1078__ = ~new_new_n1072__ & new_new_n1077__;
  assign new_new_n1079__ = new_new_n1072__ & ~new_new_n1077__;
  assign new_new_n1080__ = ~new_new_n1078__ & ~new_new_n1079__;
  assign new_new_n1081__ = new_new_n1071__ & new_new_n1080__;
  assign new_new_n1082__ = ~new_new_n1071__ & ~new_new_n1080__;
  assign new_new_n1083__ = ~new_new_n1081__ & ~new_new_n1082__;
  assign new_new_n1084__ = ~new_new_n1062__ & new_new_n1083__;
  assign new_new_n1085__ = new_new_n1062__ & ~new_new_n1083__;
  assign new_new_n1086__ = ~new_new_n1084__ & ~new_new_n1085__;
  assign new_new_n1087__ = new_new_n1061__ & new_new_n1086__;
  assign new_new_n1088__ = ~new_new_n1061__ & ~new_new_n1086__;
  assign new_new_n1089__ = ~new_new_n1087__ & ~new_new_n1088__;
  assign new_new_n1090__ = ~new_new_n1044__ & new_new_n1089__;
  assign new_new_n1091__ = new_new_n1044__ & ~new_new_n1089__;
  assign new_new_n1092__ = ~new_new_n1090__ & ~new_new_n1091__;
  assign new_new_n1093__ = ~new_new_n944__ & ~new_new_n948__;
  assign new_new_n1094__ = \a[2]  & \b[14] ;
  assign new_new_n1095__ = \a[3]  & \b[13] ;
  assign new_new_n1096__ = \a[4]  & \b[12] ;
  assign new_new_n1097__ = ~new_new_n1095__ & ~new_new_n1096__;
  assign new_new_n1098__ = new_new_n1095__ & new_new_n1096__;
  assign new_new_n1099__ = ~new_new_n1097__ & ~new_new_n1098__;
  assign new_new_n1100__ = new_new_n1094__ & new_new_n1099__;
  assign new_new_n1101__ = ~new_new_n1094__ & ~new_new_n1099__;
  assign new_new_n1102__ = ~new_new_n1100__ & ~new_new_n1101__;
  assign new_new_n1103__ = ~new_new_n939__ & ~new_new_n941__;
  assign new_new_n1104__ = \a[5]  & \b[11] ;
  assign new_new_n1105__ = \a[6]  & \b[10] ;
  assign new_new_n1106__ = \a[7]  & \b[9] ;
  assign new_new_n1107__ = ~new_new_n1105__ & ~new_new_n1106__;
  assign new_new_n1108__ = new_new_n1105__ & new_new_n1106__;
  assign new_new_n1109__ = ~new_new_n1107__ & ~new_new_n1108__;
  assign new_new_n1110__ = new_new_n1104__ & new_new_n1109__;
  assign new_new_n1111__ = ~new_new_n1104__ & ~new_new_n1109__;
  assign new_new_n1112__ = ~new_new_n1110__ & ~new_new_n1111__;
  assign new_new_n1113__ = ~new_new_n1103__ & new_new_n1112__;
  assign new_new_n1114__ = new_new_n1103__ & ~new_new_n1112__;
  assign new_new_n1115__ = ~new_new_n1113__ & ~new_new_n1114__;
  assign new_new_n1116__ = ~new_new_n1102__ & ~new_new_n1115__;
  assign new_new_n1117__ = new_new_n1102__ & new_new_n1115__;
  assign new_new_n1118__ = ~new_new_n1116__ & ~new_new_n1117__;
  assign new_new_n1119__ = ~new_new_n969__ & ~new_new_n972__;
  assign new_new_n1120__ = new_new_n1118__ & ~new_new_n1119__;
  assign new_new_n1121__ = ~new_new_n1118__ & new_new_n1119__;
  assign new_new_n1122__ = ~new_new_n1120__ & ~new_new_n1121__;
  assign new_new_n1123__ = ~new_new_n1093__ & new_new_n1122__;
  assign new_new_n1124__ = new_new_n1093__ & ~new_new_n1122__;
  assign new_new_n1125__ = ~new_new_n1123__ & ~new_new_n1124__;
  assign new_new_n1126__ = new_new_n1092__ & new_new_n1125__;
  assign new_new_n1127__ = ~new_new_n1092__ & ~new_new_n1125__;
  assign new_new_n1128__ = ~new_new_n1126__ & ~new_new_n1127__;
  assign new_new_n1129__ = ~new_new_n1043__ & new_new_n1128__;
  assign new_new_n1130__ = new_new_n1043__ & ~new_new_n1128__;
  assign new_new_n1131__ = ~new_new_n1129__ & ~new_new_n1130__;
  assign new_new_n1132__ = new_new_n1042__ & new_new_n1131__;
  assign new_new_n1133__ = ~new_new_n1042__ & ~new_new_n1131__;
  assign new_new_n1134__ = ~new_new_n1132__ & ~new_new_n1133__;
  assign new_new_n1135__ = ~new_new_n1033__ & new_new_n1134__;
  assign new_new_n1136__ = new_new_n1033__ & ~new_new_n1134__;
  assign new_new_n1137__ = ~new_new_n1135__ & ~new_new_n1136__;
  assign new_new_n1138__ = ~new_new_n1032__ & new_new_n1137__;
  assign new_new_n1139__ = new_new_n1032__ & ~new_new_n1137__;
  assign new_new_n1140__ = ~new_new_n1138__ & ~new_new_n1139__;
  assign new_new_n1141__ = new_new_n1031__ & ~new_new_n1140__;
  assign new_new_n1142__ = ~new_new_n1031__ & new_new_n1140__;
  assign new_new_n1143__ = ~new_new_n1141__ & ~new_new_n1142__;
  assign new_new_n1144__ = new_new_n908__ & new_new_n1027__;
  assign new_new_n1145__ = new_new_n798__ & new_new_n1144__;
  assign new_new_n1146__ = new_new_n800__ & new_new_n1144__;
  assign new_new_n1147__ = ~new_new_n904__ & ~new_new_n906__;
  assign new_new_n1148__ = new_new_n1024__ & ~new_new_n1147__;
  assign new_new_n1149__ = ~new_new_n1146__ & ~new_new_n1148__;
  assign new_new_n1150__ = ~new_new_n1145__ & new_new_n1149__;
  assign new_new_n1151__ = new_new_n1143__ & ~new_new_n1150__;
  assign new_new_n1152__ = ~new_new_n1143__ & new_new_n1150__;
  assign \r[16]  = ~new_new_n1151__ & ~new_new_n1152__;
  assign new_new_n1154__ = ~new_new_n1142__ & ~new_new_n1151__;
  assign new_new_n1155__ = ~new_new_n1135__ & ~new_new_n1138__;
  assign new_new_n1156__ = ~new_new_n1037__ & ~new_new_n1040__;
  assign new_new_n1157__ = ~new_new_n1129__ & ~new_new_n1132__;
  assign new_new_n1158__ = \a[2]  & \b[15] ;
  assign new_new_n1159__ = ~new_new_n1098__ & ~new_new_n1100__;
  assign new_new_n1160__ = ~new_new_n1120__ & ~new_new_n1123__;
  assign new_new_n1161__ = ~new_new_n1159__ & ~new_new_n1160__;
  assign new_new_n1162__ = new_new_n1159__ & new_new_n1160__;
  assign new_new_n1163__ = ~new_new_n1161__ & ~new_new_n1162__;
  assign new_new_n1164__ = new_new_n1158__ & new_new_n1163__;
  assign new_new_n1165__ = ~new_new_n1158__ & ~new_new_n1163__;
  assign new_new_n1166__ = ~new_new_n1164__ & ~new_new_n1165__;
  assign new_new_n1167__ = ~new_new_n1090__ & ~new_new_n1126__;
  assign new_new_n1168__ = ~new_new_n1084__ & ~new_new_n1087__;
  assign new_new_n1169__ = ~new_new_n1050__ & ~new_new_n1053__;
  assign new_new_n1170__ = \a[9]  & \b[8] ;
  assign new_new_n1171__ = \a[10]  & \b[7] ;
  assign new_new_n1172__ = \a[11]  & \b[6] ;
  assign new_new_n1173__ = ~new_new_n1171__ & ~new_new_n1172__;
  assign new_new_n1174__ = new_new_n1171__ & new_new_n1172__;
  assign new_new_n1175__ = ~new_new_n1173__ & ~new_new_n1174__;
  assign new_new_n1176__ = ~new_new_n1170__ & ~new_new_n1175__;
  assign new_new_n1177__ = new_new_n1170__ & new_new_n1175__;
  assign new_new_n1178__ = ~new_new_n1176__ & ~new_new_n1177__;
  assign new_new_n1179__ = ~new_new_n1067__ & ~new_new_n1069__;
  assign new_new_n1180__ = new_new_n1178__ & ~new_new_n1179__;
  assign new_new_n1181__ = ~new_new_n1178__ & new_new_n1179__;
  assign new_new_n1182__ = ~new_new_n1180__ & ~new_new_n1181__;
  assign new_new_n1183__ = ~new_new_n1169__ & new_new_n1182__;
  assign new_new_n1184__ = new_new_n1169__ & ~new_new_n1182__;
  assign new_new_n1185__ = ~new_new_n1183__ & ~new_new_n1184__;
  assign new_new_n1186__ = ~new_new_n1078__ & ~new_new_n1081__;
  assign new_new_n1187__ = \a[12]  & \b[5] ;
  assign new_new_n1188__ = \a[13]  & \b[4] ;
  assign new_new_n1189__ = \a[15]  & \b[2] ;
  assign new_new_n1190__ = ~new_new_n1188__ & ~new_new_n1189__;
  assign new_new_n1191__ = new_new_n1188__ & new_new_n1189__;
  assign new_new_n1192__ = ~new_new_n1190__ & ~new_new_n1191__;
  assign new_new_n1193__ = new_new_n1187__ & new_new_n1192__;
  assign new_new_n1194__ = ~new_new_n1187__ & ~new_new_n1192__;
  assign new_new_n1195__ = ~new_new_n1193__ & ~new_new_n1194__;
  assign new_new_n1196__ = \a[14]  & \b[3] ;
  assign new_new_n1197__ = ~new_new_n1076__ & ~new_new_n1196__;
  assign new_new_n1198__ = \a[14]  & new_new_n1076__;
  assign new_new_n1199__ = ~new_new_n1197__ & ~new_new_n1198__;
  assign new_new_n1200__ = new_new_n1195__ & new_new_n1199__;
  assign new_new_n1201__ = ~new_new_n1195__ & ~new_new_n1199__;
  assign new_new_n1202__ = ~new_new_n1200__ & ~new_new_n1201__;
  assign new_new_n1203__ = ~new_new_n1186__ & new_new_n1202__;
  assign new_new_n1204__ = new_new_n1186__ & ~new_new_n1202__;
  assign new_new_n1205__ = ~new_new_n1203__ & ~new_new_n1204__;
  assign new_new_n1206__ = new_new_n1185__ & new_new_n1205__;
  assign new_new_n1207__ = ~new_new_n1185__ & ~new_new_n1205__;
  assign new_new_n1208__ = ~new_new_n1206__ & ~new_new_n1207__;
  assign new_new_n1209__ = ~new_new_n1168__ & new_new_n1208__;
  assign new_new_n1210__ = new_new_n1168__ & ~new_new_n1208__;
  assign new_new_n1211__ = ~new_new_n1209__ & ~new_new_n1210__;
  assign new_new_n1212__ = ~new_new_n1113__ & ~new_new_n1117__;
  assign new_new_n1213__ = \a[3]  & \b[14] ;
  assign new_new_n1214__ = \a[4]  & \b[13] ;
  assign new_new_n1215__ = \a[5]  & \b[12] ;
  assign new_new_n1216__ = ~new_new_n1214__ & ~new_new_n1215__;
  assign new_new_n1217__ = new_new_n1214__ & new_new_n1215__;
  assign new_new_n1218__ = ~new_new_n1216__ & ~new_new_n1217__;
  assign new_new_n1219__ = new_new_n1213__ & new_new_n1218__;
  assign new_new_n1220__ = ~new_new_n1213__ & ~new_new_n1218__;
  assign new_new_n1221__ = ~new_new_n1219__ & ~new_new_n1220__;
  assign new_new_n1222__ = ~new_new_n1108__ & ~new_new_n1110__;
  assign new_new_n1223__ = \a[6]  & \b[11] ;
  assign new_new_n1224__ = \a[7]  & \b[10] ;
  assign new_new_n1225__ = \a[8]  & \b[9] ;
  assign new_new_n1226__ = ~new_new_n1224__ & ~new_new_n1225__;
  assign new_new_n1227__ = new_new_n1224__ & new_new_n1225__;
  assign new_new_n1228__ = ~new_new_n1226__ & ~new_new_n1227__;
  assign new_new_n1229__ = new_new_n1223__ & new_new_n1228__;
  assign new_new_n1230__ = ~new_new_n1223__ & ~new_new_n1228__;
  assign new_new_n1231__ = ~new_new_n1229__ & ~new_new_n1230__;
  assign new_new_n1232__ = ~new_new_n1222__ & new_new_n1231__;
  assign new_new_n1233__ = new_new_n1222__ & ~new_new_n1231__;
  assign new_new_n1234__ = ~new_new_n1232__ & ~new_new_n1233__;
  assign new_new_n1235__ = ~new_new_n1221__ & ~new_new_n1234__;
  assign new_new_n1236__ = new_new_n1221__ & new_new_n1234__;
  assign new_new_n1237__ = ~new_new_n1235__ & ~new_new_n1236__;
  assign new_new_n1238__ = ~new_new_n1056__ & ~new_new_n1059__;
  assign new_new_n1239__ = new_new_n1237__ & ~new_new_n1238__;
  assign new_new_n1240__ = ~new_new_n1237__ & new_new_n1238__;
  assign new_new_n1241__ = ~new_new_n1239__ & ~new_new_n1240__;
  assign new_new_n1242__ = ~new_new_n1212__ & new_new_n1241__;
  assign new_new_n1243__ = new_new_n1212__ & ~new_new_n1241__;
  assign new_new_n1244__ = ~new_new_n1242__ & ~new_new_n1243__;
  assign new_new_n1245__ = new_new_n1211__ & new_new_n1244__;
  assign new_new_n1246__ = ~new_new_n1211__ & ~new_new_n1244__;
  assign new_new_n1247__ = ~new_new_n1245__ & ~new_new_n1246__;
  assign new_new_n1248__ = ~new_new_n1167__ & new_new_n1247__;
  assign new_new_n1249__ = new_new_n1167__ & ~new_new_n1247__;
  assign new_new_n1250__ = ~new_new_n1248__ & ~new_new_n1249__;
  assign new_new_n1251__ = new_new_n1166__ & new_new_n1250__;
  assign new_new_n1252__ = ~new_new_n1166__ & ~new_new_n1250__;
  assign new_new_n1253__ = ~new_new_n1251__ & ~new_new_n1252__;
  assign new_new_n1254__ = ~new_new_n1157__ & new_new_n1253__;
  assign new_new_n1255__ = new_new_n1157__ & ~new_new_n1253__;
  assign new_new_n1256__ = ~new_new_n1254__ & ~new_new_n1255__;
  assign new_new_n1257__ = ~new_new_n1156__ & new_new_n1256__;
  assign new_new_n1258__ = new_new_n1156__ & ~new_new_n1256__;
  assign new_new_n1259__ = ~new_new_n1257__ & ~new_new_n1258__;
  assign new_new_n1260__ = ~new_new_n1155__ & new_new_n1259__;
  assign new_new_n1261__ = new_new_n1155__ & ~new_new_n1259__;
  assign new_new_n1262__ = ~new_new_n1260__ & ~new_new_n1261__;
  assign new_new_n1263__ = new_new_n1154__ & new_new_n1262__;
  assign new_new_n1264__ = ~new_new_n1154__ & ~new_new_n1262__;
  assign \r[17]  = new_new_n1263__ | new_new_n1264__;
  assign new_new_n1266__ = ~new_new_n1254__ & ~new_new_n1257__;
  assign new_new_n1267__ = ~new_new_n1161__ & ~new_new_n1164__;
  assign new_new_n1268__ = ~new_new_n1248__ & ~new_new_n1251__;
  assign new_new_n1269__ = \a[3]  & \b[15] ;
  assign new_new_n1270__ = ~new_new_n1217__ & ~new_new_n1219__;
  assign new_new_n1271__ = ~new_new_n1239__ & ~new_new_n1242__;
  assign new_new_n1272__ = ~new_new_n1270__ & ~new_new_n1271__;
  assign new_new_n1273__ = new_new_n1270__ & new_new_n1271__;
  assign new_new_n1274__ = ~new_new_n1272__ & ~new_new_n1273__;
  assign new_new_n1275__ = new_new_n1269__ & new_new_n1274__;
  assign new_new_n1276__ = ~new_new_n1269__ & ~new_new_n1274__;
  assign new_new_n1277__ = ~new_new_n1275__ & ~new_new_n1276__;
  assign new_new_n1278__ = ~new_new_n1209__ & ~new_new_n1245__;
  assign new_new_n1279__ = ~new_new_n1203__ & ~new_new_n1206__;
  assign new_new_n1280__ = ~new_new_n1174__ & ~new_new_n1177__;
  assign new_new_n1281__ = \a[10]  & \b[8] ;
  assign new_new_n1282__ = \a[11]  & \b[7] ;
  assign new_new_n1283__ = \a[12]  & \b[6] ;
  assign new_new_n1284__ = ~new_new_n1282__ & ~new_new_n1283__;
  assign new_new_n1285__ = new_new_n1282__ & new_new_n1283__;
  assign new_new_n1286__ = ~new_new_n1284__ & ~new_new_n1285__;
  assign new_new_n1287__ = ~new_new_n1281__ & ~new_new_n1286__;
  assign new_new_n1288__ = new_new_n1281__ & new_new_n1286__;
  assign new_new_n1289__ = ~new_new_n1287__ & ~new_new_n1288__;
  assign new_new_n1290__ = ~new_new_n1191__ & ~new_new_n1193__;
  assign new_new_n1291__ = new_new_n1289__ & ~new_new_n1290__;
  assign new_new_n1292__ = ~new_new_n1289__ & new_new_n1290__;
  assign new_new_n1293__ = ~new_new_n1291__ & ~new_new_n1292__;
  assign new_new_n1294__ = ~new_new_n1280__ & new_new_n1293__;
  assign new_new_n1295__ = new_new_n1280__ & ~new_new_n1293__;
  assign new_new_n1296__ = ~new_new_n1294__ & ~new_new_n1295__;
  assign new_new_n1297__ = ~new_new_n1198__ & ~new_new_n1200__;
  assign new_new_n1298__ = \a[15]  & \b[3] ;
  assign new_new_n1299__ = \a[14]  & \b[4] ;
  assign new_new_n1300__ = \a[13]  & \b[5] ;
  assign new_new_n1301__ = ~new_new_n1299__ & ~new_new_n1300__;
  assign new_new_n1302__ = new_new_n1299__ & new_new_n1300__;
  assign new_new_n1303__ = ~new_new_n1301__ & ~new_new_n1302__;
  assign new_new_n1304__ = new_new_n1298__ & new_new_n1303__;
  assign new_new_n1305__ = ~new_new_n1298__ & ~new_new_n1303__;
  assign new_new_n1306__ = ~new_new_n1304__ & ~new_new_n1305__;
  assign new_new_n1307__ = ~new_new_n1297__ & new_new_n1306__;
  assign new_new_n1308__ = new_new_n1297__ & ~new_new_n1306__;
  assign new_new_n1309__ = ~new_new_n1307__ & ~new_new_n1308__;
  assign new_new_n1310__ = new_new_n1296__ & new_new_n1309__;
  assign new_new_n1311__ = ~new_new_n1296__ & ~new_new_n1309__;
  assign new_new_n1312__ = ~new_new_n1310__ & ~new_new_n1311__;
  assign new_new_n1313__ = ~new_new_n1279__ & new_new_n1312__;
  assign new_new_n1314__ = new_new_n1279__ & ~new_new_n1312__;
  assign new_new_n1315__ = ~new_new_n1313__ & ~new_new_n1314__;
  assign new_new_n1316__ = ~new_new_n1232__ & ~new_new_n1236__;
  assign new_new_n1317__ = \a[4]  & \b[14] ;
  assign new_new_n1318__ = \a[5]  & \b[13] ;
  assign new_new_n1319__ = \a[6]  & \b[12] ;
  assign new_new_n1320__ = ~new_new_n1318__ & ~new_new_n1319__;
  assign new_new_n1321__ = new_new_n1318__ & new_new_n1319__;
  assign new_new_n1322__ = ~new_new_n1320__ & ~new_new_n1321__;
  assign new_new_n1323__ = new_new_n1317__ & new_new_n1322__;
  assign new_new_n1324__ = ~new_new_n1317__ & ~new_new_n1322__;
  assign new_new_n1325__ = ~new_new_n1323__ & ~new_new_n1324__;
  assign new_new_n1326__ = ~new_new_n1227__ & ~new_new_n1229__;
  assign new_new_n1327__ = \a[7]  & \b[11] ;
  assign new_new_n1328__ = \a[8]  & \b[10] ;
  assign new_new_n1329__ = \a[9]  & \b[9] ;
  assign new_new_n1330__ = ~new_new_n1328__ & ~new_new_n1329__;
  assign new_new_n1331__ = new_new_n1328__ & new_new_n1329__;
  assign new_new_n1332__ = ~new_new_n1330__ & ~new_new_n1331__;
  assign new_new_n1333__ = new_new_n1327__ & new_new_n1332__;
  assign new_new_n1334__ = ~new_new_n1327__ & ~new_new_n1332__;
  assign new_new_n1335__ = ~new_new_n1333__ & ~new_new_n1334__;
  assign new_new_n1336__ = ~new_new_n1326__ & new_new_n1335__;
  assign new_new_n1337__ = new_new_n1326__ & ~new_new_n1335__;
  assign new_new_n1338__ = ~new_new_n1336__ & ~new_new_n1337__;
  assign new_new_n1339__ = ~new_new_n1325__ & ~new_new_n1338__;
  assign new_new_n1340__ = new_new_n1325__ & new_new_n1338__;
  assign new_new_n1341__ = ~new_new_n1339__ & ~new_new_n1340__;
  assign new_new_n1342__ = ~new_new_n1180__ & ~new_new_n1183__;
  assign new_new_n1343__ = new_new_n1341__ & ~new_new_n1342__;
  assign new_new_n1344__ = ~new_new_n1341__ & new_new_n1342__;
  assign new_new_n1345__ = ~new_new_n1343__ & ~new_new_n1344__;
  assign new_new_n1346__ = ~new_new_n1316__ & new_new_n1345__;
  assign new_new_n1347__ = new_new_n1316__ & ~new_new_n1345__;
  assign new_new_n1348__ = ~new_new_n1346__ & ~new_new_n1347__;
  assign new_new_n1349__ = new_new_n1315__ & new_new_n1348__;
  assign new_new_n1350__ = ~new_new_n1315__ & ~new_new_n1348__;
  assign new_new_n1351__ = ~new_new_n1349__ & ~new_new_n1350__;
  assign new_new_n1352__ = ~new_new_n1278__ & new_new_n1351__;
  assign new_new_n1353__ = new_new_n1278__ & ~new_new_n1351__;
  assign new_new_n1354__ = ~new_new_n1352__ & ~new_new_n1353__;
  assign new_new_n1355__ = new_new_n1277__ & new_new_n1354__;
  assign new_new_n1356__ = ~new_new_n1277__ & ~new_new_n1354__;
  assign new_new_n1357__ = ~new_new_n1355__ & ~new_new_n1356__;
  assign new_new_n1358__ = ~new_new_n1268__ & new_new_n1357__;
  assign new_new_n1359__ = new_new_n1268__ & ~new_new_n1357__;
  assign new_new_n1360__ = ~new_new_n1358__ & ~new_new_n1359__;
  assign new_new_n1361__ = ~new_new_n1267__ & new_new_n1360__;
  assign new_new_n1362__ = new_new_n1267__ & ~new_new_n1360__;
  assign new_new_n1363__ = ~new_new_n1361__ & ~new_new_n1362__;
  assign new_new_n1364__ = ~new_new_n1266__ & new_new_n1363__;
  assign new_new_n1365__ = new_new_n1266__ & ~new_new_n1363__;
  assign new_new_n1366__ = ~new_new_n1364__ & ~new_new_n1365__;
  assign new_new_n1367__ = ~new_new_n1142__ & ~new_new_n1260__;
  assign new_new_n1368__ = ~new_new_n1261__ & ~new_new_n1367__;
  assign new_new_n1369__ = new_new_n1143__ & new_new_n1262__;
  assign new_new_n1370__ = ~new_new_n1150__ & new_new_n1369__;
  assign new_new_n1371__ = ~new_new_n1368__ & ~new_new_n1370__;
  assign new_new_n1372__ = new_new_n1366__ & ~new_new_n1371__;
  assign new_new_n1373__ = ~new_new_n1366__ & new_new_n1371__;
  assign \r[18]  = ~new_new_n1372__ & ~new_new_n1373__;
  assign new_new_n1375__ = ~new_new_n1364__ & ~new_new_n1372__;
  assign new_new_n1376__ = ~new_new_n1358__ & ~new_new_n1361__;
  assign new_new_n1377__ = ~new_new_n1272__ & ~new_new_n1275__;
  assign new_new_n1378__ = ~new_new_n1352__ & ~new_new_n1355__;
  assign new_new_n1379__ = \a[4]  & \b[15] ;
  assign new_new_n1380__ = ~new_new_n1321__ & ~new_new_n1323__;
  assign new_new_n1381__ = ~new_new_n1343__ & ~new_new_n1346__;
  assign new_new_n1382__ = ~new_new_n1380__ & ~new_new_n1381__;
  assign new_new_n1383__ = new_new_n1380__ & new_new_n1381__;
  assign new_new_n1384__ = ~new_new_n1382__ & ~new_new_n1383__;
  assign new_new_n1385__ = new_new_n1379__ & new_new_n1384__;
  assign new_new_n1386__ = ~new_new_n1379__ & ~new_new_n1384__;
  assign new_new_n1387__ = ~new_new_n1385__ & ~new_new_n1386__;
  assign new_new_n1388__ = ~new_new_n1313__ & ~new_new_n1349__;
  assign new_new_n1389__ = ~new_new_n1307__ & ~new_new_n1310__;
  assign new_new_n1390__ = ~new_new_n1285__ & ~new_new_n1288__;
  assign new_new_n1391__ = \a[11]  & \b[8] ;
  assign new_new_n1392__ = \a[12]  & \b[7] ;
  assign new_new_n1393__ = \a[13]  & \b[6] ;
  assign new_new_n1394__ = ~new_new_n1392__ & ~new_new_n1393__;
  assign new_new_n1395__ = new_new_n1392__ & new_new_n1393__;
  assign new_new_n1396__ = ~new_new_n1394__ & ~new_new_n1395__;
  assign new_new_n1397__ = ~new_new_n1391__ & ~new_new_n1396__;
  assign new_new_n1398__ = new_new_n1391__ & new_new_n1396__;
  assign new_new_n1399__ = ~new_new_n1397__ & ~new_new_n1398__;
  assign new_new_n1400__ = new_new_n1302__ & new_new_n1399__;
  assign new_new_n1401__ = ~new_new_n1302__ & ~new_new_n1399__;
  assign new_new_n1402__ = ~new_new_n1400__ & ~new_new_n1401__;
  assign new_new_n1403__ = ~new_new_n1390__ & new_new_n1402__;
  assign new_new_n1404__ = new_new_n1390__ & ~new_new_n1402__;
  assign new_new_n1405__ = ~new_new_n1403__ & ~new_new_n1404__;
  assign new_new_n1406__ = \a[15]  & \b[4] ;
  assign new_new_n1407__ = \a[14]  & \b[5] ;
  assign new_new_n1408__ = ~new_new_n1406__ & ~new_new_n1407__;
  assign new_new_n1409__ = new_new_n1406__ & new_new_n1407__;
  assign new_new_n1410__ = ~new_new_n1408__ & ~new_new_n1409__;
  assign new_new_n1411__ = new_new_n1304__ & new_new_n1410__;
  assign new_new_n1412__ = ~new_new_n1304__ & ~new_new_n1410__;
  assign new_new_n1413__ = ~new_new_n1411__ & ~new_new_n1412__;
  assign new_new_n1414__ = new_new_n1405__ & new_new_n1413__;
  assign new_new_n1415__ = ~new_new_n1405__ & ~new_new_n1413__;
  assign new_new_n1416__ = ~new_new_n1414__ & ~new_new_n1415__;
  assign new_new_n1417__ = ~new_new_n1389__ & new_new_n1416__;
  assign new_new_n1418__ = new_new_n1389__ & ~new_new_n1416__;
  assign new_new_n1419__ = ~new_new_n1417__ & ~new_new_n1418__;
  assign new_new_n1420__ = ~new_new_n1336__ & ~new_new_n1340__;
  assign new_new_n1421__ = \a[5]  & \b[14] ;
  assign new_new_n1422__ = \a[6]  & \b[13] ;
  assign new_new_n1423__ = \a[7]  & \b[12] ;
  assign new_new_n1424__ = ~new_new_n1422__ & ~new_new_n1423__;
  assign new_new_n1425__ = new_new_n1422__ & new_new_n1423__;
  assign new_new_n1426__ = ~new_new_n1424__ & ~new_new_n1425__;
  assign new_new_n1427__ = new_new_n1421__ & new_new_n1426__;
  assign new_new_n1428__ = ~new_new_n1421__ & ~new_new_n1426__;
  assign new_new_n1429__ = ~new_new_n1427__ & ~new_new_n1428__;
  assign new_new_n1430__ = ~new_new_n1331__ & ~new_new_n1333__;
  assign new_new_n1431__ = \a[8]  & \b[11] ;
  assign new_new_n1432__ = \a[9]  & \b[10] ;
  assign new_new_n1433__ = \a[10]  & \b[9] ;
  assign new_new_n1434__ = ~new_new_n1432__ & ~new_new_n1433__;
  assign new_new_n1435__ = new_new_n1432__ & new_new_n1433__;
  assign new_new_n1436__ = ~new_new_n1434__ & ~new_new_n1435__;
  assign new_new_n1437__ = new_new_n1431__ & new_new_n1436__;
  assign new_new_n1438__ = ~new_new_n1431__ & ~new_new_n1436__;
  assign new_new_n1439__ = ~new_new_n1437__ & ~new_new_n1438__;
  assign new_new_n1440__ = ~new_new_n1430__ & new_new_n1439__;
  assign new_new_n1441__ = new_new_n1430__ & ~new_new_n1439__;
  assign new_new_n1442__ = ~new_new_n1440__ & ~new_new_n1441__;
  assign new_new_n1443__ = ~new_new_n1429__ & ~new_new_n1442__;
  assign new_new_n1444__ = new_new_n1429__ & new_new_n1442__;
  assign new_new_n1445__ = ~new_new_n1443__ & ~new_new_n1444__;
  assign new_new_n1446__ = ~new_new_n1291__ & ~new_new_n1294__;
  assign new_new_n1447__ = new_new_n1445__ & ~new_new_n1446__;
  assign new_new_n1448__ = ~new_new_n1445__ & new_new_n1446__;
  assign new_new_n1449__ = ~new_new_n1447__ & ~new_new_n1448__;
  assign new_new_n1450__ = ~new_new_n1420__ & new_new_n1449__;
  assign new_new_n1451__ = new_new_n1420__ & ~new_new_n1449__;
  assign new_new_n1452__ = ~new_new_n1450__ & ~new_new_n1451__;
  assign new_new_n1453__ = new_new_n1419__ & new_new_n1452__;
  assign new_new_n1454__ = ~new_new_n1419__ & ~new_new_n1452__;
  assign new_new_n1455__ = ~new_new_n1453__ & ~new_new_n1454__;
  assign new_new_n1456__ = ~new_new_n1388__ & new_new_n1455__;
  assign new_new_n1457__ = new_new_n1388__ & ~new_new_n1455__;
  assign new_new_n1458__ = ~new_new_n1456__ & ~new_new_n1457__;
  assign new_new_n1459__ = new_new_n1387__ & new_new_n1458__;
  assign new_new_n1460__ = ~new_new_n1387__ & ~new_new_n1458__;
  assign new_new_n1461__ = ~new_new_n1459__ & ~new_new_n1460__;
  assign new_new_n1462__ = ~new_new_n1378__ & new_new_n1461__;
  assign new_new_n1463__ = new_new_n1378__ & ~new_new_n1461__;
  assign new_new_n1464__ = ~new_new_n1462__ & ~new_new_n1463__;
  assign new_new_n1465__ = ~new_new_n1377__ & new_new_n1464__;
  assign new_new_n1466__ = new_new_n1377__ & ~new_new_n1464__;
  assign new_new_n1467__ = ~new_new_n1465__ & ~new_new_n1466__;
  assign new_new_n1468__ = ~new_new_n1376__ & new_new_n1467__;
  assign new_new_n1469__ = new_new_n1376__ & ~new_new_n1467__;
  assign new_new_n1470__ = ~new_new_n1468__ & ~new_new_n1469__;
  assign new_new_n1471__ = new_new_n1375__ & new_new_n1470__;
  assign new_new_n1472__ = ~new_new_n1375__ & ~new_new_n1470__;
  assign \r[19]  = new_new_n1471__ | new_new_n1472__;
  assign new_new_n1474__ = new_new_n1366__ & new_new_n1470__;
  assign new_new_n1475__ = new_new_n1369__ & new_new_n1474__;
  assign new_new_n1476__ = ~new_new_n1150__ & new_new_n1475__;
  assign new_new_n1477__ = new_new_n1364__ & ~new_new_n1469__;
  assign new_new_n1478__ = new_new_n1368__ & new_new_n1474__;
  assign new_new_n1479__ = ~new_new_n1468__ & ~new_new_n1477__;
  assign new_new_n1480__ = ~new_new_n1478__ & new_new_n1479__;
  assign new_new_n1481__ = ~new_new_n1476__ & new_new_n1480__;
  assign new_new_n1482__ = ~new_new_n1462__ & ~new_new_n1465__;
  assign new_new_n1483__ = ~new_new_n1382__ & ~new_new_n1385__;
  assign new_new_n1484__ = ~new_new_n1456__ & ~new_new_n1459__;
  assign new_new_n1485__ = \a[5]  & \b[15] ;
  assign new_new_n1486__ = ~new_new_n1425__ & ~new_new_n1427__;
  assign new_new_n1487__ = ~new_new_n1447__ & ~new_new_n1450__;
  assign new_new_n1488__ = ~new_new_n1486__ & ~new_new_n1487__;
  assign new_new_n1489__ = new_new_n1486__ & new_new_n1487__;
  assign new_new_n1490__ = ~new_new_n1488__ & ~new_new_n1489__;
  assign new_new_n1491__ = new_new_n1485__ & new_new_n1490__;
  assign new_new_n1492__ = ~new_new_n1485__ & ~new_new_n1490__;
  assign new_new_n1493__ = ~new_new_n1491__ & ~new_new_n1492__;
  assign new_new_n1494__ = ~new_new_n1417__ & ~new_new_n1453__;
  assign new_new_n1495__ = ~new_new_n1440__ & ~new_new_n1444__;
  assign new_new_n1496__ = \a[6]  & \b[14] ;
  assign new_new_n1497__ = \a[7]  & \b[13] ;
  assign new_new_n1498__ = \a[8]  & \b[12] ;
  assign new_new_n1499__ = ~new_new_n1497__ & ~new_new_n1498__;
  assign new_new_n1500__ = new_new_n1497__ & new_new_n1498__;
  assign new_new_n1501__ = ~new_new_n1499__ & ~new_new_n1500__;
  assign new_new_n1502__ = new_new_n1496__ & new_new_n1501__;
  assign new_new_n1503__ = ~new_new_n1496__ & ~new_new_n1501__;
  assign new_new_n1504__ = ~new_new_n1502__ & ~new_new_n1503__;
  assign new_new_n1505__ = ~new_new_n1435__ & ~new_new_n1437__;
  assign new_new_n1506__ = \a[9]  & \b[11] ;
  assign new_new_n1507__ = \a[10]  & \b[10] ;
  assign new_new_n1508__ = \a[11]  & \b[9] ;
  assign new_new_n1509__ = ~new_new_n1507__ & ~new_new_n1508__;
  assign new_new_n1510__ = new_new_n1507__ & new_new_n1508__;
  assign new_new_n1511__ = ~new_new_n1509__ & ~new_new_n1510__;
  assign new_new_n1512__ = new_new_n1506__ & new_new_n1511__;
  assign new_new_n1513__ = ~new_new_n1506__ & ~new_new_n1511__;
  assign new_new_n1514__ = ~new_new_n1512__ & ~new_new_n1513__;
  assign new_new_n1515__ = ~new_new_n1505__ & new_new_n1514__;
  assign new_new_n1516__ = new_new_n1505__ & ~new_new_n1514__;
  assign new_new_n1517__ = ~new_new_n1515__ & ~new_new_n1516__;
  assign new_new_n1518__ = ~new_new_n1504__ & ~new_new_n1517__;
  assign new_new_n1519__ = new_new_n1504__ & new_new_n1517__;
  assign new_new_n1520__ = ~new_new_n1518__ & ~new_new_n1519__;
  assign new_new_n1521__ = ~new_new_n1400__ & ~new_new_n1403__;
  assign new_new_n1522__ = new_new_n1520__ & ~new_new_n1521__;
  assign new_new_n1523__ = ~new_new_n1520__ & new_new_n1521__;
  assign new_new_n1524__ = ~new_new_n1522__ & ~new_new_n1523__;
  assign new_new_n1525__ = ~new_new_n1495__ & new_new_n1524__;
  assign new_new_n1526__ = new_new_n1495__ & ~new_new_n1524__;
  assign new_new_n1527__ = ~new_new_n1525__ & ~new_new_n1526__;
  assign new_new_n1528__ = ~new_new_n1411__ & ~new_new_n1414__;
  assign new_new_n1529__ = \a[15]  & \b[5] ;
  assign new_new_n1530__ = ~new_new_n1395__ & ~new_new_n1398__;
  assign new_new_n1531__ = \a[12]  & \b[8] ;
  assign new_new_n1532__ = \a[13]  & \b[7] ;
  assign new_new_n1533__ = \a[14]  & \b[6] ;
  assign new_new_n1534__ = ~new_new_n1532__ & ~new_new_n1533__;
  assign new_new_n1535__ = new_new_n1532__ & new_new_n1533__;
  assign new_new_n1536__ = ~new_new_n1534__ & ~new_new_n1535__;
  assign new_new_n1537__ = new_new_n1531__ & new_new_n1536__;
  assign new_new_n1538__ = ~new_new_n1531__ & ~new_new_n1536__;
  assign new_new_n1539__ = ~new_new_n1537__ & ~new_new_n1538__;
  assign new_new_n1540__ = new_new_n1409__ & new_new_n1539__;
  assign new_new_n1541__ = ~new_new_n1409__ & ~new_new_n1539__;
  assign new_new_n1542__ = ~new_new_n1540__ & ~new_new_n1541__;
  assign new_new_n1543__ = new_new_n1530__ & ~new_new_n1542__;
  assign new_new_n1544__ = ~new_new_n1530__ & new_new_n1542__;
  assign new_new_n1545__ = ~new_new_n1543__ & ~new_new_n1544__;
  assign new_new_n1546__ = new_new_n1529__ & new_new_n1545__;
  assign new_new_n1547__ = ~new_new_n1529__ & ~new_new_n1545__;
  assign new_new_n1548__ = ~new_new_n1546__ & ~new_new_n1547__;
  assign new_new_n1549__ = ~new_new_n1528__ & new_new_n1548__;
  assign new_new_n1550__ = new_new_n1528__ & ~new_new_n1548__;
  assign new_new_n1551__ = ~new_new_n1549__ & ~new_new_n1550__;
  assign new_new_n1552__ = new_new_n1527__ & new_new_n1551__;
  assign new_new_n1553__ = ~new_new_n1527__ & ~new_new_n1551__;
  assign new_new_n1554__ = ~new_new_n1552__ & ~new_new_n1553__;
  assign new_new_n1555__ = ~new_new_n1494__ & new_new_n1554__;
  assign new_new_n1556__ = new_new_n1494__ & ~new_new_n1554__;
  assign new_new_n1557__ = ~new_new_n1555__ & ~new_new_n1556__;
  assign new_new_n1558__ = new_new_n1493__ & new_new_n1557__;
  assign new_new_n1559__ = ~new_new_n1493__ & ~new_new_n1557__;
  assign new_new_n1560__ = ~new_new_n1558__ & ~new_new_n1559__;
  assign new_new_n1561__ = ~new_new_n1484__ & new_new_n1560__;
  assign new_new_n1562__ = new_new_n1484__ & ~new_new_n1560__;
  assign new_new_n1563__ = ~new_new_n1561__ & ~new_new_n1562__;
  assign new_new_n1564__ = ~new_new_n1483__ & new_new_n1563__;
  assign new_new_n1565__ = new_new_n1483__ & ~new_new_n1563__;
  assign new_new_n1566__ = ~new_new_n1564__ & ~new_new_n1565__;
  assign new_new_n1567__ = ~new_new_n1482__ & new_new_n1566__;
  assign new_new_n1568__ = new_new_n1482__ & ~new_new_n1566__;
  assign new_new_n1569__ = ~new_new_n1567__ & ~new_new_n1568__;
  assign new_new_n1570__ = ~new_new_n1481__ & new_new_n1569__;
  assign new_new_n1571__ = new_new_n1481__ & ~new_new_n1569__;
  assign \r[20]  = ~new_new_n1570__ & ~new_new_n1571__;
  assign new_new_n1573__ = ~new_new_n1567__ & ~new_new_n1570__;
  assign new_new_n1574__ = ~new_new_n1561__ & ~new_new_n1564__;
  assign new_new_n1575__ = ~new_new_n1488__ & ~new_new_n1491__;
  assign new_new_n1576__ = ~new_new_n1555__ & ~new_new_n1558__;
  assign new_new_n1577__ = \a[6]  & \b[15] ;
  assign new_new_n1578__ = ~new_new_n1500__ & ~new_new_n1502__;
  assign new_new_n1579__ = ~new_new_n1522__ & ~new_new_n1525__;
  assign new_new_n1580__ = ~new_new_n1578__ & ~new_new_n1579__;
  assign new_new_n1581__ = new_new_n1578__ & new_new_n1579__;
  assign new_new_n1582__ = ~new_new_n1580__ & ~new_new_n1581__;
  assign new_new_n1583__ = new_new_n1577__ & new_new_n1582__;
  assign new_new_n1584__ = ~new_new_n1577__ & ~new_new_n1582__;
  assign new_new_n1585__ = ~new_new_n1583__ & ~new_new_n1584__;
  assign new_new_n1586__ = ~new_new_n1549__ & ~new_new_n1552__;
  assign new_new_n1587__ = ~new_new_n1515__ & ~new_new_n1519__;
  assign new_new_n1588__ = \a[7]  & \b[14] ;
  assign new_new_n1589__ = \a[8]  & \b[13] ;
  assign new_new_n1590__ = \a[9]  & \b[12] ;
  assign new_new_n1591__ = ~new_new_n1589__ & ~new_new_n1590__;
  assign new_new_n1592__ = new_new_n1589__ & new_new_n1590__;
  assign new_new_n1593__ = ~new_new_n1591__ & ~new_new_n1592__;
  assign new_new_n1594__ = new_new_n1588__ & new_new_n1593__;
  assign new_new_n1595__ = ~new_new_n1588__ & ~new_new_n1593__;
  assign new_new_n1596__ = ~new_new_n1594__ & ~new_new_n1595__;
  assign new_new_n1597__ = ~new_new_n1510__ & ~new_new_n1512__;
  assign new_new_n1598__ = \a[10]  & \b[11] ;
  assign new_new_n1599__ = \a[11]  & \b[10] ;
  assign new_new_n1600__ = \a[12]  & \b[9] ;
  assign new_new_n1601__ = ~new_new_n1599__ & ~new_new_n1600__;
  assign new_new_n1602__ = new_new_n1599__ & new_new_n1600__;
  assign new_new_n1603__ = ~new_new_n1601__ & ~new_new_n1602__;
  assign new_new_n1604__ = new_new_n1598__ & new_new_n1603__;
  assign new_new_n1605__ = ~new_new_n1598__ & ~new_new_n1603__;
  assign new_new_n1606__ = ~new_new_n1604__ & ~new_new_n1605__;
  assign new_new_n1607__ = ~new_new_n1597__ & new_new_n1606__;
  assign new_new_n1608__ = new_new_n1597__ & ~new_new_n1606__;
  assign new_new_n1609__ = ~new_new_n1607__ & ~new_new_n1608__;
  assign new_new_n1610__ = ~new_new_n1596__ & ~new_new_n1609__;
  assign new_new_n1611__ = new_new_n1596__ & new_new_n1609__;
  assign new_new_n1612__ = ~new_new_n1610__ & ~new_new_n1611__;
  assign new_new_n1613__ = ~new_new_n1540__ & ~new_new_n1544__;
  assign new_new_n1614__ = new_new_n1612__ & ~new_new_n1613__;
  assign new_new_n1615__ = ~new_new_n1612__ & new_new_n1613__;
  assign new_new_n1616__ = ~new_new_n1614__ & ~new_new_n1615__;
  assign new_new_n1617__ = ~new_new_n1587__ & new_new_n1616__;
  assign new_new_n1618__ = new_new_n1587__ & ~new_new_n1616__;
  assign new_new_n1619__ = ~new_new_n1617__ & ~new_new_n1618__;
  assign new_new_n1620__ = ~new_new_n1535__ & ~new_new_n1537__;
  assign new_new_n1621__ = \a[13]  & \b[8] ;
  assign new_new_n1622__ = \a[14]  & \b[7] ;
  assign new_new_n1623__ = \a[15]  & \b[6] ;
  assign new_new_n1624__ = ~new_new_n1622__ & ~new_new_n1623__;
  assign new_new_n1625__ = new_new_n1622__ & new_new_n1623__;
  assign new_new_n1626__ = ~new_new_n1624__ & ~new_new_n1625__;
  assign new_new_n1627__ = new_new_n1621__ & new_new_n1626__;
  assign new_new_n1628__ = ~new_new_n1621__ & ~new_new_n1626__;
  assign new_new_n1629__ = ~new_new_n1627__ & ~new_new_n1628__;
  assign new_new_n1630__ = ~new_new_n1620__ & new_new_n1629__;
  assign new_new_n1631__ = new_new_n1620__ & ~new_new_n1629__;
  assign new_new_n1632__ = ~new_new_n1630__ & ~new_new_n1631__;
  assign new_new_n1633__ = new_new_n1546__ & new_new_n1632__;
  assign new_new_n1634__ = ~new_new_n1546__ & ~new_new_n1632__;
  assign new_new_n1635__ = ~new_new_n1633__ & ~new_new_n1634__;
  assign new_new_n1636__ = new_new_n1619__ & new_new_n1635__;
  assign new_new_n1637__ = ~new_new_n1619__ & ~new_new_n1635__;
  assign new_new_n1638__ = ~new_new_n1636__ & ~new_new_n1637__;
  assign new_new_n1639__ = ~new_new_n1586__ & new_new_n1638__;
  assign new_new_n1640__ = new_new_n1586__ & ~new_new_n1638__;
  assign new_new_n1641__ = ~new_new_n1639__ & ~new_new_n1640__;
  assign new_new_n1642__ = new_new_n1585__ & new_new_n1641__;
  assign new_new_n1643__ = ~new_new_n1585__ & ~new_new_n1641__;
  assign new_new_n1644__ = ~new_new_n1642__ & ~new_new_n1643__;
  assign new_new_n1645__ = ~new_new_n1576__ & new_new_n1644__;
  assign new_new_n1646__ = new_new_n1576__ & ~new_new_n1644__;
  assign new_new_n1647__ = ~new_new_n1645__ & ~new_new_n1646__;
  assign new_new_n1648__ = ~new_new_n1575__ & new_new_n1647__;
  assign new_new_n1649__ = new_new_n1575__ & ~new_new_n1647__;
  assign new_new_n1650__ = ~new_new_n1648__ & ~new_new_n1649__;
  assign new_new_n1651__ = ~new_new_n1574__ & new_new_n1650__;
  assign new_new_n1652__ = new_new_n1574__ & ~new_new_n1650__;
  assign new_new_n1653__ = ~new_new_n1651__ & ~new_new_n1652__;
  assign new_new_n1654__ = new_new_n1573__ & new_new_n1653__;
  assign new_new_n1655__ = ~new_new_n1573__ & ~new_new_n1653__;
  assign \r[21]  = new_new_n1654__ | new_new_n1655__;
  assign new_new_n1657__ = ~new_new_n1645__ & ~new_new_n1648__;
  assign new_new_n1658__ = ~new_new_n1580__ & ~new_new_n1583__;
  assign new_new_n1659__ = ~new_new_n1639__ & ~new_new_n1642__;
  assign new_new_n1660__ = \a[7]  & \b[15] ;
  assign new_new_n1661__ = ~new_new_n1592__ & ~new_new_n1594__;
  assign new_new_n1662__ = ~new_new_n1614__ & ~new_new_n1617__;
  assign new_new_n1663__ = ~new_new_n1661__ & ~new_new_n1662__;
  assign new_new_n1664__ = new_new_n1661__ & new_new_n1662__;
  assign new_new_n1665__ = ~new_new_n1663__ & ~new_new_n1664__;
  assign new_new_n1666__ = new_new_n1660__ & new_new_n1665__;
  assign new_new_n1667__ = ~new_new_n1660__ & ~new_new_n1665__;
  assign new_new_n1668__ = ~new_new_n1666__ & ~new_new_n1667__;
  assign new_new_n1669__ = ~new_new_n1633__ & ~new_new_n1636__;
  assign new_new_n1670__ = ~new_new_n1607__ & ~new_new_n1611__;
  assign new_new_n1671__ = \a[8]  & \b[14] ;
  assign new_new_n1672__ = \a[9]  & \b[13] ;
  assign new_new_n1673__ = \a[10]  & \b[12] ;
  assign new_new_n1674__ = ~new_new_n1672__ & ~new_new_n1673__;
  assign new_new_n1675__ = new_new_n1672__ & new_new_n1673__;
  assign new_new_n1676__ = ~new_new_n1674__ & ~new_new_n1675__;
  assign new_new_n1677__ = new_new_n1671__ & new_new_n1676__;
  assign new_new_n1678__ = ~new_new_n1671__ & ~new_new_n1676__;
  assign new_new_n1679__ = ~new_new_n1677__ & ~new_new_n1678__;
  assign new_new_n1680__ = ~new_new_n1602__ & ~new_new_n1604__;
  assign new_new_n1681__ = \a[11]  & \b[11] ;
  assign new_new_n1682__ = \a[12]  & \b[10] ;
  assign new_new_n1683__ = \a[13]  & \b[9] ;
  assign new_new_n1684__ = ~new_new_n1682__ & ~new_new_n1683__;
  assign new_new_n1685__ = new_new_n1682__ & new_new_n1683__;
  assign new_new_n1686__ = ~new_new_n1684__ & ~new_new_n1685__;
  assign new_new_n1687__ = new_new_n1681__ & new_new_n1686__;
  assign new_new_n1688__ = ~new_new_n1681__ & ~new_new_n1686__;
  assign new_new_n1689__ = ~new_new_n1687__ & ~new_new_n1688__;
  assign new_new_n1690__ = ~new_new_n1680__ & new_new_n1689__;
  assign new_new_n1691__ = new_new_n1680__ & ~new_new_n1689__;
  assign new_new_n1692__ = ~new_new_n1690__ & ~new_new_n1691__;
  assign new_new_n1693__ = ~new_new_n1679__ & ~new_new_n1692__;
  assign new_new_n1694__ = new_new_n1679__ & new_new_n1692__;
  assign new_new_n1695__ = ~new_new_n1693__ & ~new_new_n1694__;
  assign new_new_n1696__ = new_new_n1630__ & new_new_n1695__;
  assign new_new_n1697__ = ~new_new_n1630__ & ~new_new_n1695__;
  assign new_new_n1698__ = ~new_new_n1696__ & ~new_new_n1697__;
  assign new_new_n1699__ = new_new_n1670__ & ~new_new_n1698__;
  assign new_new_n1700__ = ~new_new_n1670__ & new_new_n1698__;
  assign new_new_n1701__ = ~new_new_n1699__ & ~new_new_n1700__;
  assign new_new_n1702__ = ~new_new_n1625__ & ~new_new_n1627__;
  assign new_new_n1703__ = \a[15]  & \b[7] ;
  assign new_new_n1704__ = \a[14]  & \b[8] ;
  assign new_new_n1705__ = ~new_new_n1703__ & ~new_new_n1704__;
  assign new_new_n1706__ = new_new_n1703__ & new_new_n1704__;
  assign new_new_n1707__ = ~new_new_n1705__ & ~new_new_n1706__;
  assign new_new_n1708__ = new_new_n1702__ & ~new_new_n1707__;
  assign new_new_n1709__ = ~new_new_n1702__ & new_new_n1707__;
  assign new_new_n1710__ = ~new_new_n1708__ & ~new_new_n1709__;
  assign new_new_n1711__ = new_new_n1701__ & new_new_n1710__;
  assign new_new_n1712__ = ~new_new_n1701__ & ~new_new_n1710__;
  assign new_new_n1713__ = ~new_new_n1711__ & ~new_new_n1712__;
  assign new_new_n1714__ = ~new_new_n1669__ & new_new_n1713__;
  assign new_new_n1715__ = new_new_n1669__ & ~new_new_n1713__;
  assign new_new_n1716__ = ~new_new_n1714__ & ~new_new_n1715__;
  assign new_new_n1717__ = new_new_n1668__ & new_new_n1716__;
  assign new_new_n1718__ = ~new_new_n1668__ & ~new_new_n1716__;
  assign new_new_n1719__ = ~new_new_n1717__ & ~new_new_n1718__;
  assign new_new_n1720__ = ~new_new_n1659__ & new_new_n1719__;
  assign new_new_n1721__ = new_new_n1659__ & ~new_new_n1719__;
  assign new_new_n1722__ = ~new_new_n1720__ & ~new_new_n1721__;
  assign new_new_n1723__ = ~new_new_n1658__ & new_new_n1722__;
  assign new_new_n1724__ = new_new_n1658__ & ~new_new_n1722__;
  assign new_new_n1725__ = ~new_new_n1723__ & ~new_new_n1724__;
  assign new_new_n1726__ = ~new_new_n1657__ & new_new_n1725__;
  assign new_new_n1727__ = new_new_n1657__ & ~new_new_n1725__;
  assign new_new_n1728__ = ~new_new_n1726__ & ~new_new_n1727__;
  assign new_new_n1729__ = new_new_n1573__ & ~new_new_n1651__;
  assign new_new_n1730__ = ~new_new_n1652__ & ~new_new_n1729__;
  assign new_new_n1731__ = new_new_n1728__ & new_new_n1730__;
  assign new_new_n1732__ = ~new_new_n1728__ & ~new_new_n1730__;
  assign \r[22]  = ~new_new_n1731__ & ~new_new_n1732__;
  assign new_new_n1734__ = ~new_new_n1726__ & ~new_new_n1731__;
  assign new_new_n1735__ = ~new_new_n1720__ & ~new_new_n1723__;
  assign new_new_n1736__ = ~new_new_n1663__ & ~new_new_n1666__;
  assign new_new_n1737__ = ~new_new_n1714__ & ~new_new_n1717__;
  assign new_new_n1738__ = \a[8]  & \b[15] ;
  assign new_new_n1739__ = ~new_new_n1675__ & ~new_new_n1677__;
  assign new_new_n1740__ = ~new_new_n1696__ & ~new_new_n1700__;
  assign new_new_n1741__ = ~new_new_n1739__ & ~new_new_n1740__;
  assign new_new_n1742__ = new_new_n1739__ & new_new_n1740__;
  assign new_new_n1743__ = ~new_new_n1741__ & ~new_new_n1742__;
  assign new_new_n1744__ = new_new_n1738__ & new_new_n1743__;
  assign new_new_n1745__ = ~new_new_n1738__ & ~new_new_n1743__;
  assign new_new_n1746__ = ~new_new_n1744__ & ~new_new_n1745__;
  assign new_new_n1747__ = ~new_new_n1690__ & ~new_new_n1694__;
  assign new_new_n1748__ = \a[9]  & \b[14] ;
  assign new_new_n1749__ = \a[10]  & \b[13] ;
  assign new_new_n1750__ = \a[11]  & \b[12] ;
  assign new_new_n1751__ = ~new_new_n1749__ & ~new_new_n1750__;
  assign new_new_n1752__ = new_new_n1749__ & new_new_n1750__;
  assign new_new_n1753__ = ~new_new_n1751__ & ~new_new_n1752__;
  assign new_new_n1754__ = new_new_n1748__ & new_new_n1753__;
  assign new_new_n1755__ = ~new_new_n1748__ & ~new_new_n1753__;
  assign new_new_n1756__ = ~new_new_n1754__ & ~new_new_n1755__;
  assign new_new_n1757__ = ~new_new_n1685__ & ~new_new_n1687__;
  assign new_new_n1758__ = \a[12]  & \b[11] ;
  assign new_new_n1759__ = \a[13]  & \b[10] ;
  assign new_new_n1760__ = \a[14]  & \b[9] ;
  assign new_new_n1761__ = ~new_new_n1759__ & ~new_new_n1760__;
  assign new_new_n1762__ = new_new_n1759__ & new_new_n1760__;
  assign new_new_n1763__ = ~new_new_n1761__ & ~new_new_n1762__;
  assign new_new_n1764__ = new_new_n1758__ & new_new_n1763__;
  assign new_new_n1765__ = ~new_new_n1758__ & ~new_new_n1763__;
  assign new_new_n1766__ = ~new_new_n1764__ & ~new_new_n1765__;
  assign new_new_n1767__ = ~new_new_n1757__ & new_new_n1766__;
  assign new_new_n1768__ = new_new_n1757__ & ~new_new_n1766__;
  assign new_new_n1769__ = ~new_new_n1767__ & ~new_new_n1768__;
  assign new_new_n1770__ = ~new_new_n1756__ & ~new_new_n1769__;
  assign new_new_n1771__ = new_new_n1756__ & new_new_n1769__;
  assign new_new_n1772__ = ~new_new_n1770__ & ~new_new_n1771__;
  assign new_new_n1773__ = new_new_n1709__ & new_new_n1772__;
  assign new_new_n1774__ = ~new_new_n1709__ & ~new_new_n1772__;
  assign new_new_n1775__ = ~new_new_n1773__ & ~new_new_n1774__;
  assign new_new_n1776__ = new_new_n1747__ & ~new_new_n1775__;
  assign new_new_n1777__ = ~new_new_n1747__ & new_new_n1775__;
  assign new_new_n1778__ = ~new_new_n1776__ & ~new_new_n1777__;
  assign new_new_n1779__ = \a[15]  & \b[8] ;
  assign new_new_n1780__ = ~new_new_n1622__ & new_new_n1779__;
  assign new_new_n1781__ = new_new_n1778__ & new_new_n1780__;
  assign new_new_n1782__ = ~new_new_n1778__ & ~new_new_n1780__;
  assign new_new_n1783__ = ~new_new_n1781__ & ~new_new_n1782__;
  assign new_new_n1784__ = new_new_n1711__ & new_new_n1783__;
  assign new_new_n1785__ = ~new_new_n1711__ & ~new_new_n1783__;
  assign new_new_n1786__ = ~new_new_n1784__ & ~new_new_n1785__;
  assign new_new_n1787__ = new_new_n1746__ & new_new_n1786__;
  assign new_new_n1788__ = ~new_new_n1746__ & ~new_new_n1786__;
  assign new_new_n1789__ = ~new_new_n1787__ & ~new_new_n1788__;
  assign new_new_n1790__ = ~new_new_n1737__ & new_new_n1789__;
  assign new_new_n1791__ = new_new_n1737__ & ~new_new_n1789__;
  assign new_new_n1792__ = ~new_new_n1790__ & ~new_new_n1791__;
  assign new_new_n1793__ = ~new_new_n1736__ & new_new_n1792__;
  assign new_new_n1794__ = new_new_n1736__ & ~new_new_n1792__;
  assign new_new_n1795__ = ~new_new_n1793__ & ~new_new_n1794__;
  assign new_new_n1796__ = ~new_new_n1735__ & new_new_n1795__;
  assign new_new_n1797__ = new_new_n1735__ & ~new_new_n1795__;
  assign new_new_n1798__ = ~new_new_n1796__ & ~new_new_n1797__;
  assign new_new_n1799__ = new_new_n1734__ & new_new_n1798__;
  assign new_new_n1800__ = ~new_new_n1734__ & ~new_new_n1798__;
  assign \r[23]  = new_new_n1799__ | new_new_n1800__;
  assign new_new_n1802__ = new_new_n1728__ & new_new_n1798__;
  assign new_new_n1803__ = new_new_n1569__ & new_new_n1802__;
  assign new_new_n1804__ = new_new_n1653__ & new_new_n1803__;
  assign new_new_n1805__ = new_new_n1476__ & new_new_n1804__;
  assign new_new_n1806__ = ~new_new_n1480__ & new_new_n1804__;
  assign new_new_n1807__ = new_new_n1726__ & ~new_new_n1797__;
  assign new_new_n1808__ = ~new_new_n1567__ & ~new_new_n1651__;
  assign new_new_n1809__ = ~new_new_n1652__ & new_new_n1802__;
  assign new_new_n1810__ = ~new_new_n1808__ & new_new_n1809__;
  assign new_new_n1811__ = ~new_new_n1796__ & ~new_new_n1807__;
  assign new_new_n1812__ = ~new_new_n1810__ & new_new_n1811__;
  assign new_new_n1813__ = ~new_new_n1806__ & new_new_n1812__;
  assign new_new_n1814__ = ~new_new_n1805__ & new_new_n1813__;
  assign new_new_n1815__ = ~new_new_n1790__ & ~new_new_n1793__;
  assign new_new_n1816__ = ~new_new_n1741__ & ~new_new_n1744__;
  assign new_new_n1817__ = ~new_new_n1784__ & ~new_new_n1787__;
  assign new_new_n1818__ = \a[9]  & \b[15] ;
  assign new_new_n1819__ = ~new_new_n1752__ & ~new_new_n1754__;
  assign new_new_n1820__ = ~new_new_n1773__ & ~new_new_n1777__;
  assign new_new_n1821__ = ~new_new_n1819__ & ~new_new_n1820__;
  assign new_new_n1822__ = new_new_n1819__ & new_new_n1820__;
  assign new_new_n1823__ = ~new_new_n1821__ & ~new_new_n1822__;
  assign new_new_n1824__ = new_new_n1818__ & new_new_n1823__;
  assign new_new_n1825__ = ~new_new_n1818__ & ~new_new_n1823__;
  assign new_new_n1826__ = ~new_new_n1824__ & ~new_new_n1825__;
  assign new_new_n1827__ = ~new_new_n1767__ & ~new_new_n1771__;
  assign new_new_n1828__ = \a[10]  & \b[14] ;
  assign new_new_n1829__ = \a[11]  & \b[13] ;
  assign new_new_n1830__ = \a[12]  & \b[12] ;
  assign new_new_n1831__ = ~new_new_n1829__ & ~new_new_n1830__;
  assign new_new_n1832__ = new_new_n1829__ & new_new_n1830__;
  assign new_new_n1833__ = ~new_new_n1831__ & ~new_new_n1832__;
  assign new_new_n1834__ = new_new_n1828__ & new_new_n1833__;
  assign new_new_n1835__ = ~new_new_n1828__ & ~new_new_n1833__;
  assign new_new_n1836__ = ~new_new_n1834__ & ~new_new_n1835__;
  assign new_new_n1837__ = ~new_new_n1762__ & ~new_new_n1764__;
  assign new_new_n1838__ = \a[13]  & \b[11] ;
  assign new_new_n1839__ = \a[14]  & \b[10] ;
  assign new_new_n1840__ = \a[15]  & \b[9] ;
  assign new_new_n1841__ = ~new_new_n1839__ & ~new_new_n1840__;
  assign new_new_n1842__ = new_new_n1839__ & new_new_n1840__;
  assign new_new_n1843__ = ~new_new_n1841__ & ~new_new_n1842__;
  assign new_new_n1844__ = new_new_n1838__ & new_new_n1843__;
  assign new_new_n1845__ = ~new_new_n1838__ & ~new_new_n1843__;
  assign new_new_n1846__ = ~new_new_n1844__ & ~new_new_n1845__;
  assign new_new_n1847__ = ~new_new_n1837__ & new_new_n1846__;
  assign new_new_n1848__ = new_new_n1837__ & ~new_new_n1846__;
  assign new_new_n1849__ = ~new_new_n1847__ & ~new_new_n1848__;
  assign new_new_n1850__ = ~new_new_n1836__ & ~new_new_n1849__;
  assign new_new_n1851__ = new_new_n1836__ & new_new_n1849__;
  assign new_new_n1852__ = ~new_new_n1850__ & ~new_new_n1851__;
  assign new_new_n1853__ = ~new_new_n1706__ & ~new_new_n1852__;
  assign new_new_n1854__ = new_new_n1706__ & new_new_n1852__;
  assign new_new_n1855__ = ~new_new_n1853__ & ~new_new_n1854__;
  assign new_new_n1856__ = new_new_n1827__ & ~new_new_n1855__;
  assign new_new_n1857__ = ~new_new_n1827__ & new_new_n1855__;
  assign new_new_n1858__ = ~new_new_n1856__ & ~new_new_n1857__;
  assign new_new_n1859__ = new_new_n1781__ & new_new_n1858__;
  assign new_new_n1860__ = ~new_new_n1781__ & ~new_new_n1858__;
  assign new_new_n1861__ = ~new_new_n1859__ & ~new_new_n1860__;
  assign new_new_n1862__ = new_new_n1826__ & new_new_n1861__;
  assign new_new_n1863__ = ~new_new_n1826__ & ~new_new_n1861__;
  assign new_new_n1864__ = ~new_new_n1862__ & ~new_new_n1863__;
  assign new_new_n1865__ = ~new_new_n1817__ & new_new_n1864__;
  assign new_new_n1866__ = new_new_n1817__ & ~new_new_n1864__;
  assign new_new_n1867__ = ~new_new_n1865__ & ~new_new_n1866__;
  assign new_new_n1868__ = ~new_new_n1816__ & new_new_n1867__;
  assign new_new_n1869__ = new_new_n1816__ & ~new_new_n1867__;
  assign new_new_n1870__ = ~new_new_n1868__ & ~new_new_n1869__;
  assign new_new_n1871__ = ~new_new_n1815__ & new_new_n1870__;
  assign new_new_n1872__ = new_new_n1815__ & ~new_new_n1870__;
  assign new_new_n1873__ = ~new_new_n1871__ & ~new_new_n1872__;
  assign new_new_n1874__ = ~new_new_n1814__ & new_new_n1873__;
  assign new_new_n1875__ = new_new_n1814__ & ~new_new_n1873__;
  assign \r[24]  = ~new_new_n1874__ & ~new_new_n1875__;
  assign new_new_n1877__ = ~new_new_n1871__ & ~new_new_n1874__;
  assign new_new_n1878__ = ~new_new_n1865__ & ~new_new_n1868__;
  assign new_new_n1879__ = ~new_new_n1821__ & ~new_new_n1824__;
  assign new_new_n1880__ = ~new_new_n1859__ & ~new_new_n1862__;
  assign new_new_n1881__ = \a[10]  & \b[15] ;
  assign new_new_n1882__ = ~new_new_n1832__ & ~new_new_n1834__;
  assign new_new_n1883__ = ~new_new_n1854__ & ~new_new_n1857__;
  assign new_new_n1884__ = new_new_n1882__ & new_new_n1883__;
  assign new_new_n1885__ = ~new_new_n1882__ & ~new_new_n1883__;
  assign new_new_n1886__ = ~new_new_n1884__ & ~new_new_n1885__;
  assign new_new_n1887__ = new_new_n1881__ & new_new_n1886__;
  assign new_new_n1888__ = ~new_new_n1881__ & ~new_new_n1886__;
  assign new_new_n1889__ = ~new_new_n1887__ & ~new_new_n1888__;
  assign new_new_n1890__ = ~new_new_n1847__ & ~new_new_n1851__;
  assign new_new_n1891__ = \a[11]  & \b[14] ;
  assign new_new_n1892__ = \a[12]  & \b[13] ;
  assign new_new_n1893__ = \a[13]  & \b[12] ;
  assign new_new_n1894__ = ~new_new_n1892__ & ~new_new_n1893__;
  assign new_new_n1895__ = new_new_n1892__ & new_new_n1893__;
  assign new_new_n1896__ = ~new_new_n1894__ & ~new_new_n1895__;
  assign new_new_n1897__ = new_new_n1891__ & new_new_n1896__;
  assign new_new_n1898__ = ~new_new_n1891__ & ~new_new_n1896__;
  assign new_new_n1899__ = ~new_new_n1897__ & ~new_new_n1898__;
  assign new_new_n1900__ = ~new_new_n1842__ & ~new_new_n1844__;
  assign new_new_n1901__ = \a[15]  & \b[10] ;
  assign new_new_n1902__ = \a[14]  & \b[11] ;
  assign new_new_n1903__ = ~new_new_n1901__ & ~new_new_n1902__;
  assign new_new_n1904__ = new_new_n1901__ & new_new_n1902__;
  assign new_new_n1905__ = ~new_new_n1903__ & ~new_new_n1904__;
  assign new_new_n1906__ = ~new_new_n1900__ & new_new_n1905__;
  assign new_new_n1907__ = new_new_n1900__ & ~new_new_n1905__;
  assign new_new_n1908__ = ~new_new_n1906__ & ~new_new_n1907__;
  assign new_new_n1909__ = new_new_n1899__ & new_new_n1908__;
  assign new_new_n1910__ = ~new_new_n1899__ & ~new_new_n1908__;
  assign new_new_n1911__ = ~new_new_n1909__ & ~new_new_n1910__;
  assign new_new_n1912__ = new_new_n1890__ & ~new_new_n1911__;
  assign new_new_n1913__ = ~new_new_n1890__ & new_new_n1911__;
  assign new_new_n1914__ = ~new_new_n1912__ & ~new_new_n1913__;
  assign new_new_n1915__ = new_new_n1889__ & new_new_n1914__;
  assign new_new_n1916__ = ~new_new_n1889__ & ~new_new_n1914__;
  assign new_new_n1917__ = ~new_new_n1915__ & ~new_new_n1916__;
  assign new_new_n1918__ = ~new_new_n1880__ & new_new_n1917__;
  assign new_new_n1919__ = new_new_n1880__ & ~new_new_n1917__;
  assign new_new_n1920__ = ~new_new_n1918__ & ~new_new_n1919__;
  assign new_new_n1921__ = ~new_new_n1879__ & new_new_n1920__;
  assign new_new_n1922__ = new_new_n1879__ & ~new_new_n1920__;
  assign new_new_n1923__ = ~new_new_n1921__ & ~new_new_n1922__;
  assign new_new_n1924__ = new_new_n1878__ & ~new_new_n1923__;
  assign new_new_n1925__ = ~new_new_n1878__ & new_new_n1923__;
  assign new_new_n1926__ = ~new_new_n1924__ & ~new_new_n1925__;
  assign new_new_n1927__ = new_new_n1877__ & new_new_n1926__;
  assign new_new_n1928__ = ~new_new_n1877__ & ~new_new_n1926__;
  assign \r[25]  = new_new_n1927__ | new_new_n1928__;
  assign new_new_n1930__ = ~new_new_n1918__ & ~new_new_n1921__;
  assign new_new_n1931__ = ~new_new_n1885__ & ~new_new_n1887__;
  assign new_new_n1932__ = \a[11]  & \b[15] ;
  assign new_new_n1933__ = ~new_new_n1895__ & ~new_new_n1897__;
  assign new_new_n1934__ = ~new_new_n1913__ & new_new_n1933__;
  assign new_new_n1935__ = new_new_n1913__ & ~new_new_n1933__;
  assign new_new_n1936__ = ~new_new_n1934__ & ~new_new_n1935__;
  assign new_new_n1937__ = new_new_n1932__ & new_new_n1936__;
  assign new_new_n1938__ = ~new_new_n1932__ & ~new_new_n1936__;
  assign new_new_n1939__ = ~new_new_n1937__ & ~new_new_n1938__;
  assign new_new_n1940__ = ~new_new_n1906__ & ~new_new_n1909__;
  assign new_new_n1941__ = \a[12]  & \b[14] ;
  assign new_new_n1942__ = \a[13]  & \b[13] ;
  assign new_new_n1943__ = \a[14]  & \b[12] ;
  assign new_new_n1944__ = ~new_new_n1942__ & ~new_new_n1943__;
  assign new_new_n1945__ = new_new_n1942__ & new_new_n1943__;
  assign new_new_n1946__ = ~new_new_n1944__ & ~new_new_n1945__;
  assign new_new_n1947__ = new_new_n1941__ & new_new_n1946__;
  assign new_new_n1948__ = ~new_new_n1941__ & ~new_new_n1946__;
  assign new_new_n1949__ = ~new_new_n1947__ & ~new_new_n1948__;
  assign new_new_n1950__ = \a[15]  & \b[11] ;
  assign new_new_n1951__ = ~new_new_n1839__ & new_new_n1950__;
  assign new_new_n1952__ = ~new_new_n1949__ & ~new_new_n1951__;
  assign new_new_n1953__ = new_new_n1949__ & new_new_n1951__;
  assign new_new_n1954__ = ~new_new_n1952__ & ~new_new_n1953__;
  assign new_new_n1955__ = new_new_n1940__ & ~new_new_n1954__;
  assign new_new_n1956__ = ~new_new_n1940__ & new_new_n1954__;
  assign new_new_n1957__ = ~new_new_n1955__ & ~new_new_n1956__;
  assign new_new_n1958__ = new_new_n1939__ & new_new_n1957__;
  assign new_new_n1959__ = ~new_new_n1939__ & ~new_new_n1957__;
  assign new_new_n1960__ = ~new_new_n1958__ & ~new_new_n1959__;
  assign new_new_n1961__ = new_new_n1915__ & new_new_n1960__;
  assign new_new_n1962__ = ~new_new_n1915__ & ~new_new_n1960__;
  assign new_new_n1963__ = ~new_new_n1961__ & ~new_new_n1962__;
  assign new_new_n1964__ = ~new_new_n1931__ & new_new_n1963__;
  assign new_new_n1965__ = new_new_n1931__ & ~new_new_n1963__;
  assign new_new_n1966__ = ~new_new_n1964__ & ~new_new_n1965__;
  assign new_new_n1967__ = ~new_new_n1930__ & new_new_n1966__;
  assign new_new_n1968__ = new_new_n1930__ & ~new_new_n1966__;
  assign new_new_n1969__ = ~new_new_n1967__ & ~new_new_n1968__;
  assign new_new_n1970__ = ~new_new_n1871__ & ~new_new_n1925__;
  assign new_new_n1971__ = ~new_new_n1874__ & new_new_n1970__;
  assign new_new_n1972__ = ~new_new_n1924__ & ~new_new_n1971__;
  assign new_new_n1973__ = new_new_n1969__ & new_new_n1972__;
  assign new_new_n1974__ = ~new_new_n1969__ & ~new_new_n1972__;
  assign \r[26]  = ~new_new_n1973__ & ~new_new_n1974__;
  assign new_new_n1976__ = ~new_new_n1967__ & ~new_new_n1973__;
  assign new_new_n1977__ = ~new_new_n1961__ & ~new_new_n1964__;
  assign new_new_n1978__ = ~new_new_n1935__ & ~new_new_n1937__;
  assign new_new_n1979__ = \a[12]  & \b[15] ;
  assign new_new_n1980__ = ~new_new_n1945__ & ~new_new_n1947__;
  assign new_new_n1981__ = ~new_new_n1956__ & new_new_n1980__;
  assign new_new_n1982__ = new_new_n1956__ & ~new_new_n1980__;
  assign new_new_n1983__ = ~new_new_n1981__ & ~new_new_n1982__;
  assign new_new_n1984__ = new_new_n1979__ & new_new_n1983__;
  assign new_new_n1985__ = ~new_new_n1979__ & ~new_new_n1983__;
  assign new_new_n1986__ = ~new_new_n1984__ & ~new_new_n1985__;
  assign new_new_n1987__ = ~new_new_n1904__ & ~new_new_n1953__;
  assign new_new_n1988__ = \a[13]  & \b[14] ;
  assign new_new_n1989__ = \a[14]  & \b[13] ;
  assign new_new_n1990__ = \a[15]  & \b[12] ;
  assign new_new_n1991__ = ~new_new_n1989__ & ~new_new_n1990__;
  assign new_new_n1992__ = new_new_n1989__ & new_new_n1990__;
  assign new_new_n1993__ = ~new_new_n1991__ & ~new_new_n1992__;
  assign new_new_n1994__ = new_new_n1988__ & new_new_n1993__;
  assign new_new_n1995__ = ~new_new_n1988__ & ~new_new_n1993__;
  assign new_new_n1996__ = ~new_new_n1994__ & ~new_new_n1995__;
  assign new_new_n1997__ = new_new_n1987__ & ~new_new_n1996__;
  assign new_new_n1998__ = ~new_new_n1987__ & new_new_n1996__;
  assign new_new_n1999__ = ~new_new_n1997__ & ~new_new_n1998__;
  assign new_new_n2000__ = new_new_n1986__ & new_new_n1999__;
  assign new_new_n2001__ = ~new_new_n1986__ & ~new_new_n1999__;
  assign new_new_n2002__ = ~new_new_n2000__ & ~new_new_n2001__;
  assign new_new_n2003__ = new_new_n1958__ & new_new_n2002__;
  assign new_new_n2004__ = ~new_new_n1958__ & ~new_new_n2002__;
  assign new_new_n2005__ = ~new_new_n2003__ & ~new_new_n2004__;
  assign new_new_n2006__ = ~new_new_n1978__ & new_new_n2005__;
  assign new_new_n2007__ = new_new_n1978__ & ~new_new_n2005__;
  assign new_new_n2008__ = ~new_new_n2006__ & ~new_new_n2007__;
  assign new_new_n2009__ = new_new_n1977__ & ~new_new_n2008__;
  assign new_new_n2010__ = ~new_new_n1977__ & new_new_n2008__;
  assign new_new_n2011__ = ~new_new_n2009__ & ~new_new_n2010__;
  assign new_new_n2012__ = new_new_n1976__ & new_new_n2011__;
  assign new_new_n2013__ = ~new_new_n1976__ & ~new_new_n2011__;
  assign \r[27]  = new_new_n2012__ | new_new_n2013__;
  assign new_new_n2015__ = new_new_n1969__ & new_new_n2011__;
  assign new_new_n2016__ = new_new_n1873__ & new_new_n1926__;
  assign new_new_n2017__ = new_new_n2015__ & new_new_n2016__;
  assign new_new_n2018__ = ~new_new_n1814__ & new_new_n2017__;
  assign new_new_n2019__ = new_new_n1967__ & ~new_new_n2009__;
  assign new_new_n2020__ = ~new_new_n1924__ & ~new_new_n1970__;
  assign new_new_n2021__ = new_new_n2015__ & new_new_n2020__;
  assign new_new_n2022__ = ~new_new_n2010__ & ~new_new_n2019__;
  assign new_new_n2023__ = ~new_new_n2021__ & new_new_n2022__;
  assign new_new_n2024__ = ~new_new_n2018__ & new_new_n2023__;
  assign new_new_n2025__ = ~new_new_n2003__ & ~new_new_n2006__;
  assign new_new_n2026__ = ~new_new_n1982__ & ~new_new_n1984__;
  assign new_new_n2027__ = \a[13]  & \b[15] ;
  assign new_new_n2028__ = new_new_n1992__ & new_new_n1998__;
  assign new_new_n2029__ = ~new_new_n1992__ & ~new_new_n1998__;
  assign new_new_n2030__ = ~new_new_n2028__ & ~new_new_n2029__;
  assign new_new_n2031__ = ~new_new_n1994__ & ~new_new_n2030__;
  assign new_new_n2032__ = new_new_n2027__ & ~new_new_n2031__;
  assign new_new_n2033__ = ~new_new_n2027__ & new_new_n2031__;
  assign new_new_n2034__ = ~new_new_n2032__ & ~new_new_n2033__;
  assign new_new_n2035__ = \a[15]  & \b[13] ;
  assign new_new_n2036__ = \a[14]  & \b[14] ;
  assign new_new_n2037__ = ~new_new_n2035__ & ~new_new_n2036__;
  assign new_new_n2038__ = new_new_n2035__ & new_new_n2036__;
  assign new_new_n2039__ = ~new_new_n2037__ & ~new_new_n2038__;
  assign new_new_n2040__ = ~new_new_n2034__ & ~new_new_n2039__;
  assign new_new_n2041__ = new_new_n2034__ & new_new_n2039__;
  assign new_new_n2042__ = ~new_new_n2040__ & ~new_new_n2041__;
  assign new_new_n2043__ = new_new_n2000__ & new_new_n2042__;
  assign new_new_n2044__ = ~new_new_n2000__ & ~new_new_n2042__;
  assign new_new_n2045__ = ~new_new_n2043__ & ~new_new_n2044__;
  assign new_new_n2046__ = new_new_n2026__ & ~new_new_n2045__;
  assign new_new_n2047__ = ~new_new_n2026__ & new_new_n2045__;
  assign new_new_n2048__ = ~new_new_n2046__ & ~new_new_n2047__;
  assign new_new_n2049__ = new_new_n2025__ & ~new_new_n2048__;
  assign new_new_n2050__ = ~new_new_n2025__ & new_new_n2048__;
  assign new_new_n2051__ = ~new_new_n2049__ & ~new_new_n2050__;
  assign new_new_n2052__ = ~new_new_n2024__ & new_new_n2051__;
  assign new_new_n2053__ = new_new_n2024__ & ~new_new_n2051__;
  assign \r[28]  = ~new_new_n2052__ & ~new_new_n2053__;
  assign new_new_n2055__ = ~new_new_n2050__ & ~new_new_n2052__;
  assign new_new_n2056__ = ~new_new_n2043__ & ~new_new_n2047__;
  assign new_new_n2057__ = ~new_new_n2028__ & ~new_new_n2032__;
  assign new_new_n2058__ = \a[15]  & \b[14] ;
  assign new_new_n2059__ = \a[14]  & \b[15] ;
  assign new_new_n2060__ = ~new_new_n2058__ & ~new_new_n2059__;
  assign new_new_n2061__ = new_new_n2058__ & new_new_n2059__;
  assign new_new_n2062__ = \b[13]  & new_new_n2061__;
  assign new_new_n2063__ = ~new_new_n2038__ & ~new_new_n2059__;
  assign new_new_n2064__ = new_new_n2058__ & ~new_new_n2063__;
  assign new_new_n2065__ = ~new_new_n2062__ & new_new_n2064__;
  assign new_new_n2066__ = ~new_new_n2060__ & ~new_new_n2065__;
  assign new_new_n2067__ = new_new_n2041__ & new_new_n2066__;
  assign new_new_n2068__ = ~new_new_n2041__ & ~new_new_n2066__;
  assign new_new_n2069__ = ~new_new_n2067__ & ~new_new_n2068__;
  assign new_new_n2070__ = new_new_n2057__ & ~new_new_n2069__;
  assign new_new_n2071__ = ~new_new_n2057__ & new_new_n2069__;
  assign new_new_n2072__ = ~new_new_n2070__ & ~new_new_n2071__;
  assign new_new_n2073__ = new_new_n2056__ & ~new_new_n2072__;
  assign new_new_n2074__ = ~new_new_n2056__ & new_new_n2072__;
  assign new_new_n2075__ = ~new_new_n2073__ & ~new_new_n2074__;
  assign new_new_n2076__ = new_new_n2055__ & new_new_n2075__;
  assign new_new_n2077__ = ~new_new_n2055__ & ~new_new_n2075__;
  assign \r[29]  = new_new_n2076__ | new_new_n2077__;
  assign new_new_n2079__ = new_new_n2051__ & new_new_n2075__;
  assign new_new_n2080__ = ~new_new_n2024__ & new_new_n2079__;
  assign new_new_n2081__ = ~new_new_n2050__ & ~new_new_n2074__;
  assign new_new_n2082__ = ~new_new_n2073__ & ~new_new_n2081__;
  assign new_new_n2083__ = ~new_new_n2080__ & ~new_new_n2082__;
  assign new_new_n2084__ = ~new_new_n2067__ & ~new_new_n2071__;
  assign new_new_n2085__ = \a[15]  & \b[15] ;
  assign new_new_n2086__ = ~new_new_n2064__ & ~new_new_n2085__;
  assign new_new_n2087__ = ~new_new_n2061__ & ~new_new_n2086__;
  assign new_new_n2088__ = new_new_n2084__ & ~new_new_n2087__;
  assign new_new_n2089__ = ~new_new_n2084__ & new_new_n2087__;
  assign new_new_n2090__ = ~new_new_n2088__ & ~new_new_n2089__;
  assign new_new_n2091__ = ~new_new_n2083__ & new_new_n2090__;
  assign new_new_n2092__ = new_new_n2083__ & ~new_new_n2090__;
  assign \r[30]  = ~new_new_n2091__ & ~new_new_n2092__;
  assign new_new_n2094__ = ~new_new_n2061__ & new_new_n2091__;
  assign new_new_n2095__ = ~new_new_n2061__ & ~new_new_n2089__;
  assign new_new_n2096__ = ~new_new_n2091__ & ~new_new_n2095__;
  assign \r[31]  = new_new_n2094__ | new_new_n2096__;
endmodule


