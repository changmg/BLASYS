module max_7(pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 , pi11 , po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 );
  input pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , pi10 , pi11 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 ;
  wire new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33, new_n34, new_n35, new_n36, new_n37, new_n38, new_n39, new_n40, new_n41, new_n42, new_n43, new_n44, new_n45;
  assign new_n13 = ~pi00 & pi05 ;
  assign new_n14 = pi01 & ~pi06 ;
  assign new_n15 = pi00 & ~pi05 ;
  assign new_n16 = ~new_n14 & ~new_n15 ;
  assign new_n17 = ~pi10 & new_n16 ;
  assign new_n18 = ~pi02 & pi07 ;
  assign new_n19 = ~pi01 & pi06 ;
  assign new_n20 = ~new_n18 & ~new_n19 ;
  assign new_n21 = ~new_n17 & new_n20 ;
  assign new_n22 = pi03 & ~pi08 ;
  assign new_n23 = pi02 & ~pi07 ;
  assign new_n24 = ~new_n22 & ~new_n23 ;
  assign new_n25 = ~new_n21 & new_n24 ;
  assign new_n26 = ~pi04 & pi09 ;
  assign new_n27 = ~pi03 & pi08 ;
  assign new_n28 = ~new_n26 & ~new_n27 ;
  assign new_n29 = ~new_n25 & new_n28 ;
  assign new_n30 = pi04 & ~pi09 ;
  assign new_n31 = pi04 & pi11 ;
  assign new_n32 = pi09 & ~pi11 ;
  assign new_n33 = ~new_n31 & ~new_n32 ;
  assign new_n34 = pi00 & pi11 ;
  assign new_n35 = pi05 & ~pi11 ;
  assign new_n36 = ~new_n34 & ~new_n35 ;
  assign new_n37 = pi01 & pi11 ;
  assign new_n38 = pi06 & ~pi11 ;
  assign new_n39 = ~new_n37 & ~new_n38 ;
  assign new_n40 = pi02 & pi11 ;
  assign new_n41 = pi07 & ~pi11 ;
  assign new_n42 = ~new_n40 & ~new_n41 ;
  assign new_n43 = pi03 & pi11 ;
  assign new_n44 = pi08 & ~pi11 ;
  assign new_n45 = ~new_n43 & ~new_n44 ;
  assign po0 = new_n13 ;
  assign po1 = new_n29 ;
  assign po2 = new_n30 ;
  assign po3 = new_n33 ;
  assign po4 = new_n36 ;
  assign po5 = new_n39 ;
  assign po6 = new_n42 ;
  assign po7 = new_n45 ;
endmodule
