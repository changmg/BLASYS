module max_14_2(pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 , po0 , po1 , po2 , po3 );
  input pi00 , pi01 , pi02 , pi03 , pi04 , pi05 , pi06 , pi07 , pi08 , pi09 ;
  output po0 , po1 , po2 , po3 ;
  wire new_n11, new_n12, new_n13, new_n14, new_n15, new_n16, new_n17, new_n18, new_n19, new_n20, new_n21, new_n22, new_n23, new_n24, new_n25, new_n26, new_n27, new_n28, new_n29, new_n30, new_n31, new_n32, new_n33;
  assign new_n11 = pi01 & ~pi06 ;
  assign new_n12 = ~pi07 & ~new_n11 ;
  assign new_n13 = ~pi00 & new_n12 ;
  assign new_n14 = ~pi02 & pi08 ;
  assign new_n15 = ~pi01 & pi06 ;
  assign new_n16 = ~new_n14 & ~new_n15 ;
  assign new_n17 = ~new_n13 & new_n16 ;
  assign new_n18 = pi02 & ~pi08 ;
  assign new_n19 = pi03 & ~pi09 ;
  assign new_n20 = ~new_n18 & ~new_n19 ;
  assign new_n21 = ~new_n17 & new_n20 ;
  assign new_n22 = ~pi03 & pi09 ;
  assign new_n23 = ~pi04 & ~new_n22 ;
  assign new_n24 = ~new_n21 & new_n23 ;
  assign new_n25 = ~pi01 & pi05 ;
  assign new_n26 = ~pi05 & ~pi06 ;
  assign new_n27 = ~new_n25 & ~new_n26 ;
  assign new_n28 = ~pi02 & pi05 ;
  assign new_n29 = ~pi05 & ~pi08 ;
  assign new_n30 = ~new_n28 & ~new_n29 ;
  assign new_n31 = ~pi03 & pi05 ;
  assign new_n32 = ~pi05 & ~pi09 ;
  assign new_n33 = ~new_n31 & ~new_n32 ;
  assign po0 = new_n24 ;
  assign po1 = new_n27 ;
  assign po2 = new_n30 ;
  assign po3 = new_n33 ;
endmodule
