// Benchmark "ex" written by ABC on Thu Jul 14 00:22:41 2022

module ex ( 
    a, b, c, d, e, f, g, h, i, j, k, l,
    F  );
  input  a, b, c, d, e, f, g, h, i, j, k, l;
  output F;
  assign F = ~a & f;
endmodule


